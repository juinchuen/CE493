* NGSPICE file created from top.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X12 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X13 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X14 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
.ends

.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0683 ps=0.86 w=0.65 l=0.15
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
X0 VGND A2 a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0683 ps=0.86 w=0.65 l=0.15
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A1 a_114_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X3 a_114_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.185 ps=1.87 w=0.65 l=0.15
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X8 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X10 a_285_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
X11 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
X0 a_222_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X1 VPWR A1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X2 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_222_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.186 ps=1.41 w=0.42 l=0.15
X4 VGND A2 a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X5 a_448_47# a_222_93# a_79_199# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_79_199# a_222_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X7 a_544_297# A2 a_79_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8 a_448_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.41 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 a_78_199# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2 a_493_297# A2 a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X3 VPWR a_78_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.373 pd=1.75 as=0.28 ps=2.56 w=1 l=0.15
X4 VGND A2 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X5 a_78_199# B2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.117 ps=1.24 w=1 l=0.15
X6 a_215_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_215_47# B2 a_78_199# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_292_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.117 pd=1.24 as=0.373 ps=1.75 w=1 l=0.15
X9 VGND a_78_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
X0 a_27_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_560_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2 VGND B a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0991 ps=0.955 w=0.65 l=0.15
X3 Y B a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y a_27_297# a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_474_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X7 VGND A a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_27_47# B a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_27_297# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VPWR B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X12 a_474_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_560_47# a_27_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14 VPWR A a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X15 Y a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X16 VPWR a_27_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X17 a_560_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
X0 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_470_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_470_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_470_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.106 ps=0.975 w=0.65 l=0.15
X6 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X8 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X10 a_470_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.162 ps=1.33 w=1 l=0.15
X11 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 VPWR B a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X13 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VGND A a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X16 X a_112_47# a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 a_470_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X18 X B a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 a_585_47# B1 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.119 ps=1.01 w=0.65 l=0.15
X1 VGND A2 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.137 pd=1.07 as=0.117 ps=1.01 w=0.65 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.62 as=0.26 ps=2.52 w=1 l=0.15
X3 a_81_21# C1 a_585_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.203 pd=1.27 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_266_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.312 ps=1.62 w=1 l=0.15
X6 a_368_297# A2 a_266_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.18 ps=1.36 w=1 l=0.15
X7 a_266_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.137 ps=1.07 w=0.65 l=0.15
X8 a_266_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.203 ps=1.27 w=0.65 l=0.15
X9 a_81_21# A3 a_368_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.21 ps=1.42 w=1 l=0.15
X10 a_81_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X11 VPWR B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.138 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
X0 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X1 Y a_27_93# a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_206_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X3 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X5 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 a_240_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_51_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VGND A1 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_51_297# B2 a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.412 pd=1.83 as=0.105 ps=1.21 w=1 l=0.15
X4 a_149_47# C1 a_51_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.201 ps=1.92 w=0.65 l=0.15
X5 a_240_47# B1 a_149_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0991 ps=0.955 w=0.65 l=0.15
X6 VPWR A1 a_512_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X7 X a_51_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
X8 a_149_47# B2 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_245_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X10 VPWR C1 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X11 a_512_297# A2 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.412 ps=1.83 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
X0 a_219_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.157 ps=1.17 w=0.42 l=0.15
X1 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.157 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VPWR A a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 X a_219_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_301_297# a_27_53# a_219_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5 X a_219_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X6 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_219_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
X0 VGND A2 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X1 Y B1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 VPWR A1 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15
X4 a_29_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y A2 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND A1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X7 a_112_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X8 a_112_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.14 ps=1.28 w=1 l=0.15
X9 a_29_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X11 a_29_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.127 ps=1.04 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
X0 VPWR A a_49_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VGND a_285_47# a_391_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.5
X2 X a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VGND A a_49_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VPWR a_285_47# a_391_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.5
X5 a_285_47# a_49_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X6 a_285_47# a_49_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X7 X a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.167 ps=1.43 w=0.42 l=0.15
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.139 ps=1.08 w=0.42 l=0.15
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.12 ps=1.09 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.43 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.09 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
X0 a_298_297# a_27_413# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1 a_215_297# a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.136 ps=1.1 w=0.65 l=0.15
X2 a_298_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.258 ps=1.45 w=0.65 l=0.15
X4 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6 a_382_47# A1 a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.136 pd=1.1 as=0.111 ps=1.37 w=0.42 l=0.15
X8 VPWR A1 a_298_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND A2 a_382_47# VNB sky130_fd_pr__nfet_01v8 ad=0.258 pd=1.45 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
X0 a_277_47# a_247_21# a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VGND S0 a_247_21# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_834_97# a_247_21# a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VGND A3 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X4 a_1290_413# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_834_97# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_750_97# S0 a_757_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X7 a_27_47# S0 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0852 ps=0.925 w=0.42 l=0.15
X8 X a_1478_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR A1 a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10 VPWR S0 a_247_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.108 pd=1.36 as=0.108 ps=1.36 w=0.42 l=0.15
X11 X a_1478_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X12 a_193_47# A0 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_750_97# a_1290_413# a_1478_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.269 pd=2.12 as=0.0921 ps=0.99 w=0.42 l=0.15
X14 a_1478_413# S1 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0921 pd=0.99 as=0.109 ps=1.36 w=0.42 l=0.15
X15 a_1290_413# S1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X16 a_277_47# a_247_21# a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0852 pd=0.925 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_750_97# S0 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X18 a_923_363# a_247_21# a_750_97# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0901 pd=0.995 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 a_757_363# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 VPWR A3 a_923_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0901 ps=0.995 w=0.42 l=0.15
X21 a_277_47# a_1290_413# a_1478_413# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.151 ps=1.28 w=0.42 l=0.15
X22 a_193_413# A0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X23 a_193_413# S0 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.108 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X24 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X25 a_1478_413# S1 a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0.151 pd=1.28 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 VGND A1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_510_47# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X2 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X3 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X4 a_79_21# A2 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.162 ps=1.33 w=1 l=0.15
X5 a_297_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X6 a_79_21# C1 a_510_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.114 ps=1 w=0.65 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 a_215_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.106 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.92 as=0.107 ps=0.98 w=0.65 l=0.15
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.213 ps=1.42 w=1 l=0.15
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.127 ps=1.04 w=0.65 l=0.15
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.108 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122 ps=1.08 w=0.65 l=0.15
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.0536 ps=0.675 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.172 ps=1.83 w=0.65 l=0.15
X2 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X3 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X4 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X5 a_326_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.127 ps=1.04 w=0.65 l=0.15
X6 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.635 pd=3.27 as=0.195 ps=1.39 w=1 l=0.15
X7 Y C1 a_326_47# VNB sky130_fd_pr__nfet_01v8 ad=0.393 pd=2.51 as=0.0683 ps=0.86 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 a_286_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2 a_286_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.185 ps=1.87 w=0.65 l=0.15
X3 Y A2 a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 VGND A1 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.185 ps=1.87 w=0.65 l=0.15
X6 VGND A2 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7 a_487_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 a_27_47# B1 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10 VPWR A1 a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X13 a_487_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X14 a_286_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X15 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
X0 Y A1 a_194_47# VNB sky130_fd_pr__nfet_01v8 ad=0.115 pd=1 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_194_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X2 Y C1 a_376_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.35 w=1 l=0.15
X3 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.112 ps=0.995 w=0.65 l=0.15
X5 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.115 ps=1 w=0.65 l=0.15
X6 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X7 a_376_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.165 ps=1.33 w=1 l=0.15
X8 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X2 a_193_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 Y A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 a_109_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.117 ps=1.01 w=0.65 l=0.15
X1 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.41 pd=1.82 as=0.135 ps=1.27 w=1 l=0.15
X2 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.175 ps=1.35 w=1 l=0.15
X4 a_277_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_27_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.41 ps=1.82 w=1 l=0.15
X10 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.18 ps=1.36 w=1 l=0.15
X11 a_277_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X13 Y A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.0975 ps=0.95 w=0.65 l=0.15
X14 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 Y a_61_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.183 ps=1.24 w=0.65 l=0.15
X1 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_217_297# a_61_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_479_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X4 a_217_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X5 Y a_61_47# a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VPWR A1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_61_47# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=0.15
X8 VGND A2 a_637_47# VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND a_61_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 Y A1 a_479_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0683 ps=0.86 w=0.65 l=0.15
X11 VGND B1_N a_61_47# VNB sky130_fd_pr__nfet_01v8 ad=0.183 pd=1.24 as=0.126 ps=1.44 w=0.42 l=0.15
X12 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X13 a_637_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
X0 Y a_53_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.192 ps=1.38 w=1 l=0.15
X1 a_232_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.192 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A_N a_53_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VGND A_N a_53_93# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_316_47# B a_232_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.03 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 Y a_53_93# a_316_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.125 ps=1.03 w=0.65 l=0.15
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 a_75_199# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.135 ps=1.07 w=0.65 l=0.15
X1 a_208_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.03 as=0.112 ps=0.995 w=0.65 l=0.15
X2 a_315_47# A2 a_208_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.125 ps=1.03 w=0.65 l=0.15
X3 VGND B1 a_75_199# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.07 as=0.106 ps=0.975 w=0.65 l=0.15
X4 a_75_199# A1 a_315_47# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.17 w=0.65 l=0.15
X5 a_75_199# C1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.207 ps=1.41 w=1 l=0.15
X6 a_544_297# B1 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.207 pd=1.41 as=0.162 ps=1.33 w=1 l=0.15
X7 VPWR a_75_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X8 a_201_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.142 ps=1.28 w=1 l=0.15
X9 VPWR A2 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.165 ps=1.33 w=1 l=0.15
X10 a_201_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.305 ps=1.61 w=1 l=0.15
X11 VGND a_75_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 a_388_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.25 as=0.153 ps=1.3 w=1 l=0.15
X1 a_105_352# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_297_47# a_105_352# Y VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VPWR A1 a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.127 ps=1.25 w=1 l=0.15
X5 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X6 VPWR B1_N a_105_352# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X7 Y a_105_352# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.178 ps=1.4 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 a_77_199# B2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.06 as=0.127 ps=1.04 w=0.65 l=0.15
X1 a_323_297# A2 a_227_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X2 a_227_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_227_47# B1 a_77_199# VNB sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.133 ps=1.06 w=0.65 l=0.15
X4 VGND a_77_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VPWR B1 a_539_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.205 ps=1.41 w=1 l=0.15
X6 a_227_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X7 VPWR a_77_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X8 a_77_199# A3 a_323_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X9 VGND A2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.107 ps=0.98 w=0.65 l=0.15
X10 a_227_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_539_297# B2 a_77_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.195 ps=1.39 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X9 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X12 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X14 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X15 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X16 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X17 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X18 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X22 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X23 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X24 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X25 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X26 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X27 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X29 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
X0 a_109_93# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 a_215_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VGND a_109_93# a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3 VGND A a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VPWR A a_369_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 a_369_297# B a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_215_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X7 a_297_297# a_109_93# a_215_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_109_93# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X9 X a_215_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.1 ps=0.985 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_206_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.146 ps=1.34 w=0.42 l=0.15
X1 a_206_369# A2_N a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X2 VGND B2 a_489_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_585_369# B2 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0672 ps=0.74 w=0.42 l=0.15
X4 a_489_47# a_206_369# a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_489_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VPWR A2_N a_206_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.209 pd=1.35 as=0.129 ps=1.18 w=0.42 l=0.15
X7 a_76_199# a_206_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.209 ps=1.35 w=0.42 l=0.15
X8 a_205_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0662 pd=0.735 as=0.0986 ps=0.98 w=0.42 l=0.15
X9 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X10 VPWR B1 a_585_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.0986 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
X0 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_806_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_806_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_806_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 X B a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 X a_112_47# a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_806_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND A a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 X B a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 VGND A a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_806_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.272 ps=2.56 w=1 l=0.15
X15 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X17 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X19 a_806_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR B a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 VPWR B a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X24 a_806_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 a_806_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X28 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 a_806_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.257 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X30 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 VPWR A a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 X a_112_47# a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X35 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 a_806_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X38 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X39 VPWR A a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 a_676_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.213 ps=1.42 w=1 l=0.15
X1 a_512_47# B1 a_409_47# VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.26 as=0.119 ps=1.01 w=0.65 l=0.15
X2 a_306_47# D1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.198 ps=1.91 w=0.65 l=0.15
X3 VGND A2 a_512_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.198 ps=1.26 w=0.65 l=0.15
X4 VPWR C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.218 ps=1.43 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.42 as=0.305 ps=1.61 w=1 l=0.15
X6 VPWR A1 a_676_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X7 a_512_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_409_47# C1 a_306_47# VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.119 ps=1.01 w=0.65 l=0.15
X9 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.382 pd=1.76 as=0.26 ps=2.52 w=1 l=0.15
X10 a_79_21# D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=1.43 as=0.382 ps=1.76 w=1 l=0.15
X11 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 a_300_297# a_27_413# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=0.15
X3 Y a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.102 ps=0.99 w=0.65 l=0.15
X4 VPWR A1 a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 a_384_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.143 ps=1.09 w=0.65 l=0.15
X6 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.111 ps=1.37 w=0.42 l=0.15
X7 a_300_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 VPWR a_38_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A1 a_497_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X2 X a_38_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X3 a_141_47# B2 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_497_297# A2 a_38_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.387 ps=1.77 w=1 l=0.15
X5 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR C1 a_38_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.325 ps=2.65 w=1 l=0.15
X7 a_237_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.112 pd=1.23 as=0.165 ps=1.33 w=1 l=0.15
X8 a_38_47# B2 a_237_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.387 pd=1.77 as=0.112 ps=1.23 w=1 l=0.15
X9 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 X a_38_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_141_47# C1 a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.237 ps=2.03 w=0.65 l=0.15
X12 VGND a_38_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_225_47# B1 a_141_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
X0 a_121_297# B a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_39_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=1 w=0.65 l=0.15
X2 VPWR a_39_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_39_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.156 ps=1.36 w=1 l=0.15
X4 VGND a_39_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.156 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VGND A a_39_297# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=1 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_39_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X1 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_215_297# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_392_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0452 pd=0.635 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 a_465_297# B a_392_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.064 pd=0.725 as=0.0452 ps=0.635 w=0.42 l=0.15
X6 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR A a_465_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.064 ps=0.725 w=0.42 l=0.15
X8 a_297_297# a_109_53# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.064 ps=0.725 w=0.42 l=0.15
X11 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 VGND A2 a_660_47# VNB sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X1 VGND C1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X2 a_414_297# C1 a_334_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X3 VGND a_85_193# X VNB sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X4 a_334_297# D1 a_85_193# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X5 a_516_297# B1 a_414_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X6 a_516_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7 a_660_47# A1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X8 a_85_193# D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X9 VPWR A1 a_516_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X10 a_85_193# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X11 VPWR a_85_193# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 a_465_47# A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VGND A4 a_561_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X2 VPWR A3 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3 a_297_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4 a_297_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X5 VPWR A1 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_381_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.184 ps=1.22 w=0.65 l=0.15
X7 a_297_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9 a_79_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.184 pd=1.22 as=0.161 ps=1.14 w=0.65 l=0.15
X10 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.161 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_561_47# A3 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
X0 VPWR S a_591_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X1 a_591_369# A0 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.131 ps=1.05 w=0.64 l=0.15
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.41 as=0.135 ps=1.27 w=1 l=0.15
X3 a_79_21# A1 a_306_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.131 pd=1.05 as=0.229 ps=1.36 w=0.64 l=0.15
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND S a_578_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0578 ps=0.695 w=0.42 l=0.15
X6 a_306_369# a_257_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.229 pd=1.36 as=0.178 ps=1.41 w=0.64 l=0.15
X7 a_79_21# A0 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=0.173 pd=1.25 as=0.0683 ps=0.745 w=0.42 l=0.15
X8 a_288_47# a_257_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X9 a_257_199# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_578_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.173 ps=1.25 w=0.42 l=0.15
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 a_257_199# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.173 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
X0 VGND C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_277_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_27_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X8 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_277_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X1 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X3 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_381_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VGND A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.0683 ps=0.86 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
X0 VGND A a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 Y a_38_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_38_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_820_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR a_38_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X5 VGND A a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND B a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND B a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y B a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_38_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_38_297# B a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VGND A a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_902_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_820_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_902_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 VPWR A a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 Y a_38_297# a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 Y a_38_297# a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 a_38_47# B a_38_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_38_47# B a_38_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 a_38_297# B a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X21 a_38_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 VPWR B a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X23 a_38_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X24 a_902_47# a_38_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 a_902_47# a_38_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 Y B a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_38_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 a_820_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VPWR A a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 VGND A a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 VPWR A a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 a_902_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X33 a_820_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 Y a_38_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X35 a_902_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X36 a_38_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 VPWR A a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X38 VPWR a_38_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X39 VPWR B a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.198 ps=1.26 w=0.65 l=0.15
X1 Y A3 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.393 pd=1.78 as=0.135 ps=1.27 w=1 l=0.15
X2 a_193_297# A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.393 ps=1.78 w=1 l=0.15
X5 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.26 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 Y A1 a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.119 ps=1.01 w=0.65 l=0.15
X1 a_181_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.0683 ps=0.86 w=0.65 l=0.15
X2 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.106 ps=0.975 w=0.65 l=0.15
X3 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.162 ps=1.33 w=1 l=0.15
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.153 ps=1.3 w=1 l=0.15
X6 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0483 pd=0.65 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X6 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X7 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.17 as=0.218 ps=2.2 w=0.84 l=0.15
X8 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X9 a_1224_47# a_27_47# a_1032_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VGND a_1032_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X12 VPWR a_1182_261# a_1140_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X13 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X14 a_1032_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X15 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.125 ps=1.17 w=0.42 l=0.15
X16 a_1296_47# a_1182_261# a_1224_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0483 pd=0.65 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X19 VPWR SET_B a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X20 a_1032_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0483 ps=0.65 w=0.42 l=0.15
X21 a_1182_261# a_1032_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.123 ps=1.17 w=0.84 l=0.15
X22 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1140_413# a_193_47# a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VPWR a_1032_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X26 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X27 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X28 a_1182_261# a_1032_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.6 as=0.114 ps=1.01 w=0.54 l=0.15
X29 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X30 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X31 VGND SET_B a_1296_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1.01 as=0.0483 ps=0.65 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0894 ps=0.925 w=0.65 l=0.15
X1 a_191_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X2 VPWR A a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.119 ps=1.01 w=0.65 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_297_297# B a_191_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X6 a_109_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.115 ps=1 w=0.65 l=0.15
X1 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.115 pd=1 as=0.0926 ps=0.935 w=0.65 l=0.15
X2 VPWR A1 a_307_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.105 ps=1.21 w=1 l=0.15
X3 a_307_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.233 ps=1.47 w=1 l=0.15
X4 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.233 pd=1.47 as=0.112 ps=1.23 w=1 l=0.15
X6 a_109_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.112 pd=1.23 as=0.26 ps=2.52 w=1 l=0.15
X7 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR A1 a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.16 ps=1.32 w=1 l=0.15
X1 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.4 ps=1.8 w=1 l=0.15
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0894 ps=0.925 w=0.65 l=0.15
X3 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_470_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=1.8 as=0.138 ps=1.27 w=1 l=0.15
X6 a_384_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X7 a_384_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.104 ps=0.97 w=0.65 l=0.15
X8 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 VGND A2 a_485_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 VPWR A1 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 a_37_297# B1 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_485_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_292_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X7 VPWR A2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8 a_485_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X11 a_37_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 Y A1 a_485_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X13 Y C1 a_37_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X14 a_292_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X15 a_292_297# B1 a_37_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_467_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_467_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A1 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_109_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND A2 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
X0 VPWR a_30_53# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.315 pd=2.63 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND a_30_53# X VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 X a_30_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148 ps=1.34 w=1 l=0.15
X3 a_112_297# C a_30_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4 X a_30_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X5 VGND A a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_30_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VGND C a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_184_297# B a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X9 VPWR A a_184_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_294_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0662 pd=0.735 as=0.0986 ps=0.98 w=0.42 l=0.15
X1 VPWR A2_N a_295_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.227 pd=1.35 as=0.173 ps=1.4 w=0.64 l=0.15
X2 VPWR B1 a_665_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.0986 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.185 ps=1.87 w=0.65 l=0.15
X5 a_581_47# a_295_369# a_84_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X7 a_665_369# B2 a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0928 ps=0.93 w=0.64 l=0.15
X8 VGND B2 a_581_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_295_369# A2_N a_294_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X10 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.285 ps=2.57 w=1 l=0.15
X11 a_84_21# a_295_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0928 pd=0.93 as=0.227 ps=1.35 w=0.64 l=0.15
X12 a_295_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.173 pd=1.4 as=0.154 ps=1.34 w=0.64 l=0.15
X13 a_581_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 a_109_47# B1 a_213_123# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.165 ps=1.82 w=0.65 l=0.15
X1 Y B2 a_295_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.12 ps=1.24 w=1 l=0.15
X2 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3 a_213_123# B2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_295_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12 pd=1.24 as=0.38 ps=1.76 w=1 l=0.15
X5 a_493_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.225 ps=1.45 w=1 l=0.15
X6 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=1.76 as=0.28 ps=2.56 w=1 l=0.15
X7 VGND A2 a_213_123# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.117 ps=1.01 w=0.65 l=0.15
X8 a_213_123# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_109_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
X0 VPWR A a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_218_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.156 ps=1.16 w=0.42 l=0.15
X2 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.156 pd=1.16 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_300_297# a_27_53# a_218_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4 X a_218_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X5 VPWR a_218_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X6 X a_218_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148 ps=1.34 w=1 l=0.15
X7 VGND a_218_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X9 VGND A a_218_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
X0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X7 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X13 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X14 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X16 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X17 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X18 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X19 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X20 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X21 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X22 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X23 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X9 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X12 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X15 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X16 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X17 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X18 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X19 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X28 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X29 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X30 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X31 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X32 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X33 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14 ps=1.28 w=1 l=0.15
X1 VGND A3 a_383_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X2 a_309_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0715 pd=0.87 as=0.153 ps=1.12 w=0.65 l=0.15
X3 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.153 pd=1.12 as=0.0747 ps=0.88 w=0.65 l=0.15
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X5 a_383_47# A2 a_309_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0715 ps=0.87 w=0.65 l=0.15
X6 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X7 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=1.67 w=1 l=0.15
X1 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0.194 pd=1.95 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VGND B a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 Y a_27_93# a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 a_229_47# a_27_93# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y a_27_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.147 ps=1.34 w=1 l=0.15
X6 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.165 ps=1.33 w=1 l=0.15
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X8 a_229_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 a_465_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_204_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0699 pd=0.865 as=0.106 ps=0.975 w=0.65 l=0.15
X4 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.91 as=0.0991 ps=0.955 w=0.65 l=0.15
X5 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.26 ps=2.52 w=1 l=0.15
X6 Y B1 a_204_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0699 ps=0.865 w=0.65 l=0.15
X7 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.153 ps=1.3 w=1 l=0.15
X8 a_109_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X11 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X18 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
X0 a_28_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 a_462_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 Y B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_462_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_28_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 a_462_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X7 Y B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y A1 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X11 a_28_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.145 ps=1.29 w=1 l=0.15
X12 VPWR A2 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X14 VGND A2 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X15 a_28_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X16 VPWR A1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X17 a_28_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 VGND A2 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X19 VPWR A2 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.155 ps=1.31 w=1 l=0.15
X20 a_28_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X21 Y A1 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X22 a_462_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X23 VPWR A1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
X0 a_297_47# a_27_47# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.103 ps=1 w=0.65 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0.103 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X6 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X8 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.128 ps=1.03 w=0.42 l=0.15
X9 a_193_413# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X11 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
X0 VPWR a_29_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_29_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.151 ps=1.35 w=1 l=0.15
X2 VPWR A a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3 VGND a_29_311# X VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_184_53# B a_112_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 VPWR C a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.151 pd=1.35 as=0.0744 ps=0.815 w=0.42 l=0.15
X6 X a_29_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.13 ps=1.11 w=0.65 l=0.15
X7 a_112_53# A a_29_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_29_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 VGND C a_184_53# VNB sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.11 as=0.0536 ps=0.675 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X2 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.338 pd=1.67 as=0.135 ps=1.27 w=1 l=0.15
X5 a_1249_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_1249_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.252 pd=1.5 as=0.338 ps=1.67 w=1 l=0.15
X12 a_803_47# A2 a_1249_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X16 a_803_47# A2 a_1249_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X20 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X21 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 a_1249_47# A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.133 ps=1.06 w=0.65 l=0.15
X23 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 a_1249_47# A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.252 ps=1.5 w=1 l=0.15
X28 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.06 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X30 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X32 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X33 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X35 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 VGND A3 a_1249_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X37 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X38 VGND A3 a_1249_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X39 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 a_56_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR A2 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
X3 a_139_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.266 ps=2.12 w=0.65 l=0.15
X4 a_311_297# B1 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X5 Y C1 a_311_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X6 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X7 Y A1 a_139_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
X0 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X1 a_471_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.42 pd=2.84 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_27_47# C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=1.67 w=1 l=0.15
X8 a_277_47# B a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X9 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.135 ps=1.27 w=1 l=0.15
X10 Y A a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_277_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X13 a_471_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 a_79_21# C1 a_635_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.21 ps=1.42 w=1 l=0.15
X1 VPWR A2 a_319_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.17 ps=1.34 w=1 l=0.15
X2 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.08 as=0.133 ps=1.06 w=0.65 l=0.15
X3 a_417_47# A2 a_319_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.02 as=0.111 ps=0.99 w=0.65 l=0.15
X4 a_79_21# A1 a_417_47# VNB sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.06 as=0.12 ps=1.02 w=0.65 l=0.15
X5 a_319_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.111 pd=0.99 as=0.156 ps=1.13 w=0.65 l=0.15
X6 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.24 pd=1.48 as=0.135 ps=1.27 w=1 l=0.15
X7 a_319_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.185 ps=1.37 w=1 l=0.15
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.156 pd=1.13 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_319_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.34 as=0.24 ps=1.48 w=1 l=0.15
X10 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.14 ps=1.08 w=0.65 l=0.15
X11 a_635_297# B1 a_319_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.21 ps=1.42 w=1 l=0.15
X12 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
X0 Y a_74_47# a_265_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR B_N a_74_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.39 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_265_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.157 ps=1.39 w=1 l=0.15
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X4 VGND B_N a_74_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VGND a_74_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.91 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148 ps=1.34 w=1 l=0.15
X9 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
X0 a_600_345# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1 a_788_316# S1 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VPWR A3 a_372_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.164 ps=1.33 w=0.64 l=0.15
X3 a_872_316# a_600_345# a_788_316# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X4 VPWR S0 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5 a_1279_413# S0 a_872_316# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=0.995 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND a_788_316# X VNB sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_1060_369# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.16 as=0.166 ps=1.8 w=0.64 l=0.15
X8 a_872_316# a_27_47# a_1060_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.138 ps=1.16 w=0.42 l=0.15
X9 a_1281_47# a_27_47# a_872_316# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.072 ps=0.76 w=0.36 l=0.15
X10 a_193_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_1064_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0786 pd=0.805 as=0.109 ps=1.36 w=0.42 l=0.15
X12 a_872_316# S1 a_788_316# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.6 as=0.0729 ps=0.81 w=0.54 l=0.15
X13 a_872_316# S0 a_1064_47# VNB sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0786 ps=0.805 w=0.36 l=0.15
X14 X a_788_316# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=1 w=0.65 l=0.15
X15 a_788_316# a_600_345# a_288_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0729 pd=0.81 as=0.14 ps=1.6 w=0.54 l=0.15
X16 a_372_413# a_27_47# a_288_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.164 pd=1.33 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VGND A3 a_397_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.0671 ps=0.75 w=0.42 l=0.15
X18 a_600_345# S1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0819 ps=0.81 w=0.42 l=0.15
X19 a_193_369# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0957 pd=0.965 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 VPWR a_788_316# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.135 ps=1.27 w=1 l=0.15
X21 a_288_47# S0 a_193_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0957 ps=0.965 w=0.42 l=0.15
X22 a_397_47# S0 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X23 VGND A0 a_1281_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=1 as=0.066 ps=0.745 w=0.42 l=0.15
X24 a_288_47# a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X25 X a_788_316# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.154 ps=1.34 w=1 l=0.15
X26 VGND S0 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X27 VPWR A0 a_1279_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.105 ps=0.995 w=0.64 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR a_80_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1 X a_80_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 VGND a_80_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.111 pd=0.99 as=0.091 ps=0.93 w=0.65 l=0.15
X3 a_386_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X4 X a_80_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X5 a_80_199# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.162 pd=1.15 as=0.111 ps=0.99 w=0.65 l=0.15
X6 a_386_297# B1 a_80_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_458_47# A1 a_80_199# VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.162 ps=1.15 w=0.65 l=0.15
X8 VPWR A1 a_386_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X9 VGND A2 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.123 ps=1.03 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
X0 VPWR A1 a_485_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_485_297# a_297_93# a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 a_297_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.108 ps=1.01 w=0.42 l=0.15
X3 a_581_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.01 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_79_21# a_297_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6 VGND A2 a_581_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.51 as=0.14 ps=1.28 w=1 l=0.15
X8 a_297_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.182 ps=1.51 w=0.42 l=0.15
X9 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X10 a_485_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_475_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR A1 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X9 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.27 pd=1.48 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X12 a_475_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 Y A2 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X14 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.27 ps=1.48 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 Y A2 a_734_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_300_47# B2 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 a_300_47# B1 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_300_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_734_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X7 a_28_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y C1 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR B1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X11 a_382_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_28_47# B1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_28_47# B2 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VGND A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X15 Y B2 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 VPWR A1 a_734_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND A2 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 a_382_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X19 a_734_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 a_281_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1 a_281_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.26 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X7 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X9 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.127 ps=1.04 w=0.65 l=0.15
X10 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.198 ps=1.26 w=0.65 l=0.15
X11 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.127 ps=1.04 w=0.65 l=0.15
X12 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 Y A3 a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.195 ps=1.39 w=1 l=0.15
X15 a_27_297# A2 a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
X0 VPWR D a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_223_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.5 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 a_515_93# a_223_47# a_429_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 a_223_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.134 pd=1.48 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X5 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X6 X a_343_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.46 w=1 l=0.15
X7 a_429_93# a_27_47# a_343_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.118 ps=1.4 w=0.42 l=0.15
X8 VGND D a_615_93# VNB sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.11 as=0.0777 ps=0.79 w=0.42 l=0.15
X9 a_343_93# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X10 a_343_93# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X11 a_615_93# C a_515_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X12 X a_343_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.82 as=0.126 ps=1.11 w=0.65 l=0.15
X13 VPWR a_223_47# a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
X0 VGND a_91_199# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VPWR A a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X3 a_91_199# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_245_297# B a_161_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_91_199# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.146 ps=1.34 w=0.42 l=0.15
X7 a_161_297# a_91_199# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
X0 VGND A a_311_413# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 VPWR A a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0598 ps=0.705 w=0.42 l=0.15
X2 a_393_413# a_205_93# a_311_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X3 VGND C_N a_27_410# VNB sky130_fd_pr__nfet_01v8 ad=0.0619 pd=0.715 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VPWR C_N a_27_410# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.32 as=0.109 ps=1.36 w=0.42 l=0.15
X5 X a_311_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X6 VGND a_27_410# a_311_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0598 ps=0.705 w=0.42 l=0.15
X7 a_561_297# B a_489_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0598 pd=0.705 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 a_205_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0619 ps=0.715 w=0.42 l=0.15
X9 a_205_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.123 ps=1.32 w=0.42 l=0.15
X10 a_489_297# a_27_410# a_393_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.122 ps=1.33 w=0.42 l=0.15
X11 a_311_413# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_311_413# a_205_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0598 pd=0.705 as=0.109 ps=1.36 w=0.42 l=0.15
X13 X a_311_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.102 ps=0.99 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 a_1224_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VPWR A1 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.183 ps=1.37 w=1 l=0.15
X2 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_806_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.205 ps=1.28 w=0.65 l=0.15
X8 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.205 pd=1.28 as=0.14 ps=1.08 w=0.65 l=0.15
X10 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_806_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 Y A3 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 Y A3 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X19 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.119 ps=1.01 w=0.65 l=0.15
X22 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0926 ps=0.935 w=0.65 l=0.15
X24 a_806_297# A2 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X25 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.142 ps=1.28 w=1 l=0.15
X28 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.08 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 a_1224_297# A2 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 a_1224_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.135 ps=1.27 w=1 l=0.15
X32 a_806_297# A2 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 VPWR A1 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X35 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X36 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X37 a_1224_297# A2 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X38 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X39 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
X0 a_149_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_757_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_757_47# A3 a_567_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VPWR A3 a_149_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=1.77 as=0.145 ps=1.29 w=1 l=0.15
X4 Y B1 a_149_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_567_47# A3 a_757_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VGND A4 a_757_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A4 a_149_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_149_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_317_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_317_47# A2 a_567_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_149_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.385 ps=1.77 w=1 l=0.15
X13 a_149_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X14 Y A1 a_317_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 VPWR A2 a_149_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_567_47# A2 a_317_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 a_149_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 VPWR A1 a_149_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.192 ps=1.38 w=1 l=0.15
X1 a_232_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.118 ps=1.04 w=0.65 l=0.15
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.192 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A_N a_41_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VPWR a_41_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.195 ps=1.39 w=1 l=0.15
X5 a_316_47# C a_232_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.03 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 Y a_41_93# a_423_47# VNB sky130_fd_pr__nfet_01v8 ad=0.228 pd=2 as=0.127 ps=1.04 w=0.65 l=0.15
X7 a_423_47# B a_316_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.125 ps=1.03 w=0.65 l=0.15
X8 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X9 VGND A_N a_41_93# VNB sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.04 as=0.111 ps=1.37 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.14 ps=1.28 w=1 l=0.15
X1 a_235_47# C1 a_163_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.0683 ps=0.86 w=0.65 l=0.15
X2 a_343_47# B1 a_235_47# VNB sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.05 as=0.127 ps=1.04 w=0.65 l=0.15
X3 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.203 pd=1.4 as=0.195 ps=1.39 w=1 l=0.15
X4 a_454_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.203 ps=1.4 w=1 l=0.15
X5 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6 VPWR A1 a_454_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.195 ps=1.39 w=1 l=0.15
X7 a_163_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X8 VGND A2 a_343_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.132 ps=1.05 w=0.65 l=0.15
X9 a_343_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.127 ps=1.04 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
X0 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
X0 VPWR a_212_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_297_47# a_27_413# a_212_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_212_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.229 ps=1.75 w=1 l=0.15
X3 X a_212_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_212_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0767 ps=0.785 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VPWR B a_212_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.229 pd=1.75 as=0.0609 ps=0.71 w=0.42 l=0.15
X7 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND a_212_413# X VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 a_467_297# B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X1 a_287_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 VPWR A2 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X3 a_923_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.112 ps=0.995 w=0.65 l=0.15
X4 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.127 ps=1.04 w=0.65 l=0.15
X5 a_28_297# B1 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.185 ps=1.87 w=0.65 l=0.15
X7 a_28_297# C1 a_287_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X8 Y A1 a_923_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND A2 a_684_47# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.179 ps=1.2 w=0.65 l=0.15
X10 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X11 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.106 ps=0.975 w=0.65 l=0.15
X12 Y D1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 a_467_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=2.67 as=0.16 ps=1.32 w=1 l=0.15
X14 VGND D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X15 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.127 ps=1.04 w=0.65 l=0.15
X16 VPWR A1 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X17 a_115_297# C1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X18 a_467_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 a_684_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.2 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 VPWR a_82_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X1 a_646_47# B2 a_82_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_574_369# a_313_47# a_82_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0976 pd=0.945 as=0.166 ps=1.8 w=0.64 l=0.15
X3 a_574_369# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4 VGND a_82_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.09 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR B2 a_574_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0976 ps=0.945 w=0.64 l=0.15
X6 X a_82_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X7 X a_82_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X8 a_313_47# A2_N a_313_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.0672 ps=0.85 w=0.64 l=0.15
X9 a_313_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.12 ps=1.09 w=0.42 l=0.15
X10 a_313_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.186 ps=1.43 w=0.64 l=0.15
X11 VGND A2_N a_313_47# VNB sky130_fd_pr__nfet_01v8 ad=0.142 pd=1.1 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_82_21# a_313_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.142 ps=1.1 w=0.42 l=0.15
X13 VGND B1 a_646_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
X0 Y a_251_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y a_251_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X5 VGND a_251_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 VPWR B_N a_251_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X8 VGND B_N a_251_21# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_27_297# a_251_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X3 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X17 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X30 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X31 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 a_397_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR B1_N a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X2 Y A2 a_397_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 VGND A2 a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VGND A1 a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_28_297# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X6 Y a_28_297# a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VPWR a_28_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 a_397_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X9 a_229_47# a_28_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 Y a_28_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X11 a_229_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_229_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VPWR A1 a_397_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 a_298_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VGND A1 a_497_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3 a_664_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND A2 a_497_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 a_298_47# B1 a_497_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.176 ps=1.84 w=0.65 l=0.15
X7 a_497_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 Y D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.224 ps=1.99 w=0.65 l=0.15
X9 a_497_47# B1 a_298_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 Y A2 a_664_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.295 ps=2.59 w=1 l=0.15
X12 a_27_47# C1 a_298_47# VNB sky130_fd_pr__nfet_01v8 ad=0.192 pd=1.89 as=0.091 ps=0.93 w=0.65 l=0.15
X13 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X15 a_27_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X16 a_497_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.091 ps=0.93 w=0.65 l=0.15
X17 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X18 VPWR A1 a_664_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 a_664_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 VPWR A1 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 a_806_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.101 ps=0.96 w=0.65 l=0.15
X3 a_110_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VPWR A1 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X10 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_47# B1 a_1314_47# VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=2.09 as=0.104 ps=0.97 w=0.65 l=0.15
X12 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X14 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X17 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.0943 ps=0.94 w=0.65 l=0.15
X19 Y C1 a_978_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 Y C1 a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X22 a_27_47# B1 a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X23 a_110_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 a_806_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.675 pd=3.35 as=0.135 ps=1.27 w=1 l=0.15
X26 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.091 ps=0.93 w=0.65 l=0.15
X27 a_978_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.091 ps=0.93 w=0.65 l=0.15
X28 a_1314_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X31 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 a_27_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_27_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=1.77 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X9 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.385 ps=1.77 w=1 l=0.15
X14 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X21 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X24 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 a_445_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_445_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X28 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X31 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_47# C a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y A a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.107 ps=0.98 w=0.65 l=0.15
X5 a_277_47# B a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.219 pd=1.33 as=0.101 ps=0.96 w=0.65 l=0.15
X1 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.219 ps=1.33 w=0.65 l=0.15
X2 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.105 ps=1.21 w=1 l=0.15
X3 a_333_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.245 pd=1.49 as=0.305 ps=1.61 w=1 l=0.15
X4 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.106 ps=0.975 w=0.65 l=0.15
X6 VPWR A1 a_461_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X7 a_109_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X8 a_461_297# A2 a_333_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.245 ps=1.49 w=1 l=0.15
X9 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 a_316_297# C1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.172 ps=1.35 w=1 l=0.15
X1 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.03 as=0.481 ps=2.78 w=0.65 l=0.15
X2 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.02 as=0.125 ps=1.03 w=0.65 l=0.15
X3 a_420_297# B1 a_316_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=1.58 as=0.185 ps=1.37 w=1 l=0.15
X4 VPWR A1 a_420_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.29 ps=1.58 w=1 l=0.15
X5 VGND A2 a_568_47# VNB sky130_fd_pr__nfet_01v8 ad=0.192 pd=1.89 as=0.0845 ps=0.91 w=0.65 l=0.15
X6 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.192 pd=1.24 as=0.12 ps=1.02 w=0.65 l=0.15
X7 a_420_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.138 ps=1.27 w=1 l=0.15
X8 a_217_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.755 ps=3.51 w=1 l=0.15
X9 a_568_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0845 pd=0.91 as=0.192 ps=1.24 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
X0 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
X0 Y A a_150_67# VNB sky130_fd_pr__nfet_01v8 ad=0.157 pd=1.67 as=0.066 ps=0.79 w=0.55 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=2.78 as=0.14 ps=1.28 w=1 l=0.25
X2 a_150_67# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.79 as=0.157 ps=1.67 w=0.55 l=0.15
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
.ends

.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 Y A1 a_478_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.377 ps=1.75 w=1 l=0.15
X2 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.305 ps=1.61 w=1 l=0.15
X3 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.335 ps=1.67 w=1 l=0.15
X4 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.138 ps=1.27 w=1 l=0.15
X5 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.377 pd=1.75 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_478_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_478_47# A2 a_730_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VGND A3 a_730_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12 ps=1.02 w=0.65 l=0.15
X10 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_730_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.02 as=0.205 ps=1.93 w=0.65 l=0.15
X16 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.15 ps=1.3 w=1 l=0.15
X18 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X19 a_730_47# A2 a_478_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
.ends

.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 a_301_47# B2 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VGND A2 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.123 ps=1.03 w=0.65 l=0.15
X2 a_383_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.39 ps=1.78 w=1 l=0.15
X3 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=1.78 as=0.135 ps=1.27 w=1 l=0.15
X4 a_301_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 X a_81_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_81_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X8 VPWR A1 a_579_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X9 a_81_21# B1 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_579_297# A2 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X11 a_81_21# B2 a_383_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.105 ps=1.21 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
X0 Y A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_641_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=1.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_109_297# B1 a_641_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X5 a_277_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR A3 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_27_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.17 w=0.65 l=0.15
X11 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X12 a_641_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13 a_277_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0975 ps=0.95 w=0.65 l=0.15
X15 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 Y C1 a_641_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=1.52 w=1 l=0.15
X18 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X19 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt top VGND VPWR angle_in[0] angle_in[10] angle_in[11] angle_in[12] angle_in[13]
+ angle_in[14] angle_in[15] angle_in[1] angle_in[2] angle_in[3] angle_in[4] angle_in[5]
+ angle_in[6] angle_in[7] angle_in[8] angle_in[9] clk currA_in[0] currA_in[10] currA_in[11]
+ currA_in[12] currA_in[13] currA_in[14] currA_in[15] currA_in[1] currA_in[2] currA_in[3]
+ currA_in[4] currA_in[5] currA_in[6] currA_in[7] currA_in[8] currA_in[9] currB_in[0]
+ currB_in[10] currB_in[11] currB_in[12] currB_in[13] currB_in[14] currB_in[15] currB_in[1]
+ currB_in[2] currB_in[3] currB_in[4] currB_in[5] currB_in[6] currB_in[7] currB_in[8]
+ currB_in[9] currC_in[0] currC_in[10] currC_in[11] currC_in[12] currC_in[13] currC_in[14]
+ currC_in[15] currC_in[1] currC_in[2] currC_in[3] currC_in[4] currC_in[5] currC_in[6]
+ currC_in[7] currC_in[8] currC_in[9] currT_in[0] currT_in[10] currT_in[11] currT_in[12]
+ currT_in[13] currT_in[14] currT_in[15] currT_in[1] currT_in[2] currT_in[3] currT_in[4]
+ currT_in[5] currT_in[6] currT_in[7] currT_in[8] currT_in[9] periodTop[0] periodTop[10]
+ periodTop[11] periodTop[12] periodTop[13] periodTop[14] periodTop[15] periodTop[1]
+ periodTop[2] periodTop[3] periodTop[4] periodTop[5] periodTop[6] periodTop[7] periodTop[8]
+ periodTop[9] pid_d_addr[0] pid_d_addr[10] pid_d_addr[11] pid_d_addr[12] pid_d_addr[13]
+ pid_d_addr[14] pid_d_addr[15] pid_d_addr[1] pid_d_addr[2] pid_d_addr[3] pid_d_addr[4]
+ pid_d_addr[5] pid_d_addr[6] pid_d_addr[7] pid_d_addr[8] pid_d_addr[9] pid_d_data[0]
+ pid_d_data[10] pid_d_data[11] pid_d_data[12] pid_d_data[13] pid_d_data[14] pid_d_data[15]
+ pid_d_data[1] pid_d_data[2] pid_d_data[3] pid_d_data[4] pid_d_data[5] pid_d_data[6]
+ pid_d_data[7] pid_d_data[8] pid_d_data[9] pid_d_wen pid_q_addr[0] pid_q_addr[10]
+ pid_q_addr[11] pid_q_addr[12] pid_q_addr[13] pid_q_addr[14] pid_q_addr[15] pid_q_addr[1]
+ pid_q_addr[2] pid_q_addr[3] pid_q_addr[4] pid_q_addr[5] pid_q_addr[6] pid_q_addr[7]
+ pid_q_addr[8] pid_q_addr[9] pid_q_data[0] pid_q_data[10] pid_q_data[11] pid_q_data[12]
+ pid_q_data[13] pid_q_data[14] pid_q_data[15] pid_q_data[1] pid_q_data[2] pid_q_data[3]
+ pid_q_data[4] pid_q_data[5] pid_q_data[6] pid_q_data[7] pid_q_data[8] pid_q_data[9]
+ pid_q_wen pwmA_out pwmB_out pwmC_out ready rstb valid
XFILLER_0_193_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18869_ _10709_ _10710_ VGND VGND VPWR VPWR _10711_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20900_ _00895_ _00914_ _00915_ VGND VGND VPWR VPWR _00916_ sky130_fd_sc_hd__a21o_1
X_21880_ _01780_ _01790_ _01886_ _01888_ VGND VGND VPWR VPWR _01889_ sky130_fd_sc_hd__a22o_1
X_20831_ _12548_ _12549_ _12550_ VGND VGND VPWR VPWR _00847_ sky130_fd_sc_hd__o21a_1
XFILLER_0_178_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23550_ _03322_ _03323_ _03324_ VGND VGND VPWR VPWR _03418_ sky130_fd_sc_hd__o21a_1
X_20762_ _12530_ net2485 VGND VGND VPWR VPWR _12533_ sky130_fd_sc_hd__nor2_1
Xmax_length5429 net5423 VGND VGND VPWR VPWR net5429 sky130_fd_sc_hd__buf_1
Xmax_length4706 net4707 VGND VGND VPWR VPWR net4706 sky130_fd_sc_hd__clkbuf_1
X_22501_ _02438_ _02501_ VGND VGND VPWR VPWR _02502_ sky130_fd_sc_hd__nand2_1
X_23481_ net4727 net4876 VGND VGND VPWR VPWR _03350_ sky130_fd_sc_hd__nand2_2
X_20693_ _12466_ _12467_ VGND VGND VPWR VPWR _12468_ sky130_fd_sc_hd__xor2_1
Xmax_length4728 net4729 VGND VGND VPWR VPWR net4728 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22432_ _02229_ _02300_ _02433_ VGND VGND VPWR VPWR _02434_ sky130_fd_sc_hd__or3_1
X_25220_ clknet_leaf_59_clk _00109_ net8693 VGND VGND VPWR VPWR svm0.vC\[8\] sky130_fd_sc_hd__dfrtp_1
Xwire709 net710 VGND VGND VPWR VPWR net709 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25151_ clknet_leaf_44_clk _00040_ net8781 VGND VGND VPWR VPWR pid_q.target\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_22363_ _02364_ _02365_ VGND VGND VPWR VPWR _02366_ sky130_fd_sc_hd__and2b_1
XFILLER_0_165_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24102_ net4980 net4484 VGND VGND VPWR VPWR _03964_ sky130_fd_sc_hd__nand2_2
X_21314_ _01325_ net758 VGND VGND VPWR VPWR _01329_ sky130_fd_sc_hd__nand2_1
X_25082_ _04826_ _04827_ net1994 VGND VGND VPWR VPWR _04828_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_103_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22294_ _02215_ _02216_ _02217_ VGND VGND VPWR VPWR _02298_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4005 _09376_ VGND VGND VPWR VPWR net4005 sky130_fd_sc_hd__clkbuf_1
X_24033_ _03894_ _03895_ VGND VGND VPWR VPWR _03896_ sky130_fd_sc_hd__xnor2_1
Xwire4027 _09223_ VGND VGND VPWR VPWR net4027 sky130_fd_sc_hd__buf_1
XFILLER_0_130_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21245_ _01258_ _01259_ VGND VGND VPWR VPWR _01260_ sky130_fd_sc_hd__xnor2_1
Xwire4038 _09054_ VGND VGND VPWR VPWR net4038 sky130_fd_sc_hd__buf_1
Xwire3304 _09093_ VGND VGND VPWR VPWR net3304 sky130_fd_sc_hd__clkbuf_1
Xwire4049 _08949_ VGND VGND VPWR VPWR net4049 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3315 net3316 VGND VGND VPWR VPWR net3315 sky130_fd_sc_hd__clkbuf_1
X_21176_ _01150_ _01151_ VGND VGND VPWR VPWR _01192_ sky130_fd_sc_hd__nand2_1
Xwire3337 net3338 VGND VGND VPWR VPWR net3337 sky130_fd_sc_hd__buf_1
Xwire2603 _08988_ VGND VGND VPWR VPWR net2603 sky130_fd_sc_hd__clkbuf_1
Xwire3348 _08914_ VGND VGND VPWR VPWR net3348 sky130_fd_sc_hd__buf_1
Xwire2614 net2615 VGND VGND VPWR VPWR net2614 sky130_fd_sc_hd__clkbuf_1
Xwire3359 _08909_ VGND VGND VPWR VPWR net3359 sky130_fd_sc_hd__buf_1
X_20127_ net1055 _11953_ VGND VGND VPWR VPWR _11955_ sky130_fd_sc_hd__and2_1
Xwire2625 net2626 VGND VGND VPWR VPWR net2625 sky130_fd_sc_hd__buf_1
Xwire2636 net2637 VGND VGND VPWR VPWR net2636 sky130_fd_sc_hd__buf_1
Xwire1902 net1903 VGND VGND VPWR VPWR net1902 sky130_fd_sc_hd__buf_1
Xwire2647 _07780_ VGND VGND VPWR VPWR net2647 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1913 net1914 VGND VGND VPWR VPWR net1913 sky130_fd_sc_hd__clkbuf_1
Xwire2658 _07724_ VGND VGND VPWR VPWR net2658 sky130_fd_sc_hd__clkbuf_1
Xwire1924 net1925 VGND VGND VPWR VPWR net1924 sky130_fd_sc_hd__clkbuf_1
Xwire2669 _07713_ VGND VGND VPWR VPWR net2669 sky130_fd_sc_hd__clkbuf_1
Xwire1935 net1936 VGND VGND VPWR VPWR net1935 sky130_fd_sc_hd__clkbuf_1
X_24935_ _04717_ VGND VGND VPWR VPWR _00752_ sky130_fd_sc_hd__clkbuf_1
X_20058_ net6134 _11883_ _11886_ VGND VGND VPWR VPWR _11887_ sky130_fd_sc_hd__a21oi_2
Xwire1946 _05487_ VGND VGND VPWR VPWR net1946 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1957 _05064_ VGND VGND VPWR VPWR net1957 sky130_fd_sc_hd__clkbuf_2
Xmax_length8011 pid_q.target\[5\] VGND VGND VPWR VPWR net8011 sky130_fd_sc_hd__clkbuf_1
Xwire1968 _04932_ VGND VGND VPWR VPWR net1968 sky130_fd_sc_hd__buf_1
XFILLER_0_99_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1979 net1980 VGND VGND VPWR VPWR net1979 sky130_fd_sc_hd__buf_1
X_24866_ _04667_ net4724 net1997 VGND VGND VPWR VPWR _04669_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12880_ net1336 _05100_ VGND VGND VPWR VPWR _05153_ sky130_fd_sc_hd__nor2_1
X_23817_ net4542 net4991 VGND VGND VPWR VPWR _03682_ sky130_fd_sc_hd__nand2_1
XFILLER_0_185_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24797_ _04619_ _04620_ _04618_ VGND VGND VPWR VPWR _04622_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14550_ net5250 _06710_ _06712_ VGND VGND VPWR VPWR _06728_ sky130_fd_sc_hd__o21ai_1
X_23748_ _03588_ _03613_ VGND VGND VPWR VPWR _03614_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13501_ net504 _05773_ VGND VGND VPWR VPWR _05774_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14481_ net7361 net5305 _06663_ VGND VGND VPWR VPWR _06666_ sky130_fd_sc_hd__a21oi_1
X_23679_ _03455_ _03457_ _03458_ VGND VGND VPWR VPWR _03546_ sky130_fd_sc_hd__a21o_1
Xmax_length5952 net5948 VGND VGND VPWR VPWR net5952 sky130_fd_sc_hd__buf_1
XFILLER_0_82_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16220_ _08193_ _08198_ _08284_ VGND VGND VPWR VPWR _08285_ sky130_fd_sc_hd__o21a_1
X_13432_ net7834 net1587 _05607_ _05610_ VGND VGND VPWR VPWR _05705_ sky130_fd_sc_hd__a22o_1
X_25418_ clknet_leaf_91_clk _00301_ net8428 VGND VGND VPWR VPWR matmul0.cos\[5\] sky130_fd_sc_hd__dfrtp_1
Xmax_length5985 pid_d.curr_int\[1\] VGND VGND VPWR VPWR net5985 sky130_fd_sc_hd__buf_1
XFILLER_0_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16151_ net2802 _08216_ VGND VGND VPWR VPWR _08217_ sky130_fd_sc_hd__nor2_1
X_13363_ net732 _05550_ _05551_ VGND VGND VPWR VPWR _05636_ sky130_fd_sc_hd__o21ba_1
X_25349_ clknet_leaf_82_clk _00232_ net8503 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15102_ _07172_ _07173_ _07175_ VGND VGND VPWR VPWR _07176_ sky130_fd_sc_hd__o21ai_1
Xfanout5156 pid_q.mult0.b\[0\] VGND VGND VPWR VPWR net5156 sky130_fd_sc_hd__buf_1
X_16082_ _08147_ _08148_ VGND VGND VPWR VPWR _08149_ sky130_fd_sc_hd__xnor2_1
X_13294_ net732 _05552_ VGND VGND VPWR VPWR _05567_ sky130_fd_sc_hd__xor2_1
Xwire5240 net5241 VGND VGND VPWR VPWR net5240 sky130_fd_sc_hd__clkbuf_1
Xwire5251 net5252 VGND VGND VPWR VPWR net5251 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19910_ _11667_ _11739_ _11741_ VGND VGND VPWR VPWR _11742_ sky130_fd_sc_hd__o21ai_1
X_15033_ net4181 net4179 VGND VGND VPWR VPWR _07107_ sky130_fd_sc_hd__nor2_1
Xwire5262 net5263 VGND VGND VPWR VPWR net5262 sky130_fd_sc_hd__clkbuf_2
Xwire5273 net5274 VGND VGND VPWR VPWR net5273 sky130_fd_sc_hd__buf_1
Xwire5284 net5285 VGND VGND VPWR VPWR net5284 sky130_fd_sc_hd__buf_1
XFILLER_0_20_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4550 pid_q.mult0.a\[12\] VGND VGND VPWR VPWR net4550 sky130_fd_sc_hd__buf_1
Xwire5295 net5296 VGND VGND VPWR VPWR net5295 sky130_fd_sc_hd__clkbuf_1
Xwire4561 net4562 VGND VGND VPWR VPWR net4561 sky130_fd_sc_hd__buf_1
X_19841_ _11631_ _11653_ _11673_ VGND VGND VPWR VPWR _11674_ sky130_fd_sc_hd__a21oi_2
Xwire4572 net4573 VGND VGND VPWR VPWR net4572 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4583 net4584 VGND VGND VPWR VPWR net4583 sky130_fd_sc_hd__clkbuf_1
Xwire3871 net3872 VGND VGND VPWR VPWR net3871 sky130_fd_sc_hd__clkbuf_1
X_16984_ _08824_ _08926_ net4051 net6019 VGND VGND VPWR VPWR _08946_ sky130_fd_sc_hd__a22o_1
X_19772_ _11534_ net1057 _11532_ VGND VGND VPWR VPWR _11607_ sky130_fd_sc_hd__a21o_1
Xwire3882 _10983_ VGND VGND VPWR VPWR net3882 sky130_fd_sc_hd__clkbuf_1
Xwire3893 net3894 VGND VGND VPWR VPWR net3893 sky130_fd_sc_hd__buf_1
XFILLER_0_155_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15935_ _07911_ _07912_ VGND VGND VPWR VPWR _08004_ sky130_fd_sc_hd__nor2_1
X_18723_ net9016 net1203 _10568_ net1771 VGND VGND VPWR VPWR _00444_ sky130_fd_sc_hd__a22o_1
X_18654_ _10453_ _10499_ _10461_ VGND VGND VPWR VPWR _10501_ sky130_fd_sc_hd__or3_1
X_15866_ net3550 net3434 VGND VGND VPWR VPWR _07935_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17605_ svm0.tB\[9\] VGND VGND VPWR VPWR _09486_ sky130_fd_sc_hd__inv_2
X_14817_ net9026 net2877 net2854 _06925_ VGND VGND VPWR VPWR _00180_ sky130_fd_sc_hd__o22a_1
X_18585_ net3225 _10432_ VGND VGND VPWR VPWR _10433_ sky130_fd_sc_hd__xnor2_1
X_15797_ net3546 _07866_ VGND VGND VPWR VPWR _07867_ sky130_fd_sc_hd__nor2_1
XFILLER_0_175_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17536_ svm0.counter\[15\] _09268_ _09417_ VGND VGND VPWR VPWR _09419_ sky130_fd_sc_hd__or3_1
XFILLER_0_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14748_ net7454 _06880_ net2857 VGND VGND VPWR VPWR _06881_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17467_ _09287_ _09354_ _09359_ VGND VGND VPWR VPWR _09360_ sky130_fd_sc_hd__o21a_1
XFILLER_0_188_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14679_ net7433 net2869 net2263 net2864 VGND VGND VPWR VPWR _00138_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19206_ _11028_ _11041_ _11042_ VGND VGND VPWR VPWR _11043_ sky130_fd_sc_hd__o21ba_1
X_16418_ net723 _08479_ VGND VGND VPWR VPWR _08480_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_13_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17398_ svm0.delta\[7\] _09300_ VGND VGND VPWR VPWR _09304_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19137_ _10971_ net3185 VGND VGND VPWR VPWR _10974_ sky130_fd_sc_hd__xor2_2
X_16349_ net1079 _08411_ VGND VGND VPWR VPWR _08412_ sky130_fd_sc_hd__xnor2_1
Xfanout7092 net7093 VGND VGND VPWR VPWR net7092 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_120_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19068_ _10891_ _10892_ _10897_ net1758 _10904_ VGND VGND VPWR VPWR _10905_ sky130_fd_sc_hd__o311a_1
XFILLER_0_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18019_ net7052 net7107 VGND VGND VPWR VPWR _09870_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_11_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_196_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21030_ _01036_ _01041_ _01045_ VGND VGND VPWR VPWR _01046_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1209 _10272_ VGND VGND VPWR VPWR net1209 sky130_fd_sc_hd__clkbuf_1
X_22981_ _02858_ VGND VGND VPWR VPWR _00657_ sky130_fd_sc_hd__clkbuf_1
X_24720_ pid_q.curr_error\[3\] net1368 net1365 net1640 VGND VGND VPWR VPWR _00700_
+ sky130_fd_sc_hd__a22o_1
X_21932_ _01836_ _01841_ _01831_ VGND VGND VPWR VPWR _01940_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_69_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24651_ _04330_ _04459_ _04501_ _04383_ net195 VGND VGND VPWR VPWR _04506_ sky130_fd_sc_hd__o221a_1
X_21863_ net5812 _01868_ _01870_ _01866_ _01871_ VGND VGND VPWR VPWR _01872_ sky130_fd_sc_hd__o221a_1
XFILLER_0_179_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23602_ _03469_ _03318_ VGND VGND VPWR VPWR _03470_ sky130_fd_sc_hd__or2b_1
XFILLER_0_49_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20814_ _00826_ _00829_ VGND VGND VPWR VPWR _00830_ sky130_fd_sc_hd__xnor2_2
X_24582_ _04284_ _04437_ VGND VGND VPWR VPWR _04438_ sky130_fd_sc_hd__xnor2_2
X_21794_ _01742_ _01803_ VGND VGND VPWR VPWR _01804_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_166_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8805 net8803 VGND VGND VPWR VPWR net8805 sky130_fd_sc_hd__dlymetal6s2s_1
X_23533_ net4540 net5079 VGND VGND VPWR VPWR _03401_ sky130_fd_sc_hd__nand2_1
Xwire8816 net8817 VGND VGND VPWR VPWR net8816 sky130_fd_sc_hd__clkbuf_1
X_20745_ net5953 net5424 VGND VGND VPWR VPWR _12516_ sky130_fd_sc_hd__nand2_1
Xwire8827 net8828 VGND VGND VPWR VPWR net8827 sky130_fd_sc_hd__clkbuf_1
Xwire8838 net8839 VGND VGND VPWR VPWR net8838 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8849 net8850 VGND VGND VPWR VPWR net8849 sky130_fd_sc_hd__clkbuf_1
X_23464_ _03329_ _03332_ VGND VGND VPWR VPWR _03333_ sky130_fd_sc_hd__xnor2_1
Xwire506 net507 VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__clkbuf_1
X_20676_ net1394 _12429_ _12443_ VGND VGND VPWR VPWR _12452_ sky130_fd_sc_hd__or3_1
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4558 net4562 VGND VGND VPWR VPWR net4558 sky130_fd_sc_hd__buf_1
Xwire517 net518 VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__buf_1
Xmax_length4569 pid_q.mult0.a\[11\] VGND VGND VPWR VPWR net4569 sky130_fd_sc_hd__buf_1
Xwire528 _08720_ VGND VGND VPWR VPWR net528 sky130_fd_sc_hd__buf_1
XFILLER_0_190_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25203_ clknet_leaf_57_clk _00092_ net8715 VGND VGND VPWR VPWR matmul0.b_in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_163_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22415_ _02367_ _02345_ _02416_ VGND VGND VPWR VPWR _02417_ sky130_fd_sc_hd__o21ai_2
Xwire539 net540 VGND VGND VPWR VPWR net539 sky130_fd_sc_hd__clkbuf_1
X_23395_ net5099 net4563 VGND VGND VPWR VPWR _03265_ sky130_fd_sc_hd__nand2_2
XFILLER_0_33_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length3868 _11274_ VGND VGND VPWR VPWR net3868 sky130_fd_sc_hd__buf_1
XFILLER_0_6_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3879 _10996_ VGND VGND VPWR VPWR net3879 sky130_fd_sc_hd__buf_1
X_25134_ clknet_leaf_52_clk _00023_ net8803 VGND VGND VPWR VPWR svm0.tC\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22346_ net5720 net5745 VGND VGND VPWR VPWR _02349_ sky130_fd_sc_hd__xor2_1
XFILLER_0_61_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22277_ _02233_ net1033 _02280_ VGND VGND VPWR VPWR _02281_ sky130_fd_sc_hd__o21ai_2
X_25065_ net1627 _04812_ net2148 VGND VGND VPWR VPWR _04813_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3101 net3102 VGND VGND VPWR VPWR net3101 sky130_fd_sc_hd__clkbuf_1
X_24016_ net4987 net4500 VGND VGND VPWR VPWR _03879_ sky130_fd_sc_hd__nand2_1
X_21228_ pid_d.prev_error\[0\] net5973 VGND VGND VPWR VPWR _01244_ sky130_fd_sc_hd__xnor2_1
Xwire3112 net3113 VGND VGND VPWR VPWR net3112 sky130_fd_sc_hd__clkbuf_1
Xhold170 pid_q.prev_error\[7\] VGND VGND VPWR VPWR net9123 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3123 _12500_ VGND VGND VPWR VPWR net3123 sky130_fd_sc_hd__clkbuf_2
Xhold181 pid_d.prev_int\[15\] VGND VGND VPWR VPWR net9134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 pid_q.prev_error\[6\] VGND VGND VPWR VPWR net9145 sky130_fd_sc_hd__dlygate4sd3_1
Xwire2400 net2401 VGND VGND VPWR VPWR net2400 sky130_fd_sc_hd__clkbuf_1
Xwire2411 _03786_ VGND VGND VPWR VPWR net2411 sky130_fd_sc_hd__buf_1
Xwire3156 _11349_ VGND VGND VPWR VPWR net3156 sky130_fd_sc_hd__clkbuf_1
Xwire2422 net2423 VGND VGND VPWR VPWR net2422 sky130_fd_sc_hd__clkbuf_1
X_21159_ net5625 net5611 _01174_ net5916 net5641 VGND VGND VPWR VPWR _01175_ sky130_fd_sc_hd__a32o_1
Xwire3167 _11132_ VGND VGND VPWR VPWR net3167 sky130_fd_sc_hd__clkbuf_2
Xwire2433 _02869_ VGND VGND VPWR VPWR net2433 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3178 net3179 VGND VGND VPWR VPWR net3178 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2444 net2445 VGND VGND VPWR VPWR net2444 sky130_fd_sc_hd__clkbuf_1
Xwire3189 _10942_ VGND VGND VPWR VPWR net3189 sky130_fd_sc_hd__buf_1
Xwire1710 net1711 VGND VGND VPWR VPWR net1710 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2455 _02603_ VGND VGND VPWR VPWR net2455 sky130_fd_sc_hd__clkbuf_1
Xwire2466 net2467 VGND VGND VPWR VPWR net2466 sky130_fd_sc_hd__buf_1
Xwire1721 _01597_ VGND VGND VPWR VPWR net1721 sky130_fd_sc_hd__buf_1
X_13981_ _06244_ net1305 VGND VGND VPWR VPWR _06246_ sky130_fd_sc_hd__or2_1
Xwire2477 _01710_ VGND VGND VPWR VPWR net2477 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1732 net1733 VGND VGND VPWR VPWR net1732 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2488 net2489 VGND VGND VPWR VPWR net2488 sky130_fd_sc_hd__buf_1
Xwire1743 net1744 VGND VGND VPWR VPWR net1743 sky130_fd_sc_hd__clkbuf_1
Xwire1754 net1755 VGND VGND VPWR VPWR net1754 sky130_fd_sc_hd__clkbuf_1
Xwire2499 _11763_ VGND VGND VPWR VPWR net2499 sky130_fd_sc_hd__clkbuf_1
X_15720_ _07785_ _07790_ VGND VGND VPWR VPWR _07791_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24918_ net8867 net138 VGND VGND VPWR VPWR _04706_ sky130_fd_sc_hd__and2b_1
X_12932_ net1333 _05140_ VGND VGND VPWR VPWR _05205_ sky130_fd_sc_hd__nand2_1
Xwire1765 _10366_ VGND VGND VPWR VPWR net1765 sky130_fd_sc_hd__clkbuf_1
Xwire1776 _10120_ VGND VGND VPWR VPWR net1776 sky130_fd_sc_hd__buf_1
X_25898_ clknet_leaf_16_clk _00771_ net8627 VGND VGND VPWR VPWR pid_q.kp\[10\] sky130_fd_sc_hd__dfrtp_1
Xwire1798 _09194_ VGND VGND VPWR VPWR net1798 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_87_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15651_ net4079 net4077 VGND VGND VPWR VPWR _07723_ sky130_fd_sc_hd__nor2_1
X_24849_ _04534_ _04657_ net4821 _04642_ VGND VGND VPWR VPWR _00726_ sky130_fd_sc_hd__a2bb2o_1
X_12863_ net1957 _05111_ VGND VGND VPWR VPWR _05136_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_157_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14602_ net7209 net5194 VGND VGND VPWR VPWR _06775_ sky130_fd_sc_hd__nor2_1
X_18370_ net6858 _10169_ _10219_ net3299 _10220_ VGND VGND VPWR VPWR _10221_ sky130_fd_sc_hd__a221o_1
X_15582_ net4160 net4156 net4098 net4096 VGND VGND VPWR VPWR _07654_ sky130_fd_sc_hd__o22a_1
X_12794_ _05049_ net1144 VGND VGND VPWR VPWR _05067_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length7184 matmul0.b\[8\] VGND VGND VPWR VPWR net7184 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17321_ net4022 _09209_ _09231_ _09232_ VGND VGND VPWR VPWR _09235_ sky130_fd_sc_hd__and4_1
X_14533_ net2388 _06703_ net726 VGND VGND VPWR VPWR _06712_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6494 net6495 VGND VGND VPWR VPWR net6494 sky130_fd_sc_hd__buf_1
XFILLER_0_139_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17252_ _09185_ net218 _09190_ net9099 VGND VGND VPWR VPWR _00350_ sky130_fd_sc_hd__a22o_1
XFILLER_0_166_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14464_ net892 VGND VGND VPWR VPWR _06652_ sky130_fd_sc_hd__buf_1
XFILLER_0_37_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16203_ _08177_ _08262_ net1512 VGND VGND VPWR VPWR _08268_ sky130_fd_sc_hd__a21bo_1
X_13415_ net7900 net1327 VGND VGND VPWR VPWR _05688_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17183_ _09122_ _09123_ net1076 VGND VGND VPWR VPWR _09134_ sky130_fd_sc_hd__o21ai_1
X_14395_ _06599_ VGND VGND VPWR VPWR _00084_ sky130_fd_sc_hd__clkbuf_1
X_16134_ _08191_ _08199_ VGND VGND VPWR VPWR _08200_ sky130_fd_sc_hd__xnor2_1
X_13346_ net3682 VGND VGND VPWR VPWR _05619_ sky130_fd_sc_hd__buf_1
XFILLER_0_3_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16065_ net2205 _08049_ VGND VGND VPWR VPWR _08132_ sky130_fd_sc_hd__or2_1
X_13277_ _05547_ _05548_ net846 VGND VGND VPWR VPWR _05550_ sky130_fd_sc_hd__and3_1
Xwire5070 net5071 VGND VGND VPWR VPWR net5070 sky130_fd_sc_hd__buf_1
Xwire5081 net5082 VGND VGND VPWR VPWR net5081 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15016_ net4143 net4140 net4122 net4117 VGND VGND VPWR VPWR _07090_ sky130_fd_sc_hd__o22a_1
Xwire5092 net5093 VGND VGND VPWR VPWR net5092 sky130_fd_sc_hd__clkbuf_1
Xwire4380 net4379 VGND VGND VPWR VPWR net4380 sky130_fd_sc_hd__buf_1
Xwire4391 pid_d.prev_int\[12\] VGND VGND VPWR VPWR net4391 sky130_fd_sc_hd__buf_1
X_19824_ net6032 net1056 VGND VGND VPWR VPWR _11658_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3690 net3691 VGND VGND VPWR VPWR net3690 sky130_fd_sc_hd__clkbuf_1
X_19755_ _11588_ net3129 net6067 VGND VGND VPWR VPWR _11590_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16967_ net6123 net6082 net6501 VGND VGND VPWR VPWR _08930_ sky130_fd_sc_hd__mux2_1
X_18706_ _10520_ _10551_ VGND VGND VPWR VPWR _10552_ sky130_fd_sc_hd__xnor2_2
X_15918_ net826 _07986_ VGND VGND VPWR VPWR _07987_ sky130_fd_sc_hd__xnor2_1
X_19686_ _11520_ _11521_ VGND VGND VPWR VPWR _11522_ sky130_fd_sc_hd__nor2_2
X_16898_ cordic0.slte0.opB\[11\] VGND VGND VPWR VPWR _08862_ sky130_fd_sc_hd__inv_2
X_15849_ _07914_ _07918_ VGND VGND VPWR VPWR _07919_ sky130_fd_sc_hd__nor2_1
X_18637_ net1431 _10483_ VGND VGND VPWR VPWR _10484_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_182_Left_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18568_ _10284_ net2540 VGND VGND VPWR VPWR _10416_ sky130_fd_sc_hd__or2b_1
XFILLER_0_24_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17519_ _09319_ _09400_ net6697 VGND VGND VPWR VPWR _09404_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_19_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18499_ net6774 net2540 VGND VGND VPWR VPWR _10348_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20530_ net7088 net7042 net7074 net7010 net6489 net6514 VGND VGND VPWR VPWR _12316_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_90_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20461_ _12250_ cordic0.slte0.opA\[15\] _12252_ VGND VGND VPWR VPWR _12253_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22200_ _02141_ _02143_ _02139_ VGND VGND VPWR VPWR _02205_ sky130_fd_sc_hd__o21ba_1
X_23180_ net5115 net4737 VGND VGND VPWR VPWR _03050_ sky130_fd_sc_hd__nand2_1
XFILLER_0_171_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20392_ _12188_ _12189_ _12190_ net9188 VGND VGND VPWR VPWR _00491_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22131_ net3779 _02136_ net5764 net5389 VGND VGND VPWR VPWR _02137_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_191_Left_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22062_ _02067_ _02068_ VGND VGND VPWR VPWR _02069_ sky130_fd_sc_hd__or2b_1
XFILLER_0_100_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21013_ net1051 _01028_ VGND VGND VPWR VPWR _01029_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_26_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1006 _05116_ VGND VGND VPWR VPWR net1006 sky130_fd_sc_hd__buf_1
Xwire1017 _03768_ VGND VGND VPWR VPWR net1017 sky130_fd_sc_hd__buf_1
X_25821_ clknet_leaf_31_clk _00694_ net8686 VGND VGND VPWR VPWR pid_q.prev_error\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1028 net1029 VGND VGND VPWR VPWR net1028 sky130_fd_sc_hd__buf_1
Xwire1039 net1040 VGND VGND VPWR VPWR net1039 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25752_ clknet_leaf_13_clk _00625_ net8604 VGND VGND VPWR VPWR pid_d.kp\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22964_ matmul0.beta_pass\[1\] net3383 net6570 VGND VGND VPWR VPWR _02850_ sky130_fd_sc_hd__mux2_1
X_24703_ net4310 net3269 VGND VGND VPWR VPWR _04540_ sky130_fd_sc_hd__nor2_2
X_21915_ net599 _01922_ VGND VGND VPWR VPWR _01923_ sky130_fd_sc_hd__nand2_1
X_25683_ clknet_leaf_0_clk _00556_ net8409 VGND VGND VPWR VPWR pid_d.curr_error\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_22895_ net5354 _02785_ _02788_ VGND VGND VPWR VPWR _02789_ sky130_fd_sc_hd__mux2_1
X_24634_ _04350_ _04428_ _04488_ net4919 VGND VGND VPWR VPWR _04489_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21846_ net2474 _01854_ VGND VGND VPWR VPWR _01855_ sky130_fd_sc_hd__xor2_1
Xfanout8518 net8530 VGND VGND VPWR VPWR net8518 sky130_fd_sc_hd__buf_1
XFILLER_0_66_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24565_ net4794 _04343_ _04345_ _04418_ _04420_ VGND VGND VPWR VPWR _04421_ sky130_fd_sc_hd__o311a_1
XFILLER_0_38_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21777_ _01690_ _01691_ _01786_ VGND VGND VPWR VPWR _01787_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8613 net8614 VGND VGND VPWR VPWR net8613 sky130_fd_sc_hd__clkbuf_1
Xwire8624 net8625 VGND VGND VPWR VPWR net8624 sky130_fd_sc_hd__buf_1
Xmax_length5056 net5043 VGND VGND VPWR VPWR net5056 sky130_fd_sc_hd__clkbuf_1
X_23516_ pid_q.prev_error\[1\] net5168 VGND VGND VPWR VPWR _03385_ sky130_fd_sc_hd__xnor2_1
Xwire8635 net8636 VGND VGND VPWR VPWR net8635 sky130_fd_sc_hd__clkbuf_1
Xwire7901 net7902 VGND VGND VPWR VPWR net7901 sky130_fd_sc_hd__buf_1
X_20728_ net4390 net4346 net4324 net8906 VGND VGND VPWR VPWR _12499_ sky130_fd_sc_hd__o31a_1
Xwire8646 net8645 VGND VGND VPWR VPWR net8646 sky130_fd_sc_hd__buf_1
X_24496_ _04347_ _04352_ VGND VGND VPWR VPWR _04353_ sky130_fd_sc_hd__xnor2_2
Xwire7912 net7913 VGND VGND VPWR VPWR net7912 sky130_fd_sc_hd__clkbuf_1
Xwire8657 net8653 VGND VGND VPWR VPWR net8657 sky130_fd_sc_hd__buf_1
XFILLER_0_80_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7923 net7925 VGND VGND VPWR VPWR net7923 sky130_fd_sc_hd__buf_1
Xwire303 net304 VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__clkbuf_2
Xwire314 net315 VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__clkbuf_1
Xwire325 net326 VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__buf_1
XFILLER_0_162_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_137_Right_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8679 net8677 VGND VGND VPWR VPWR net8679 sky130_fd_sc_hd__buf_1
XFILLER_0_108_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7945 net7946 VGND VGND VPWR VPWR net7945 sky130_fd_sc_hd__clkbuf_1
X_23447_ pid_q.curr_int\[1\] pid_q.prev_int\[1\] VGND VGND VPWR VPWR _03316_ sky130_fd_sc_hd__xor2_1
Xwire336 _02277_ VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_20_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7956 net7957 VGND VGND VPWR VPWR net7956 sky130_fd_sc_hd__clkbuf_1
Xmax_length4388 pid_d.state\[1\] VGND VGND VPWR VPWR net4388 sky130_fd_sc_hd__buf_1
Xwire347 net348 VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__buf_1
X_20659_ _12435_ _12436_ VGND VGND VPWR VPWR _12437_ sky130_fd_sc_hd__nor2_1
Xwire7967 net7968 VGND VGND VPWR VPWR net7967 sky130_fd_sc_hd__buf_1
XFILLER_0_34_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13200_ _05362_ _05363_ _05472_ VGND VGND VPWR VPWR _05473_ sky130_fd_sc_hd__a21o_1
XFILLER_0_34_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire358 _08161_ VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__clkbuf_1
Xmax_length3676 net3677 VGND VGND VPWR VPWR net3676 sky130_fd_sc_hd__buf_1
Xwire369 net370 VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7978 net7979 VGND VGND VPWR VPWR net7978 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7989 pid_q.target\[9\] VGND VGND VPWR VPWR net7989 sky130_fd_sc_hd__clkbuf_1
X_14180_ net7627 net1123 _06407_ net1120 net7647 VGND VGND VPWR VPWR _06440_ sky130_fd_sc_hd__a32o_1
XFILLER_0_61_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23378_ net4833 net4773 VGND VGND VPWR VPWR _03248_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3698 _04884_ VGND VGND VPWR VPWR net3698 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13131_ net683 net848 VGND VGND VPWR VPWR _05404_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25117_ net9236 net2393 net1993 pid_d.curr_int\[5\] VGND VGND VPWR VPWR _00798_ sky130_fd_sc_hd__a22o_1
X_22329_ _02330_ _02331_ VGND VGND VPWR VPWR _02332_ sky130_fd_sc_hd__or2b_1
XFILLER_0_60_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25048_ net7473 _04797_ _04798_ net7512 net329 VGND VGND VPWR VPWR _04799_ sky130_fd_sc_hd__a32o_1
X_13062_ _05284_ _05303_ VGND VGND VPWR VPWR _05335_ sky130_fd_sc_hd__nand2_1
X_17870_ _09720_ _09602_ VGND VGND VPWR VPWR _09721_ sky130_fd_sc_hd__xnor2_1
Xwire2230 net2231 VGND VGND VPWR VPWR net2230 sky130_fd_sc_hd__clkbuf_1
Xwire2252 net2253 VGND VGND VPWR VPWR net2252 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16821_ net9233 matmul0.cos\[13\] net3368 VGND VGND VPWR VPWR _08801_ sky130_fd_sc_hd__mux2_1
Xwire2274 net2275 VGND VGND VPWR VPWR net2274 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2285 net2286 VGND VGND VPWR VPWR net2285 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1540 net1541 VGND VGND VPWR VPWR net1540 sky130_fd_sc_hd__clkbuf_1
Xwire2296 net2297 VGND VGND VPWR VPWR net2296 sky130_fd_sc_hd__buf_1
Xwire1551 net1552 VGND VGND VPWR VPWR net1551 sky130_fd_sc_hd__buf_1
X_19540_ net3153 net6098 VGND VGND VPWR VPWR _11377_ sky130_fd_sc_hd__nand2_1
X_16752_ net7561 net9230 net3380 VGND VGND VPWR VPWR _08765_ sky130_fd_sc_hd__mux2_1
X_13964_ net7718 net1571 VGND VGND VPWR VPWR _06229_ sky130_fd_sc_hd__nand2_1
Xwire1562 _05973_ VGND VGND VPWR VPWR net1562 sky130_fd_sc_hd__clkbuf_1
Xwire1573 net1574 VGND VGND VPWR VPWR net1573 sky130_fd_sc_hd__clkbuf_1
Xwire1584 _05504_ VGND VGND VPWR VPWR net1584 sky130_fd_sc_hd__buf_1
X_15703_ net1097 _07773_ VGND VGND VPWR VPWR _07774_ sky130_fd_sc_hd__xor2_1
XFILLER_0_88_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12915_ net7909 _05187_ VGND VGND VPWR VPWR _05188_ sky130_fd_sc_hd__nand2_1
Xwire1595 _05135_ VGND VGND VPWR VPWR net1595 sky130_fd_sc_hd__clkbuf_1
X_16683_ matmul0.alpha_pass\[9\] net619 net6550 VGND VGND VPWR VPWR _08715_ sky130_fd_sc_hd__mux2_1
X_19471_ net3895 net2514 _11265_ VGND VGND VPWR VPWR _11308_ sky130_fd_sc_hd__mux2_1
X_13895_ _06125_ _06135_ VGND VGND VPWR VPWR _06161_ sky130_fd_sc_hd__nor2_1
X_15634_ _07597_ _07704_ _07705_ VGND VGND VPWR VPWR _07706_ sky130_fd_sc_hd__a21o_1
X_18422_ _10155_ _10271_ VGND VGND VPWR VPWR _10272_ sky130_fd_sc_hd__nand2_1
X_12846_ _05038_ _05043_ VGND VGND VPWR VPWR _05119_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18353_ _10186_ _10189_ _10190_ VGND VGND VPWR VPWR _10204_ sky130_fd_sc_hd__a21o_1
XFILLER_0_150_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15565_ _07636_ _07637_ VGND VGND VPWR VPWR _07638_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12777_ net6673 net6678 net7275 VGND VGND VPWR VPWR _05050_ sky130_fd_sc_hd__and3b_1
X_17304_ net7661 _09213_ _09217_ net7643 VGND VGND VPWR VPWR _09218_ sky130_fd_sc_hd__o211ai_1
Xmax_length6280 net6281 VGND VGND VPWR VPWR net6280 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_185_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14516_ net7302 net5262 _06694_ _06696_ net1990 VGND VGND VPWR VPWR _06697_ sky130_fd_sc_hd__o311a_1
X_18284_ _10133_ _10055_ _10134_ VGND VGND VPWR VPWR _10135_ sky130_fd_sc_hd__a21oi_1
X_15496_ _07543_ _07563_ _07565_ _07568_ VGND VGND VPWR VPWR _07569_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_44_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17235_ net2186 _09182_ _09023_ VGND VGND VPWR VPWR _09183_ sky130_fd_sc_hd__a21o_1
X_14447_ _06639_ VGND VGND VPWR VPWR _00096_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_104_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17166_ net670 _09118_ VGND VGND VPWR VPWR _09119_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14378_ _06586_ matmul0.a_in\[13\] net899 VGND VGND VPWR VPWR _06587_ sky130_fd_sc_hd__mux2_1
Xwire870 net871 VGND VGND VPWR VPWR net870 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire881 _08446_ VGND VGND VPWR VPWR net881 sky130_fd_sc_hd__buf_1
Xwire892 net893 VGND VGND VPWR VPWR net892 sky130_fd_sc_hd__buf_1
XFILLER_0_101_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16117_ net2700 _07841_ net1515 net2630 VGND VGND VPWR VPWR _08183_ sky130_fd_sc_hd__a31o_1
X_13329_ _05598_ _05601_ VGND VGND VPWR VPWR _05602_ sky130_fd_sc_hd__xnor2_1
X_17097_ net6495 net6477 VGND VGND VPWR VPWR _09054_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16048_ net2802 net2660 VGND VGND VPWR VPWR _08115_ sky130_fd_sc_hd__nor2_1
X_19807_ _11639_ _11640_ net3150 VGND VGND VPWR VPWR _11641_ sky130_fd_sc_hd__mux2_1
X_17999_ net7135 net7118 net7109 VGND VGND VPWR VPWR _09850_ sky130_fd_sc_hd__and3b_1
XFILLER_0_193_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19738_ net6008 _11571_ net3129 VGND VGND VPWR VPWR _11573_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19669_ _11409_ _11501_ _11502_ net6066 _11504_ VGND VGND VPWR VPWR _11505_ sky130_fd_sc_hd__a221o_1
X_21700_ net5896 net3785 net3107 _01710_ VGND VGND VPWR VPWR _01711_ sky130_fd_sc_hd__a31o_1
X_22680_ _02628_ VGND VGND VPWR VPWR _00586_ sky130_fd_sc_hd__clkbuf_1
X_21631_ net4385 _01544_ net476 net4318 net1175 VGND VGND VPWR VPWR _01643_ sky130_fd_sc_hd__a221o_1
XFILLER_0_158_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24350_ _04207_ _04208_ VGND VGND VPWR VPWR _04209_ sky130_fd_sc_hd__xor2_2
XFILLER_0_35_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21562_ _01572_ _01573_ VGND VGND VPWR VPWR _01574_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7208 net7209 VGND VGND VPWR VPWR net7208 sky130_fd_sc_hd__clkbuf_1
Xwire7219 net7220 VGND VGND VPWR VPWR net7219 sky130_fd_sc_hd__clkbuf_1
X_23301_ _03160_ _03163_ _03164_ _03166_ _03170_ VGND VGND VPWR VPWR _03171_ sky130_fd_sc_hd__a32o_1
XFILLER_0_51_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20513_ net6766 net2491 net3345 VGND VGND VPWR VPWR _12300_ sky130_fd_sc_hd__mux2_1
X_24281_ _04060_ _04065_ _04140_ VGND VGND VPWR VPWR _04141_ sky130_fd_sc_hd__a21o_1
Xwire6507 net6510 VGND VGND VPWR VPWR net6507 sky130_fd_sc_hd__clkbuf_1
X_21493_ net5651 _01402_ VGND VGND VPWR VPWR _01506_ sky130_fd_sc_hd__or2_1
Xmax_length2205 net2206 VGND VGND VPWR VPWR net2205 sky130_fd_sc_hd__buf_1
Xwire6529 net6530 VGND VGND VPWR VPWR net6529 sky130_fd_sc_hd__clkbuf_1
X_23232_ _03011_ _03012_ _03101_ VGND VGND VPWR VPWR _03102_ sky130_fd_sc_hd__a21bo_1
X_20444_ _12226_ _12236_ _12237_ VGND VGND VPWR VPWR _12238_ sky130_fd_sc_hd__a21oi_1
Xwire5806 net5807 VGND VGND VPWR VPWR net5806 sky130_fd_sc_hd__buf_1
Xwire5817 net5818 VGND VGND VPWR VPWR net5817 sky130_fd_sc_hd__buf_1
Xwire5828 net5829 VGND VGND VPWR VPWR net5828 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23163_ _03027_ _03032_ VGND VGND VPWR VPWR _03033_ sky130_fd_sc_hd__xor2_2
X_20375_ net6477 net1223 VGND VGND VPWR VPWR _12174_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22114_ _02024_ _02034_ _02029_ VGND VGND VPWR VPWR _02120_ sky130_fd_sc_hd__a21bo_1
X_23094_ _02932_ _02963_ VGND VGND VPWR VPWR _02964_ sky130_fd_sc_hd__xnor2_1
X_22045_ _01941_ _01952_ net1714 VGND VGND VPWR VPWR _02052_ sky130_fd_sc_hd__o21a_1
X_25804_ clknet_leaf_30_clk _00677_ net8675 VGND VGND VPWR VPWR pid_q.curr_int\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_23996_ pid_q.curr_int\[6\] net3061 net2027 _03859_ VGND VGND VPWR VPWR _00671_ sky130_fd_sc_hd__a22o_1
X_25735_ clknet_leaf_11_clk _00608_ net8602 VGND VGND VPWR VPWR pid_d.ki\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22947_ _02388_ _02834_ _02455_ net517 VGND VGND VPWR VPWR _02835_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_15_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12700_ net7943 VGND VGND VPWR VPWR _04973_ sky130_fd_sc_hd__inv_2
X_13680_ net7810 net2947 net1939 _05947_ net3677 VGND VGND VPWR VPWR _05949_ sky130_fd_sc_hd__a311oi_1
XFILLER_0_35_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25666_ clknet_leaf_120_clk _00539_ net8397 VGND VGND VPWR VPWR pid_d.prev_error\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_22878_ net4337 _02772_ _02773_ net412 net4359 VGND VGND VPWR VPWR _02774_ sky130_fd_sc_hd__a32o_1
XFILLER_0_167_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24617_ net2018 net1649 VGND VGND VPWR VPWR _04472_ sky130_fd_sc_hd__or2_1
X_12631_ net7325 _04892_ net4278 VGND VGND VPWR VPWR _04904_ sky130_fd_sc_hd__nand3_1
X_21829_ net5703 net5515 VGND VGND VPWR VPWR _01838_ sky130_fd_sc_hd__nand2_1
X_25597_ clknet_leaf_105_clk _00470_ net8354 VGND VGND VPWR VPWR cordic0.slte0.opB\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout8348 net8370 VGND VGND VPWR VPWR net8348 sky130_fd_sc_hd__buf_1
Xfanout7614 svm0.periodTop\[15\] VGND VGND VPWR VPWR net7614 sky130_fd_sc_hd__clkbuf_1
Xfanout8359 net8374 VGND VGND VPWR VPWR net8359 sky130_fd_sc_hd__clkbuf_1
Xwire8421 net8422 VGND VGND VPWR VPWR net8421 sky130_fd_sc_hd__buf_1
X_15350_ net2832 net2726 VGND VGND VPWR VPWR _07424_ sky130_fd_sc_hd__nand2_1
Xfanout7625 net7633 VGND VGND VPWR VPWR net7625 sky130_fd_sc_hd__buf_1
X_24548_ net1649 _04354_ VGND VGND VPWR VPWR _04404_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14301_ net6451 net6456 VGND VGND VPWR VPWR _06523_ sky130_fd_sc_hd__nand2_1
Xwire8454 net8456 VGND VGND VPWR VPWR net8454 sky130_fd_sc_hd__buf_1
XFILLER_0_124_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7731 net7732 VGND VGND VPWR VPWR net7731 sky130_fd_sc_hd__clkbuf_1
X_15281_ net1877 net2703 VGND VGND VPWR VPWR _07355_ sky130_fd_sc_hd__xor2_1
Xwire8476 net8477 VGND VGND VPWR VPWR net8476 sky130_fd_sc_hd__buf_1
X_24479_ _04259_ _04260_ _04334_ _04335_ VGND VGND VPWR VPWR _04336_ sky130_fd_sc_hd__a31oi_2
Xwire7753 net7754 VGND VGND VPWR VPWR net7753 sky130_fd_sc_hd__buf_1
XFILLER_0_123_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17020_ _08977_ _08980_ VGND VGND VPWR VPWR _08981_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire155 net156 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__buf_1
X_14232_ net9091 _05779_ net154 net2373 VGND VGND VPWR VPWR _00031_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7775 net7776 VGND VGND VPWR VPWR net7775 sky130_fd_sc_hd__clkbuf_1
Xwire166 _08634_ VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length3473 _07152_ VGND VGND VPWR VPWR net3473 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire177 _04640_ VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_1
Xwire188 _06363_ VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__buf_1
Xwire7797 net7798 VGND VGND VPWR VPWR net7797 sky130_fd_sc_hd__clkbuf_1
Xwire199 net200 VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_1
X_14163_ net217 net403 _06368_ VGND VGND VPWR VPWR _06424_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13114_ _05383_ _05386_ VGND VGND VPWR VPWR _05387_ sky130_fd_sc_hd__xnor2_1
X_14094_ _06282_ _06315_ _06317_ VGND VGND VPWR VPWR _06357_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18971_ _10795_ _10806_ _10807_ VGND VGND VPWR VPWR _10808_ sky130_fd_sc_hd__a21boi_2
X_13045_ _05306_ _05310_ VGND VGND VPWR VPWR _05318_ sky130_fd_sc_hd__and2_1
Xclkbuf_4_2__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_4_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_17922_ _09665_ _09669_ _09772_ VGND VGND VPWR VPWR _09773_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17853_ net7043 net7111 VGND VGND VPWR VPWR _09704_ sky130_fd_sc_hd__nor2_1
Xwire2060 net2061 VGND VGND VPWR VPWR net2060 sky130_fd_sc_hd__clkbuf_2
Xwire2071 net2072 VGND VGND VPWR VPWR net2071 sky130_fd_sc_hd__clkbuf_1
Xwire2082 net2083 VGND VGND VPWR VPWR net2082 sky130_fd_sc_hd__clkbuf_2
X_16804_ net4287 VGND VGND VPWR VPWR _08792_ sky130_fd_sc_hd__buf_1
X_14996_ net1898 _07060_ _07069_ VGND VGND VPWR VPWR _07070_ sky130_fd_sc_hd__a21bo_1
Xwire2093 net2094 VGND VGND VPWR VPWR net2093 sky130_fd_sc_hd__clkbuf_2
X_17784_ net6986 net6942 VGND VGND VPWR VPWR _09635_ sky130_fd_sc_hd__xnor2_1
Xwire1370 _04530_ VGND VGND VPWR VPWR net1370 sky130_fd_sc_hd__buf_1
XFILLER_0_191_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1381 net1382 VGND VGND VPWR VPWR net1381 sky130_fd_sc_hd__clkbuf_1
X_19523_ _11359_ net3158 _11297_ VGND VGND VPWR VPWR _11360_ sky130_fd_sc_hd__a21o_1
X_13947_ _06159_ _06211_ _06212_ VGND VGND VPWR VPWR _06213_ sky130_fd_sc_hd__and3_1
XFILLER_0_163_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1392 _00890_ VGND VGND VPWR VPWR net1392 sky130_fd_sc_hd__buf_1
X_16735_ net9226 matmul0.b\[4\] net3703 VGND VGND VPWR VPWR _08756_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19454_ net3866 _11290_ VGND VGND VPWR VPWR _11291_ sky130_fd_sc_hd__xnor2_1
X_16666_ _08698_ _08694_ _08699_ VGND VGND VPWR VPWR _08700_ sky130_fd_sc_hd__a21o_1
X_13878_ net532 _06081_ VGND VGND VPWR VPWR _06145_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15617_ net3444 _07688_ VGND VGND VPWR VPWR _07689_ sky130_fd_sc_hd__and2_1
X_18405_ _10249_ _10255_ VGND VGND VPWR VPWR _10256_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12829_ _05093_ _05101_ VGND VGND VPWR VPWR _05102_ sky130_fd_sc_hd__xnor2_1
X_16597_ _08644_ net3389 net3388 VGND VGND VPWR VPWR _08648_ sky130_fd_sc_hd__mux2_1
X_19385_ _11220_ _11221_ VGND VGND VPWR VPWR _11222_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15548_ _07526_ _07527_ _07620_ VGND VGND VPWR VPWR _07621_ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18336_ _10121_ net1776 VGND VGND VPWR VPWR _10187_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18267_ _10044_ _10046_ VGND VGND VPWR VPWR _10118_ sky130_fd_sc_hd__or2_1
X_15479_ _07548_ _07549_ _07552_ VGND VGND VPWR VPWR _07553_ sky130_fd_sc_hd__nand3_1
XFILLER_0_4_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17218_ _09162_ _09166_ VGND VGND VPWR VPWR _09167_ sky130_fd_sc_hd__xnor2_1
X_18198_ _10044_ _10046_ net3233 _10048_ VGND VGND VPWR VPWR _10049_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_141_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17149_ net6914 _09086_ VGND VGND VPWR VPWR _09103_ sky130_fd_sc_hd__and2_1
XFILLER_0_123_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20160_ net868 _11986_ VGND VGND VPWR VPWR _11987_ sky130_fd_sc_hd__xnor2_1
X_20091_ _11841_ _11843_ _11919_ _11846_ VGND VGND VPWR VPWR _11920_ sky130_fd_sc_hd__a31o_1
XFILLER_0_196_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23850_ _03623_ _03625_ _03714_ VGND VGND VPWR VPWR _03715_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_58_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22801_ _02708_ VGND VGND VPWR VPWR _00627_ sky130_fd_sc_hd__clkbuf_1
X_23781_ _03645_ _03646_ net4748 VGND VGND VPWR VPWR _03647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20993_ net1734 _01007_ _01008_ VGND VGND VPWR VPWR _01009_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_196_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25520_ clknet_leaf_42_clk _00400_ net8773 VGND VGND VPWR VPWR svm0.counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_177_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22732_ net3718 net105 VGND VGND VPWR VPWR _02666_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25451_ clknet_leaf_119_clk _00334_ net8342 VGND VGND VPWR VPWR cordic0.vec\[1\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_177_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22663_ _02407_ net3079 net800 _02616_ net8905 VGND VGND VPWR VPWR _00581_ sky130_fd_sc_hd__o311a_1
XFILLER_0_109_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24402_ pid_q.prev_int\[11\] _04189_ VGND VGND VPWR VPWR _04260_ sky130_fd_sc_hd__or2_1
X_21614_ _01619_ _01624_ VGND VGND VPWR VPWR _01626_ sky130_fd_sc_hd__or2_1
X_25382_ clknet_leaf_74_clk _00265_ net8473 VGND VGND VPWR VPWR matmul0.b\[1\] sky130_fd_sc_hd__dfrtp_1
X_22594_ _02569_ _02570_ net3768 VGND VGND VPWR VPWR _02571_ sky130_fd_sc_hd__and3b_1
Xwire7005 net7006 VGND VGND VPWR VPWR net7005 sky130_fd_sc_hd__buf_1
XFILLER_0_29_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7016 net7017 VGND VGND VPWR VPWR net7016 sky130_fd_sc_hd__buf_1
X_24333_ _04026_ _04107_ VGND VGND VPWR VPWR _04192_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21545_ net3839 net5653 VGND VGND VPWR VPWR _01557_ sky130_fd_sc_hd__nand2_1
XFILLER_0_161_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7038 net7034 VGND VGND VPWR VPWR net7038 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_7_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6304 net6305 VGND VGND VPWR VPWR net6304 sky130_fd_sc_hd__buf_1
XFILLER_0_65_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24264_ net4580 net4836 VGND VGND VPWR VPWR _04124_ sky130_fd_sc_hd__nand2_1
X_21476_ _01373_ _01375_ _01488_ VGND VGND VPWR VPWR _01489_ sky130_fd_sc_hd__a21oi_2
Xwire5603 net5605 VGND VGND VPWR VPWR net5603 sky130_fd_sc_hd__buf_1
Xwire6348 net6349 VGND VGND VPWR VPWR net6348 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length1301 net1302 VGND VGND VPWR VPWR net1301 sky130_fd_sc_hd__buf_1
XFILLER_0_132_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6359 net6361 VGND VGND VPWR VPWR net6359 sky130_fd_sc_hd__buf_1
Xmax_length2046 net2047 VGND VGND VPWR VPWR net2046 sky130_fd_sc_hd__buf_1
X_23215_ _03082_ _03083_ _03084_ VGND VGND VPWR VPWR _03085_ sky130_fd_sc_hd__or3_1
Xfanout4829 pid_q.mult0.b\[13\] VGND VGND VPWR VPWR net4829 sky130_fd_sc_hd__buf_1
Xmax_length2068 _01779_ VGND VGND VPWR VPWR net2068 sky130_fd_sc_hd__buf_1
X_20427_ cordic0.slte0.opA\[11\] net1559 VGND VGND VPWR VPWR _12223_ sky130_fd_sc_hd__nor2_1
X_24195_ _04054_ _04055_ VGND VGND VPWR VPWR _04056_ sky130_fd_sc_hd__xor2_2
Xwire5647 net5648 VGND VGND VPWR VPWR net5647 sky130_fd_sc_hd__clkbuf_2
Xwire4913 net4915 VGND VGND VPWR VPWR net4913 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire5658 net5659 VGND VGND VPWR VPWR net5658 sky130_fd_sc_hd__clkbuf_1
Xwire4924 net4925 VGND VGND VPWR VPWR net4924 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4935 net4936 VGND VGND VPWR VPWR net4935 sky130_fd_sc_hd__clkbuf_1
X_23146_ net5112 net4697 VGND VGND VPWR VPWR _03016_ sky130_fd_sc_hd__nand2_1
Xwire4946 net4947 VGND VGND VPWR VPWR net4946 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20358_ net6458 _12158_ VGND VGND VPWR VPWR _12159_ sky130_fd_sc_hd__nor2_2
Xwire4957 net4958 VGND VGND VPWR VPWR net4957 sky130_fd_sc_hd__buf_1
XFILLER_0_105_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4968 net4969 VGND VGND VPWR VPWR net4968 sky130_fd_sc_hd__buf_1
XFILLER_0_140_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4979 pid_q.mult0.b\[7\] VGND VGND VPWR VPWR net4979 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23077_ _02880_ _02885_ VGND VGND VPWR VPWR _02947_ sky130_fd_sc_hd__nand2_1
X_20289_ net4041 _06504_ VGND VGND VPWR VPWR _12095_ sky130_fd_sc_hd__or2_1
XFILLER_0_140_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22028_ _02029_ _02034_ VGND VGND VPWR VPWR _02035_ sky130_fd_sc_hd__xnor2_1
Xhold30 pid_q.curr_error\[13\] VGND VGND VPWR VPWR net8983 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 matmul0.matmul_stage_inst.b\[5\] VGND VGND VPWR VPWR net8994 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 svm0.vC\[6\] VGND VGND VPWR VPWR net9005 sky130_fd_sc_hd__dlygate4sd3_1
X_14850_ _06942_ VGND VGND VPWR VPWR _00196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold63 cordic0.sin\[5\] VGND VGND VPWR VPWR net9016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 cordic0.sin\[1\] VGND VGND VPWR VPWR net9027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 cordic0.cos\[7\] VGND VGND VPWR VPWR net9038 sky130_fd_sc_hd__dlygate4sd3_1
X_13801_ net7810 net1319 net1923 _06068_ VGND VGND VPWR VPWR _06069_ sky130_fd_sc_hd__a22o_1
Xhold96 cordic0.cos\[0\] VGND VGND VPWR VPWR net9049 sky130_fd_sc_hd__dlygate4sd3_1
X_14781_ net7148 _06858_ _06817_ VGND VGND VPWR VPWR _06905_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_187_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23979_ _03842_ VGND VGND VPWR VPWR _03843_ sky130_fd_sc_hd__inv_2
X_16520_ _08572_ _08579_ VGND VGND VPWR VPWR _08580_ sky130_fd_sc_hd__xnor2_1
X_13732_ net503 _06000_ VGND VGND VPWR VPWR _06001_ sky130_fd_sc_hd__or2b_1
X_25718_ clknet_leaf_12_clk _00591_ net8605 VGND VGND VPWR VPWR pid_d.mult0.a\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_10__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_4_10__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16451_ net2623 net2217 VGND VGND VPWR VPWR _08512_ sky130_fd_sc_hd__nor2_1
X_13663_ _05919_ _05932_ VGND VGND VPWR VPWR _05933_ sky130_fd_sc_hd__xnor2_1
X_25649_ clknet_leaf_1_clk _00522_ net8403 VGND VGND VPWR VPWR pid_d.curr_int\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_15402_ net2838 net2768 VGND VGND VPWR VPWR _07476_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12614_ _04865_ _04887_ VGND VGND VPWR VPWR _00002_ sky130_fd_sc_hd__nor2_1
X_19170_ _11002_ _11006_ VGND VGND VPWR VPWR _11007_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16382_ _08441_ _08443_ net2629 VGND VGND VPWR VPWR _08444_ sky130_fd_sc_hd__a21o_1
X_13594_ net577 _05845_ net679 VGND VGND VPWR VPWR _05864_ sky130_fd_sc_hd__o21ba_1
Xwire8240 net8241 VGND VGND VPWR VPWR net8240 sky130_fd_sc_hd__clkbuf_1
X_18121_ _09899_ _09950_ _09971_ VGND VGND VPWR VPWR _09972_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15333_ _07124_ net1117 VGND VGND VPWR VPWR _07407_ sky130_fd_sc_hd__and2_1
XFILLER_0_108_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8251 net8252 VGND VGND VPWR VPWR net8251 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout7455 net7460 VGND VGND VPWR VPWR net7455 sky130_fd_sc_hd__buf_1
Xfanout7466 pid_q.state\[5\] VGND VGND VPWR VPWR net7466 sky130_fd_sc_hd__clkbuf_2
Xwire8262 net8263 VGND VGND VPWR VPWR net8262 sky130_fd_sc_hd__clkbuf_1
Xwire8273 net8274 VGND VGND VPWR VPWR net8273 sky130_fd_sc_hd__clkbuf_1
Xwire8284 net23 VGND VGND VPWR VPWR net8284 sky130_fd_sc_hd__clkbuf_1
Xwire8295 net8296 VGND VGND VPWR VPWR net8295 sky130_fd_sc_hd__clkbuf_1
Xwire7550 matmul0.op_in\[1\] VGND VGND VPWR VPWR net7550 sky130_fd_sc_hd__clkbuf_1
X_18052_ net7009 net7128 net3969 _09902_ VGND VGND VPWR VPWR _09903_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15264_ net1886 _07234_ _07259_ _07262_ _07337_ VGND VGND VPWR VPWR _07338_ sky130_fd_sc_hd__a311o_1
Xwire7561 matmul0.b_in\[12\] VGND VGND VPWR VPWR net7561 sky130_fd_sc_hd__clkbuf_1
Xfanout6765 cordic0.vec\[1\]\[17\] VGND VGND VPWR VPWR net6765 sky130_fd_sc_hd__clkbuf_1
Xwire7572 matmul0.b_in\[5\] VGND VGND VPWR VPWR net7572 sky130_fd_sc_hd__clkbuf_1
Xwire7583 net7584 VGND VGND VPWR VPWR net7583 sky130_fd_sc_hd__clkbuf_1
X_17003_ net7080 net1552 VGND VGND VPWR VPWR _08965_ sky130_fd_sc_hd__nor2_1
X_14215_ _06471_ _06472_ _06473_ VGND VGND VPWR VPWR _06474_ sky130_fd_sc_hd__o21ba_1
Xwire7594 matmul0.a_in\[11\] VGND VGND VPWR VPWR net7594 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6860 net6858 VGND VGND VPWR VPWR net6860 sky130_fd_sc_hd__clkbuf_2
X_15195_ _07268_ net3486 _07140_ net2845 VGND VGND VPWR VPWR _07269_ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6882 net6879 VGND VGND VPWR VPWR net6882 sky130_fd_sc_hd__buf_1
XFILLER_0_21_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6893 net6894 VGND VGND VPWR VPWR net6893 sky130_fd_sc_hd__buf_1
X_14146_ net7612 _05346_ _05709_ VGND VGND VPWR VPWR _06407_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14077_ _06221_ net1125 _06335_ net1597 _06339_ VGND VGND VPWR VPWR _06340_ sky130_fd_sc_hd__o221a_1
X_18954_ net6189 net6143 VGND VGND VPWR VPWR _10791_ sky130_fd_sc_hd__nand2_1
X_13028_ _05159_ _05300_ _05162_ _05163_ VGND VGND VPWR VPWR _05301_ sky130_fd_sc_hd__a211o_1
X_17905_ _09751_ _09755_ VGND VGND VPWR VPWR _09756_ sky130_fd_sc_hd__nor2_1
X_18885_ net657 _10726_ VGND VGND VPWR VPWR _10727_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17836_ net2559 _09686_ VGND VGND VPWR VPWR _09687_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17767_ net7092 net3996 net7116 VGND VGND VPWR VPWR _09618_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14979_ _07046_ _07052_ VGND VGND VPWR VPWR _07053_ sky130_fd_sc_hd__xnor2_1
X_19506_ _11276_ _11277_ VGND VGND VPWR VPWR _11343_ sky130_fd_sc_hd__nor2_1
X_16718_ matmul0.alpha_pass\[14\] _08744_ net6557 VGND VGND VPWR VPWR _08745_ sky130_fd_sc_hd__mux2_1
X_17698_ pid_q.state\[0\] net7521 net7463 VGND VGND VPWR VPWR _09574_ sky130_fd_sc_hd__or3_1
XFILLER_0_117_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19437_ net6147 net6155 VGND VGND VPWR VPWR _11274_ sky130_fd_sc_hd__nand2_1
X_16649_ _08685_ VGND VGND VPWR VPWR _00252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_190_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19368_ net1193 _11204_ VGND VGND VPWR VPWR _11205_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_162_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18319_ net6903 net6887 VGND VGND VPWR VPWR _10170_ sky130_fd_sc_hd__and2b_1
XFILLER_0_143_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19299_ net6319 net3191 _10986_ VGND VGND VPWR VPWR _11136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21330_ net5705 net5598 VGND VGND VPWR VPWR _01344_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21261_ _01270_ _01275_ VGND VGND VPWR VPWR _01276_ sky130_fd_sc_hd__xnor2_2
Xwire4209 _06972_ VGND VGND VPWR VPWR net4209 sky130_fd_sc_hd__clkbuf_1
X_23000_ _02869_ VGND VGND VPWR VPWR _02870_ sky130_fd_sc_hd__buf_1
X_20212_ net8953 _12034_ VGND VGND VPWR VPWR _12035_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21192_ _01189_ _01188_ VGND VGND VPWR VPWR _01208_ sky130_fd_sc_hd__or2_1
Xwire3519 net3520 VGND VGND VPWR VPWR net3519 sky130_fd_sc_hd__clkbuf_1
X_20143_ _11968_ _11949_ net2493 VGND VGND VPWR VPWR _11970_ sky130_fd_sc_hd__o21a_1
Xwire2807 _07108_ VGND VGND VPWR VPWR net2807 sky130_fd_sc_hd__buf_1
Xwire2818 net2819 VGND VGND VPWR VPWR net2818 sky130_fd_sc_hd__clkbuf_1
Xwire2829 net2830 VGND VGND VPWR VPWR net2829 sky130_fd_sc_hd__buf_1
X_24951_ net8871 net8881 VGND VGND VPWR VPWR _04728_ sky130_fd_sc_hd__and2b_1
X_20074_ net2582 _11900_ _11902_ VGND VGND VPWR VPWR _11903_ sky130_fd_sc_hd__a21o_1
XFILLER_0_148_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23902_ _03764_ _03765_ VGND VGND VPWR VPWR _03767_ sky130_fd_sc_hd__or2_1
X_24882_ _04679_ VGND VGND VPWR VPWR _00737_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23833_ _03694_ _03697_ VGND VGND VPWR VPWR _03698_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_169_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23764_ _03532_ _03534_ _03530_ VGND VGND VPWR VPWR _03630_ sky130_fd_sc_hd__a21bo_1
Xmax_length6802 net6797 VGND VGND VPWR VPWR net6802 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_170_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20976_ _00983_ _00986_ _00991_ VGND VGND VPWR VPWR _00992_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_68_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25503_ clknet_leaf_39_clk _00383_ net8771 VGND VGND VPWR VPWR svm0.delta\[8\] sky130_fd_sc_hd__dfrtp_1
X_22715_ _02651_ net5374 net3094 VGND VGND VPWR VPWR _02652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23695_ _03453_ _03460_ VGND VGND VPWR VPWR _03562_ sky130_fd_sc_hd__or2_1
Xmax_length6857 net6854 VGND VGND VPWR VPWR net6857 sky130_fd_sc_hd__buf_1
X_25434_ clknet_leaf_94_clk _00317_ net8445 VGND VGND VPWR VPWR matmul0.sin\[7\] sky130_fd_sc_hd__dfrtp_1
X_22646_ _01863_ net3077 VGND VGND VPWR VPWR _02608_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25365_ clknet_leaf_72_clk _00248_ net8478 VGND VGND VPWR VPWR matmul0.alpha_pass\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_114_clk clknet_4_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_114_clk
+ sky130_fd_sc_hd__clkbuf_16
X_22577_ net7317 _02554_ VGND VGND VPWR VPWR _02557_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout6028 net6036 VGND VGND VPWR VPWR net6028 sky130_fd_sc_hd__buf_1
Xwire6101 net6102 VGND VGND VPWR VPWR net6101 sky130_fd_sc_hd__dlymetal6s2s_1
X_24316_ _04174_ _04175_ VGND VGND VPWR VPWR _04176_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6112 net6109 VGND VGND VPWR VPWR net6112 sky130_fd_sc_hd__dlymetal6s2s_1
X_21528_ pid_d.curr_int\[3\] net3122 net2077 _01540_ VGND VGND VPWR VPWR _00522_ sky130_fd_sc_hd__a22o_1
Xwire6123 net6122 VGND VGND VPWR VPWR net6123 sky130_fd_sc_hd__buf_1
X_25296_ clknet_leaf_92_clk _00179_ net8429 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.d\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire6134 net6132 VGND VGND VPWR VPWR net6134 sky130_fd_sc_hd__buf_1
Xwire5400 net5401 VGND VGND VPWR VPWR net5400 sky130_fd_sc_hd__buf_1
Xwire6145 net6138 VGND VGND VPWR VPWR net6145 sky130_fd_sc_hd__buf_1
Xwire5411 net5412 VGND VGND VPWR VPWR net5411 sky130_fd_sc_hd__buf_1
X_24247_ _04045_ _04107_ VGND VGND VPWR VPWR _04108_ sky130_fd_sc_hd__xnor2_1
Xwire5422 pid_d.mult0.a\[13\] VGND VGND VPWR VPWR net5422 sky130_fd_sc_hd__buf_1
X_21459_ _01343_ _01345_ _01471_ VGND VGND VPWR VPWR _01472_ sky130_fd_sc_hd__a21oi_2
Xwire6167 net6164 VGND VGND VPWR VPWR net6167 sky130_fd_sc_hd__clkbuf_1
Xwire6178 net6177 VGND VGND VPWR VPWR net6178 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_32_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14000_ net529 _06264_ VGND VGND VPWR VPWR _06265_ sky130_fd_sc_hd__xnor2_2
Xwire6189 net6190 VGND VGND VPWR VPWR net6189 sky130_fd_sc_hd__buf_1
Xwire5444 net5445 VGND VGND VPWR VPWR net5444 sky130_fd_sc_hd__clkbuf_1
Xwire4710 net4711 VGND VGND VPWR VPWR net4710 sky130_fd_sc_hd__clkbuf_1
Xwire5455 net5456 VGND VGND VPWR VPWR net5455 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire5466 net5459 VGND VGND VPWR VPWR net5466 sky130_fd_sc_hd__buf_1
Xwire4732 net4733 VGND VGND VPWR VPWR net4732 sky130_fd_sc_hd__buf_1
X_24178_ _04037_ _03957_ _04038_ VGND VGND VPWR VPWR _04039_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5477 net5471 VGND VGND VPWR VPWR net5477 sky130_fd_sc_hd__clkbuf_1
Xwire4743 net4741 VGND VGND VPWR VPWR net4743 sky130_fd_sc_hd__buf_1
Xwire5488 net5478 VGND VGND VPWR VPWR net5488 sky130_fd_sc_hd__buf_1
Xwire4754 net4755 VGND VGND VPWR VPWR net4754 sky130_fd_sc_hd__buf_1
Xwire5499 net5500 VGND VGND VPWR VPWR net5499 sky130_fd_sc_hd__buf_1
Xwire4765 net4766 VGND VGND VPWR VPWR net4765 sky130_fd_sc_hd__buf_1
X_23129_ _02996_ _02997_ VGND VGND VPWR VPWR _02999_ sky130_fd_sc_hd__nor2_1
Xwire4776 net4777 VGND VGND VPWR VPWR net4776 sky130_fd_sc_hd__buf_1
XFILLER_0_128_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15951_ net2693 _07156_ VGND VGND VPWR VPWR _08019_ sky130_fd_sc_hd__nor2_1
Xinput120 pid_q_addr[15] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_1
Xinput131 pid_q_data[10] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_1
Xinput142 pid_q_data[6] VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_1
X_14902_ net6630 matmul0.matmul_stage_inst.d\[10\] net7406 net6532 VGND VGND VPWR
+ VPWR _06976_ sky130_fd_sc_hd__a22o_1
X_15882_ net3448 net3413 VGND VGND VPWR VPWR _07951_ sky130_fd_sc_hd__nor2_1
X_18670_ _10407_ _10515_ VGND VGND VPWR VPWR _10516_ sky130_fd_sc_hd__nor2_1
X_17621_ net4012 svm0.tB\[1\] VGND VGND VPWR VPWR _09502_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14833_ _06933_ VGND VGND VPWR VPWR _00188_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17552_ net4006 svm0.tC\[7\] _09433_ VGND VGND VPWR VPWR _09434_ sky130_fd_sc_hd__a21bo_1
X_14764_ net7151 _06892_ VGND VGND VPWR VPWR _06893_ sky130_fd_sc_hd__xor2_1
XFILLER_0_187_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13715_ _05961_ _05983_ VGND VGND VPWR VPWR _05984_ sky130_fd_sc_hd__xnor2_1
X_16503_ _08559_ _08562_ VGND VGND VPWR VPWR _08563_ sky130_fd_sc_hd__xor2_1
X_17483_ net3273 _09373_ net6661 VGND VGND VPWR VPWR _09374_ sky130_fd_sc_hd__o21ai_1
X_14695_ net9036 net2862 net2262 net2260 VGND VGND VPWR VPWR _00142_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19222_ _11048_ _11057_ net6139 VGND VGND VPWR VPWR _11059_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_4_Left_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13646_ _05914_ _05915_ VGND VGND VPWR VPWR _05916_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16434_ _08428_ _08480_ _08481_ _08494_ VGND VGND VPWR VPWR _08495_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19153_ net6323 _10989_ net3901 VGND VGND VPWR VPWR _10990_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16365_ _08424_ net773 VGND VGND VPWR VPWR _08428_ sky130_fd_sc_hd__nand2_2
X_13577_ _05784_ net533 VGND VGND VPWR VPWR _05848_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_105_clk clknet_4_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_105_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_54_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8070 net8071 VGND VGND VPWR VPWR net8070 sky130_fd_sc_hd__clkbuf_1
X_18104_ _09092_ _09738_ VGND VGND VPWR VPWR _09955_ sky130_fd_sc_hd__xnor2_1
X_15316_ net3495 net3553 VGND VGND VPWR VPWR _07390_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8081 net8082 VGND VGND VPWR VPWR net8081 sky130_fd_sc_hd__clkbuf_1
Xwire8092 net8093 VGND VGND VPWR VPWR net8092 sky130_fd_sc_hd__clkbuf_1
X_19084_ _10911_ _10914_ _10915_ _10916_ _10920_ VGND VGND VPWR VPWR _10921_ sky130_fd_sc_hd__o32a_1
X_16296_ net491 _08297_ _08299_ VGND VGND VPWR VPWR _08360_ sky130_fd_sc_hd__and3_1
XFILLER_0_83_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7380 matmul0.matmul_stage_inst.f\[14\] VGND VGND VPWR VPWR net7380 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18035_ net2556 _09885_ VGND VGND VPWR VPWR _09886_ sky130_fd_sc_hd__xnor2_1
X_15247_ _07319_ _07320_ net2832 net3453 VGND VGND VPWR VPWR _07321_ sky130_fd_sc_hd__o211a_1
Xfanout6584 net6586 VGND VGND VPWR VPWR net6584 sky130_fd_sc_hd__clkbuf_1
Xwire7391 matmul0.matmul_stage_inst.e\[8\] VGND VGND VPWR VPWR net7391 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5883 net5899 VGND VGND VPWR VPWR net5883 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_23_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15178_ net1883 _07250_ VGND VGND VPWR VPWR _07252_ sky130_fd_sc_hd__nor2_1
X_14129_ _06385_ _06345_ _06389_ _06291_ _06390_ VGND VGND VPWR VPWR _06391_ sky130_fd_sc_hd__o221a_1
X_19986_ _11814_ _11815_ VGND VGND VPWR VPWR _11817_ sky130_fd_sc_hd__or2_1
X_18937_ net6813 net6779 _10775_ net6830 net6796 VGND VGND VPWR VPWR _10776_ sky130_fd_sc_hd__a221o_1
XFILLER_0_158_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18868_ net6832 net3224 VGND VGND VPWR VPWR _10710_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17819_ _09666_ _09669_ VGND VGND VPWR VPWR _09670_ sky130_fd_sc_hd__nand2_1
X_18799_ net6784 _10641_ _10642_ net6800 VGND VGND VPWR VPWR _10643_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20830_ _12560_ _12561_ _00845_ VGND VGND VPWR VPWR _00846_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20761_ _12511_ _12531_ VGND VGND VPWR VPWR _12532_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_59_Left_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22500_ _02443_ _02439_ VGND VGND VPWR VPWR _02501_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23480_ _03335_ _03348_ VGND VGND VPWR VPWR _03349_ sky130_fd_sc_hd__xnor2_2
X_20692_ net3143 _12459_ _12458_ VGND VGND VPWR VPWR _12467_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_76_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22431_ net5723 net5749 _02432_ VGND VGND VPWR VPWR _02433_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_150_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25150_ clknet_leaf_41_clk _00039_ net8767 VGND VGND VPWR VPWR pid_q.target\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22362_ _02360_ _02363_ VGND VGND VPWR VPWR _02365_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24101_ net3743 _03887_ _03962_ VGND VGND VPWR VPWR _03963_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21313_ _01325_ net758 VGND VGND VPWR VPWR _01328_ sky130_fd_sc_hd__nor2_1
X_25081_ _04824_ _04825_ VGND VGND VPWR VPWR _04827_ sky130_fd_sc_hd__nand2_1
X_22293_ _02288_ _02296_ VGND VGND VPWR VPWR _02297_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4006 net4007 VGND VGND VPWR VPWR net4006 sky130_fd_sc_hd__clkbuf_2
X_24032_ net4578 net4906 VGND VGND VPWR VPWR _03895_ sky130_fd_sc_hd__nand2_1
Xwire4017 net4018 VGND VGND VPWR VPWR net4017 sky130_fd_sc_hd__buf_1
X_21244_ net5811 net5510 VGND VGND VPWR VPWR _01259_ sky130_fd_sc_hd__nand2_1
Xwire4028 net4029 VGND VGND VPWR VPWR net4028 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_68_Left_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4039 net4042 VGND VGND VPWR VPWR net4039 sky130_fd_sc_hd__buf_1
Xwire3305 _09082_ VGND VGND VPWR VPWR net3305 sky130_fd_sc_hd__buf_2
Xwire3316 net3317 VGND VGND VPWR VPWR net3316 sky130_fd_sc_hd__buf_1
XFILLER_0_159_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3327 _09006_ VGND VGND VPWR VPWR net3327 sky130_fd_sc_hd__buf_1
X_21175_ net5881 _01190_ VGND VGND VPWR VPWR _01191_ sky130_fd_sc_hd__nand2_1
Xwire3338 net3339 VGND VGND VPWR VPWR net3338 sky130_fd_sc_hd__clkbuf_1
Xwire2604 _08970_ VGND VGND VPWR VPWR net2604 sky130_fd_sc_hd__buf_1
Xwire3349 _08914_ VGND VGND VPWR VPWR net3349 sky130_fd_sc_hd__buf_1
Xwire2615 _08648_ VGND VGND VPWR VPWR net2615 sky130_fd_sc_hd__buf_1
XFILLER_0_110_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20126_ net1055 _11953_ VGND VGND VPWR VPWR _11954_ sky130_fd_sc_hd__nor2_1
Xwire2637 _07864_ VGND VGND VPWR VPWR net2637 sky130_fd_sc_hd__buf_1
XFILLER_0_102_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1903 net1904 VGND VGND VPWR VPWR net1903 sky130_fd_sc_hd__clkbuf_1
Xwire2648 net2649 VGND VGND VPWR VPWR net2648 sky130_fd_sc_hd__clkbuf_2
Xwire1914 _06508_ VGND VGND VPWR VPWR net1914 sky130_fd_sc_hd__clkbuf_1
Xwire2659 net2660 VGND VGND VPWR VPWR net2659 sky130_fd_sc_hd__dlymetal6s2s_1
X_24934_ pid_q.ki\[7\] _04716_ net1361 VGND VGND VPWR VPWR _04717_ sky130_fd_sc_hd__mux2_1
Xwire1925 _05857_ VGND VGND VPWR VPWR net1925 sky130_fd_sc_hd__buf_1
X_20057_ _11879_ _11885_ _11861_ VGND VGND VPWR VPWR _11886_ sky130_fd_sc_hd__mux2_1
Xwire1936 net1937 VGND VGND VPWR VPWR net1936 sky130_fd_sc_hd__clkbuf_1
Xwire1947 net1948 VGND VGND VPWR VPWR net1947 sky130_fd_sc_hd__buf_1
Xmax_length8001 pid_q.target\[7\] VGND VGND VPWR VPWR net8001 sky130_fd_sc_hd__clkbuf_1
Xwire1958 net1959 VGND VGND VPWR VPWR net1958 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1969 net1970 VGND VGND VPWR VPWR net1969 sky130_fd_sc_hd__buf_1
X_24865_ net2399 VGND VGND VPWR VPWR _04668_ sky130_fd_sc_hd__clkbuf_1
X_23816_ net4573 net4941 VGND VGND VPWR VPWR _03681_ sky130_fd_sc_hd__nand2_1
X_24796_ _04618_ _04619_ _04620_ VGND VGND VPWR VPWR _04621_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_77_Left_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length7355 net7356 VGND VGND VPWR VPWR net7355 sky130_fd_sc_hd__clkbuf_1
Xmax_length7377 svm0.delta\[0\] VGND VGND VPWR VPWR net7377 sky130_fd_sc_hd__dlymetal6s2s_1
X_23747_ _03611_ _03612_ VGND VGND VPWR VPWR _03613_ sky130_fd_sc_hd__and2b_1
XFILLER_0_23_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length7388 matmul0.matmul_stage_inst.e\[10\] VGND VGND VPWR VPWR net7388 sky130_fd_sc_hd__clkbuf_1
X_20959_ _00949_ _00951_ VGND VGND VPWR VPWR _00975_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13500_ net534 _05772_ VGND VGND VPWR VPWR _05773_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_166_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length6676 svm0.state\[1\] VGND VGND VPWR VPWR net6676 sky130_fd_sc_hd__clkbuf_1
X_14480_ net9095 net831 net1292 _06665_ VGND VGND VPWR VPWR _00103_ sky130_fd_sc_hd__a22o_1
X_23678_ _03441_ _03443_ _03544_ VGND VGND VPWR VPWR _03545_ sky130_fd_sc_hd__a21o_1
XFILLER_0_181_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13431_ _05700_ _05703_ VGND VGND VPWR VPWR _05704_ sky130_fd_sc_hd__xnor2_2
X_25417_ clknet_leaf_86_clk _00300_ net8531 VGND VGND VPWR VPWR matmul0.cos\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22629_ net7192 _02593_ VGND VGND VPWR VPWR _02598_ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16150_ net2662 _08114_ _08215_ VGND VGND VPWR VPWR _08216_ sky130_fd_sc_hd__a21oi_1
X_13362_ _05573_ _05634_ VGND VGND VPWR VPWR _05635_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25348_ clknet_leaf_82_clk _00231_ net8503 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult2\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xmax_length831 net832 VGND VGND VPWR VPWR net831 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_140_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15101_ _07172_ _07173_ _07174_ VGND VGND VPWR VPWR _07175_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5146 net5161 VGND VGND VPWR VPWR net5146 sky130_fd_sc_hd__clkbuf_1
X_16081_ _08018_ _08062_ _08061_ VGND VGND VPWR VPWR _08148_ sky130_fd_sc_hd__a21o_1
X_13293_ _05482_ _05564_ VGND VGND VPWR VPWR _05566_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25279_ clknet_leaf_92_clk _00162_ net8434 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.c\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_86_Left_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5230 net5231 VGND VGND VPWR VPWR net5230 sky130_fd_sc_hd__clkbuf_1
Xwire5241 net5242 VGND VGND VPWR VPWR net5241 sky130_fd_sc_hd__clkbuf_1
X_15032_ net4171 net4166 VGND VGND VPWR VPWR _07106_ sky130_fd_sc_hd__nor2_1
Xwire5252 matmul0.beta_pass\[8\] VGND VGND VPWR VPWR net5252 sky130_fd_sc_hd__clkbuf_1
Xwire5263 net5264 VGND VGND VPWR VPWR net5263 sky130_fd_sc_hd__buf_1
Xwire5274 net5275 VGND VGND VPWR VPWR net5274 sky130_fd_sc_hd__clkbuf_1
Xwire5285 net5286 VGND VGND VPWR VPWR net5285 sky130_fd_sc_hd__clkbuf_1
X_19840_ _11631_ _11653_ net953 VGND VGND VPWR VPWR _11673_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_107_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5296 net5297 VGND VGND VPWR VPWR net5296 sky130_fd_sc_hd__buf_1
Xwire4562 net4556 VGND VGND VPWR VPWR net4562 sky130_fd_sc_hd__buf_1
Xwire4573 net4574 VGND VGND VPWR VPWR net4573 sky130_fd_sc_hd__buf_1
Xwire4584 net4585 VGND VGND VPWR VPWR net4584 sky130_fd_sc_hd__clkbuf_1
Xwire4595 net4594 VGND VGND VPWR VPWR net4595 sky130_fd_sc_hd__buf_1
X_19771_ _11600_ _11605_ VGND VGND VPWR VPWR _11606_ sky130_fd_sc_hd__xnor2_2
Xwire3861 _11549_ VGND VGND VPWR VPWR net3861 sky130_fd_sc_hd__buf_1
Xwire3872 net3873 VGND VGND VPWR VPWR net3872 sky130_fd_sc_hd__clkbuf_1
X_16983_ net6502 net6522 VGND VGND VPWR VPWR _08945_ sky130_fd_sc_hd__and2b_1
Xwire3883 _10946_ VGND VGND VPWR VPWR net3883 sky130_fd_sc_hd__buf_1
Xwire3894 _10879_ VGND VGND VPWR VPWR net3894 sky130_fd_sc_hd__buf_1
X_18722_ _10517_ _10567_ VGND VGND VPWR VPWR _10568_ sky130_fd_sc_hd__xnor2_1
X_15934_ _07997_ _08002_ VGND VGND VPWR VPWR _08003_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18653_ _10453_ _10461_ _10499_ VGND VGND VPWR VPWR _10500_ sky130_fd_sc_hd__o21a_1
X_15865_ net2761 _07927_ _07931_ net2630 VGND VGND VPWR VPWR _07934_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_95_Left_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17604_ _09483_ _09484_ VGND VGND VPWR VPWR _09485_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14816_ net7441 net7167 net3627 VGND VGND VPWR VPWR _06925_ sky130_fd_sc_hd__a21o_1
X_18584_ _10430_ _10431_ VGND VGND VPWR VPWR _10432_ sky130_fd_sc_hd__xnor2_1
X_15796_ net3427 VGND VGND VPWR VPWR _07866_ sky130_fd_sc_hd__buf_1
XFILLER_0_171_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17535_ net4253 _09417_ net3388 VGND VGND VPWR VPWR _09418_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14747_ net7448 matmul0.sin\[4\] VGND VGND VPWR VPWR _06880_ sky130_fd_sc_hd__nand2_1
XFILLER_0_188_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17466_ _09287_ _09354_ net4008 VGND VGND VPWR VPWR _09359_ sky130_fd_sc_hd__a21o_1
X_14678_ net7158 _06828_ VGND VGND VPWR VPWR _06829_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_184_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19205_ net3183 _11029_ VGND VGND VPWR VPWR _11042_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13629_ _05897_ _05898_ VGND VGND VPWR VPWR _05899_ sky130_fd_sc_hd__xnor2_1
X_16417_ _08476_ _08478_ VGND VGND VPWR VPWR _08479_ sky130_fd_sc_hd__xor2_1
XFILLER_0_183_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17397_ svm0.delta\[8\] VGND VGND VPWR VPWR _09303_ sky130_fd_sc_hd__inv_2
X_19136_ net6130 _10972_ VGND VGND VPWR VPWR _10973_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16348_ net1087 net1081 net1085 VGND VGND VPWR VPWR _08411_ sky130_fd_sc_hd__o21a_1
Xfanout7093 net7097 VGND VGND VPWR VPWR net7093 sky130_fd_sc_hd__buf_1
XFILLER_0_81_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19067_ _10885_ _10903_ VGND VGND VPWR VPWR _10904_ sky130_fd_sc_hd__xnor2_1
X_16279_ net2721 net2707 net2648 _07932_ VGND VGND VPWR VPWR _08343_ sky130_fd_sc_hd__a31o_1
XFILLER_0_42_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18018_ _09697_ _09740_ VGND VGND VPWR VPWR _09869_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19969_ net6137 net6060 VGND VGND VPWR VPWR _11800_ sky130_fd_sc_hd__xnor2_2
X_22980_ net5242 net619 net6568 VGND VGND VPWR VPWR _02858_ sky130_fd_sc_hd__mux2_1
X_21931_ _01927_ _01938_ VGND VGND VPWR VPWR _01939_ sky130_fd_sc_hd__xnor2_1
X_24650_ net7496 _04504_ VGND VGND VPWR VPWR _04505_ sky130_fd_sc_hd__nand2_1
X_21862_ net5839 net5394 _01864_ VGND VGND VPWR VPWR _01871_ sky130_fd_sc_hd__or3b_1
XFILLER_0_77_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23601_ _03379_ net745 VGND VGND VPWR VPWR _03469_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_118_Right_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20813_ _00827_ _00828_ VGND VGND VPWR VPWR _00829_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_166_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24581_ _04435_ _04436_ VGND VGND VPWR VPWR _04437_ sky130_fd_sc_hd__or2b_1
X_21793_ _01714_ _01802_ VGND VGND VPWR VPWR _01803_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23532_ net4557 net5053 VGND VGND VPWR VPWR _03400_ sky130_fd_sc_hd__nand2_1
Xmax_length5227 net5219 VGND VGND VPWR VPWR net5227 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20744_ net5940 net5454 VGND VGND VPWR VPWR _12515_ sky130_fd_sc_hd__nand2_2
XFILLER_0_92_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8817 net8818 VGND VGND VPWR VPWR net8817 sky130_fd_sc_hd__clkbuf_1
Xwire8828 net8829 VGND VGND VPWR VPWR net8828 sky130_fd_sc_hd__clkbuf_1
Xmax_length4515 net4516 VGND VGND VPWR VPWR net4515 sky130_fd_sc_hd__clkbuf_2
Xwire8839 net8840 VGND VGND VPWR VPWR net8839 sky130_fd_sc_hd__buf_1
X_23463_ _03330_ _03331_ VGND VGND VPWR VPWR _03332_ sky130_fd_sc_hd__xnor2_1
Xmax_length4548 net4549 VGND VGND VPWR VPWR net4548 sky130_fd_sc_hd__buf_1
X_20675_ net6762 _12274_ _09096_ VGND VGND VPWR VPWR _12451_ sky130_fd_sc_hd__mux2_1
Xwire507 _05683_ VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire518 net519 VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__clkbuf_1
X_25202_ clknet_leaf_81_clk _00091_ net8495 VGND VGND VPWR VPWR matmul0.b_in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire529 _06258_ VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__buf_1
X_22414_ _02367_ _02345_ _02369_ VGND VGND VPWR VPWR _02416_ sky130_fd_sc_hd__a21o_1
XFILLER_0_169_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23394_ _03216_ _03227_ _03263_ VGND VGND VPWR VPWR _03264_ sky130_fd_sc_hd__a21o_1
XFILLER_0_116_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3858 net3859 VGND VGND VPWR VPWR net3858 sky130_fd_sc_hd__buf_1
XFILLER_0_162_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25133_ clknet_leaf_52_clk _00022_ net8803 VGND VGND VPWR VPWR svm0.tC\[5\] sky130_fd_sc_hd__dfrtp_1
X_22345_ net5708 net5388 VGND VGND VPWR VPWR _02348_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25064_ net3734 _04811_ VGND VGND VPWR VPWR _04812_ sky130_fd_sc_hd__xnor2_1
X_22276_ _02233_ net1033 _02207_ VGND VGND VPWR VPWR _02280_ sky130_fd_sc_hd__a21o_1
X_24015_ _03807_ _03809_ _03877_ VGND VGND VPWR VPWR _03878_ sky130_fd_sc_hd__a21bo_1
Xwire3102 net3105 VGND VGND VPWR VPWR net3102 sky130_fd_sc_hd__buf_1
Xhold160 matmul0.matmul_stage_inst.b\[8\] VGND VGND VPWR VPWR net9113 sky130_fd_sc_hd__dlygate4sd3_1
X_21227_ net5987 net4392 VGND VGND VPWR VPWR _01243_ sky130_fd_sc_hd__xor2_1
Xhold171 pid_d.prev_error\[5\] VGND VGND VPWR VPWR net9124 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3113 _00961_ VGND VGND VPWR VPWR net3113 sky130_fd_sc_hd__clkbuf_1
Xwire3124 _12313_ VGND VGND VPWR VPWR net3124 sky130_fd_sc_hd__buf_1
Xhold182 pid_d.prev_error\[2\] VGND VGND VPWR VPWR net9135 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3135 net3136 VGND VGND VPWR VPWR net3135 sky130_fd_sc_hd__buf_1
Xwire2401 net2402 VGND VGND VPWR VPWR net2401 sky130_fd_sc_hd__clkbuf_1
Xwire3146 _11409_ VGND VGND VPWR VPWR net3146 sky130_fd_sc_hd__buf_1
Xhold193 matmul0.matmul_stage_inst.c\[14\] VGND VGND VPWR VPWR net9146 sky130_fd_sc_hd__dlygate4sd3_1
Xwire2412 _03604_ VGND VGND VPWR VPWR net2412 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3157 _11330_ VGND VGND VPWR VPWR net3157 sky130_fd_sc_hd__clkbuf_2
X_21158_ net5956 net5937 VGND VGND VPWR VPWR _01174_ sky130_fd_sc_hd__and2_1
Xwire2423 _03356_ VGND VGND VPWR VPWR net2423 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2434 net2435 VGND VGND VPWR VPWR net2434 sky130_fd_sc_hd__clkbuf_1
Xwire3179 _11055_ VGND VGND VPWR VPWR net3179 sky130_fd_sc_hd__clkbuf_1
Xwire2445 net2446 VGND VGND VPWR VPWR net2445 sky130_fd_sc_hd__buf_1
Xwire1700 net1701 VGND VGND VPWR VPWR net1700 sky130_fd_sc_hd__buf_1
Xwire1711 _02063_ VGND VGND VPWR VPWR net1711 sky130_fd_sc_hd__clkbuf_1
X_20109_ net3134 _11935_ _11936_ VGND VGND VPWR VPWR _11937_ sky130_fd_sc_hd__a21o_1
Xwire2456 _02601_ VGND VGND VPWR VPWR net2456 sky130_fd_sc_hd__clkbuf_1
X_13980_ _06118_ _06173_ net7610 VGND VGND VPWR VPWR _06245_ sky130_fd_sc_hd__or3b_1
Xwire1722 _01568_ VGND VGND VPWR VPWR net1722 sky130_fd_sc_hd__buf_1
X_21089_ net5552 net5949 net5929 net5904 VGND VGND VPWR VPWR _01105_ sky130_fd_sc_hd__a22o_1
Xwire2478 _01341_ VGND VGND VPWR VPWR net2478 sky130_fd_sc_hd__clkbuf_1
Xwire1733 _01006_ VGND VGND VPWR VPWR net1733 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_189_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2489 _12502_ VGND VGND VPWR VPWR net2489 sky130_fd_sc_hd__buf_1
Xwire1744 _12354_ VGND VGND VPWR VPWR net1744 sky130_fd_sc_hd__clkbuf_1
X_12931_ _05186_ _05203_ VGND VGND VPWR VPWR _05204_ sky130_fd_sc_hd__xnor2_2
Xwire1755 _11087_ VGND VGND VPWR VPWR net1755 sky130_fd_sc_hd__clkbuf_1
X_24917_ _04705_ VGND VGND VPWR VPWR _00746_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1766 _10299_ VGND VGND VPWR VPWR net1766 sky130_fd_sc_hd__buf_1
X_25897_ clknet_leaf_14_clk _00770_ net8620 VGND VGND VPWR VPWR pid_q.kp\[9\] sky130_fd_sc_hd__dfrtp_1
Xwire1777 _10092_ VGND VGND VPWR VPWR net1777 sky130_fd_sc_hd__buf_1
Xwire1788 _09583_ VGND VGND VPWR VPWR net1788 sky130_fd_sc_hd__buf_1
Xwire1799 net1800 VGND VGND VPWR VPWR net1799 sky130_fd_sc_hd__buf_1
X_12862_ net1960 _05134_ net3688 VGND VGND VPWR VPWR _05135_ sky130_fd_sc_hd__or3b_1
X_15650_ net2776 _07720_ _07721_ VGND VGND VPWR VPWR _07722_ sky130_fd_sc_hd__o21ai_1
X_24848_ net3727 net259 net264 VGND VGND VPWR VPWR _04657_ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length7130 cordic0.vec\[1\]\[1\] VGND VGND VPWR VPWR net7130 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14601_ net7199 net5190 VGND VGND VPWR VPWR _06774_ sky130_fd_sc_hd__xnor2_1
X_15581_ _07476_ net2677 _07652_ VGND VGND VPWR VPWR _07653_ sky130_fd_sc_hd__o21a_1
X_24779_ _04604_ _04597_ net5220 _04605_ VGND VGND VPWR VPWR _04606_ sky130_fd_sc_hd__a2bb2o_1
X_12793_ _04977_ _05058_ _05062_ _05065_ VGND VGND VPWR VPWR _05066_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_29_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17320_ net4022 _09233_ VGND VGND VPWR VPWR _09234_ sky130_fd_sc_hd__nor2_1
X_14532_ net7264 net5239 VGND VGND VPWR VPWR _06711_ sky130_fd_sc_hd__xor2_4
XFILLER_0_84_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6462 net6460 VGND VGND VPWR VPWR net6462 sky130_fd_sc_hd__buf_1
XFILLER_0_141_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6495 net6496 VGND VGND VPWR VPWR net6495 sky130_fd_sc_hd__dlymetal6s2s_1
X_17251_ net2164 net190 net1799 net9219 VGND VGND VPWR VPWR _00349_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14463_ _06650_ VGND VGND VPWR VPWR _06651_ sky130_fd_sc_hd__buf_1
XFILLER_0_83_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13414_ _05686_ VGND VGND VPWR VPWR _05687_ sky130_fd_sc_hd__buf_1
X_16202_ _08185_ net981 VGND VGND VPWR VPWR _08267_ sky130_fd_sc_hd__xor2_2
X_17182_ net5997 net3344 _09096_ VGND VGND VPWR VPWR _09133_ sky130_fd_sc_hd__mux2_1
X_14394_ _06598_ matmul0.b_in\[1\] net900 VGND VGND VPWR VPWR _06599_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16133_ _08193_ _08198_ VGND VGND VPWR VPWR _08199_ sky130_fd_sc_hd__xnor2_1
X_13345_ net3679 net3675 net3682 net7923 _05617_ VGND VGND VPWR VPWR _05618_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_84_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16064_ net1093 _08130_ VGND VGND VPWR VPWR _08131_ sky130_fd_sc_hd__xnor2_1
X_13276_ _05463_ _05449_ _05448_ VGND VGND VPWR VPWR _05549_ sky130_fd_sc_hd__a21boi_1
Xwire5060 pid_q.mult0.b\[4\] VGND VGND VPWR VPWR net5060 sky130_fd_sc_hd__clkbuf_1
X_15015_ net6610 net7434 matmul0.matmul_stage_inst.a\[1\] net6582 VGND VGND VPWR VPWR
+ _07089_ sky130_fd_sc_hd__a22o_1
Xwire5071 net5067 VGND VGND VPWR VPWR net5071 sky130_fd_sc_hd__buf_1
Xwire5082 net5072 VGND VGND VPWR VPWR net5082 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5093 net5095 VGND VGND VPWR VPWR net5093 sky130_fd_sc_hd__clkbuf_1
Xwire4370 net4372 VGND VGND VPWR VPWR net4370 sky130_fd_sc_hd__buf_1
X_19823_ net6037 net1056 net3141 VGND VGND VPWR VPWR _11657_ sky130_fd_sc_hd__a21o_1
Xwire4381 net4382 VGND VGND VPWR VPWR net4381 sky130_fd_sc_hd__buf_1
Xwire4392 pid_d.prev_int\[0\] VGND VGND VPWR VPWR net4392 sky130_fd_sc_hd__buf_1
Xwire3680 net3681 VGND VGND VPWR VPWR net3680 sky130_fd_sc_hd__clkbuf_1
Xwire3691 net3692 VGND VGND VPWR VPWR net3691 sky130_fd_sc_hd__clkbuf_1
X_19754_ _11588_ net3129 net3146 VGND VGND VPWR VPWR _11589_ sky130_fd_sc_hd__a21o_1
X_16966_ _08844_ _08928_ net6519 VGND VGND VPWR VPWR _08929_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18705_ _10549_ _10550_ VGND VGND VPWR VPWR _10551_ sky130_fd_sc_hd__and2b_1
X_15917_ _07984_ _07985_ VGND VGND VPWR VPWR _07986_ sky130_fd_sc_hd__nand2_1
X_19685_ net6151 net3175 VGND VGND VPWR VPWR _11521_ sky130_fd_sc_hd__nor2_1
X_16897_ net6402 net6372 VGND VGND VPWR VPWR _08861_ sky130_fd_sc_hd__and2b_1
XFILLER_0_190_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18636_ net2127 _10482_ VGND VGND VPWR VPWR _10483_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_177_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15848_ _07730_ _07916_ _07917_ VGND VGND VPWR VPWR _07918_ sky130_fd_sc_hd__a21o_1
XFILLER_0_91_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18567_ net1071 _10380_ _10414_ VGND VGND VPWR VPWR _10415_ sky130_fd_sc_hd__o21ai_1
X_15779_ net3390 _07848_ VGND VGND VPWR VPWR _07849_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17518_ net6697 _09402_ _09403_ _09401_ VGND VGND VPWR VPWR _00403_ sky130_fd_sc_hd__a22o_1
X_18498_ _10284_ _10287_ VGND VGND VPWR VPWR _10347_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17449_ net3274 _09344_ net6656 VGND VGND VPWR VPWR _09345_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20460_ _12244_ net809 _12251_ VGND VGND VPWR VPWR _12252_ sky130_fd_sc_hd__o21a_1
XFILLER_0_171_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19119_ _10954_ _10885_ _10955_ VGND VGND VPWR VPWR _10956_ sky130_fd_sc_hd__mux2_1
X_20391_ net1399 _12188_ net8053 VGND VGND VPWR VPWR _12190_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22130_ net5779 net5799 VGND VGND VPWR VPWR _02136_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22061_ net1038 _02066_ VGND VGND VPWR VPWR _02068_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21012_ _00995_ _01004_ VGND VGND VPWR VPWR _01028_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25820_ clknet_leaf_31_clk _00693_ net8686 VGND VGND VPWR VPWR pid_q.prev_error\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1007 _05049_ VGND VGND VPWR VPWR net1007 sky130_fd_sc_hd__buf_1
Xwire1018 _03540_ VGND VGND VPWR VPWR net1018 sky130_fd_sc_hd__buf_1
XFILLER_0_96_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1029 net1030 VGND VGND VPWR VPWR net1029 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25751_ clknet_leaf_11_clk _00624_ net8602 VGND VGND VPWR VPWR pid_d.kp\[9\] sky130_fd_sc_hd__dfrtp_1
X_22963_ _02849_ VGND VGND VPWR VPWR _00648_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_94_clk clknet_4_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_94_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24702_ net8028 _04538_ VGND VGND VPWR VPWR _04539_ sky130_fd_sc_hd__xnor2_1
X_21914_ _01905_ VGND VGND VPWR VPWR _01922_ sky130_fd_sc_hd__inv_2
X_25682_ clknet_leaf_120_clk _00555_ net8395 VGND VGND VPWR VPWR pid_d.curr_error\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_22894_ net5976 _02787_ VGND VGND VPWR VPWR _02788_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_179_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24633_ net4894 net4871 _04428_ VGND VGND VPWR VPWR _04488_ sky130_fd_sc_hd__a21o_1
X_21845_ _01764_ _01765_ _01853_ VGND VGND VPWR VPWR _01854_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_194_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24564_ net4538 net3046 _04419_ VGND VGND VPWR VPWR _04420_ sky130_fd_sc_hd__or3_1
XFILLER_0_72_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21776_ _01690_ _01691_ _01692_ VGND VGND VPWR VPWR _01786_ sky130_fd_sc_hd__o21a_1
Xwire8603 net8604 VGND VGND VPWR VPWR net8603 sky130_fd_sc_hd__buf_1
Xwire8614 net8608 VGND VGND VPWR VPWR net8614 sky130_fd_sc_hd__buf_1
XFILLER_0_154_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8625 net8623 VGND VGND VPWR VPWR net8625 sky130_fd_sc_hd__clkbuf_2
X_23515_ _03309_ _03383_ VGND VGND VPWR VPWR _03384_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20727_ _12472_ _12491_ _12493_ _12495_ _12498_ VGND VGND VPWR VPWR _00518_ sky130_fd_sc_hd__a311o_1
XFILLER_0_65_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length5068 net5069 VGND VGND VPWR VPWR net5068 sky130_fd_sc_hd__clkbuf_1
Xwire8636 net8637 VGND VGND VPWR VPWR net8636 sky130_fd_sc_hd__clkbuf_1
X_24495_ net4871 _04349_ _04351_ VGND VGND VPWR VPWR _04352_ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7902 net7903 VGND VGND VPWR VPWR net7902 sky130_fd_sc_hd__clkbuf_1
Xwire8647 net8648 VGND VGND VPWR VPWR net8647 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_65_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7913 net7905 VGND VGND VPWR VPWR net7913 sky130_fd_sc_hd__clkbuf_1
Xwire304 _08377_ VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__clkbuf_1
Xwire315 net316 VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_190_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23446_ pid_q.curr_int\[0\] pid_q.prev_int\[0\] VGND VGND VPWR VPWR _03315_ sky130_fd_sc_hd__nand2_1
Xwire326 _05775_ VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__clkbuf_1
X_20658_ _12431_ _12434_ VGND VGND VPWR VPWR _12436_ sky130_fd_sc_hd__nor2_1
Xwire7946 net7947 VGND VGND VPWR VPWR net7946 sky130_fd_sc_hd__buf_1
Xwire337 _02260_ VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__buf_1
Xwire7957 net7958 VGND VGND VPWR VPWR net7957 sky130_fd_sc_hd__clkbuf_1
Xwire348 net349 VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__clkbuf_1
Xwire7968 net7969 VGND VGND VPWR VPWR net7968 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire359 net360 VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__buf_1
Xwire7979 pid_q.target\[11\] VGND VGND VPWR VPWR net7979 sky130_fd_sc_hd__clkbuf_1
Xmax_length3666 _06510_ VGND VGND VPWR VPWR net3666 sky130_fd_sc_hd__clkbuf_1
X_23377_ _03186_ _03187_ _03246_ VGND VGND VPWR VPWR _03247_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_162_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20589_ _12370_ _12371_ VGND VGND VPWR VPWR _12372_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13130_ _05398_ _05399_ net848 VGND VGND VPWR VPWR _05403_ sky130_fd_sc_hd__or3_1
X_25116_ net9209 net2393 net1993 pid_d.curr_int\[4\] VGND VGND VPWR VPWR _00797_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22328_ pid_d.curr_int\[13\] pid_d.prev_int\[13\] VGND VGND VPWR VPWR _02331_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length2976 _04956_ VGND VGND VPWR VPWR net2976 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25047_ _04795_ _04796_ VGND VGND VPWR VPWR _04798_ sky130_fd_sc_hd__or2_1
X_13061_ _05147_ _05150_ _05320_ _05333_ VGND VGND VPWR VPWR _05334_ sky130_fd_sc_hd__o31a_1
XFILLER_0_103_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22259_ pid_d.prev_error\[12\] pid_d.curr_error\[12\] VGND VGND VPWR VPWR _02263_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_178_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2220 _07896_ VGND VGND VPWR VPWR net2220 sky130_fd_sc_hd__buf_1
XFILLER_0_178_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2231 net2232 VGND VGND VPWR VPWR net2231 sky130_fd_sc_hd__clkbuf_1
X_16820_ _08800_ VGND VGND VPWR VPWR _00308_ sky130_fd_sc_hd__clkbuf_1
Xwire2242 _07231_ VGND VGND VPWR VPWR net2242 sky130_fd_sc_hd__buf_1
Xwire2253 net2254 VGND VGND VPWR VPWR net2253 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2264 _06519_ VGND VGND VPWR VPWR net2264 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2275 net2276 VGND VGND VPWR VPWR net2275 sky130_fd_sc_hd__clkbuf_1
Xwire1530 net1531 VGND VGND VPWR VPWR net1530 sky130_fd_sc_hd__clkbuf_2
Xwire2286 _06502_ VGND VGND VPWR VPWR net2286 sky130_fd_sc_hd__clkbuf_1
Xwire1541 _07380_ VGND VGND VPWR VPWR net1541 sky130_fd_sc_hd__clkbuf_1
X_16751_ _08764_ VGND VGND VPWR VPWR _00275_ sky130_fd_sc_hd__clkbuf_1
X_13963_ net7703 net1324 VGND VGND VPWR VPWR _06228_ sky130_fd_sc_hd__nand2_1
Xwire2297 net2298 VGND VGND VPWR VPWR net2297 sky130_fd_sc_hd__buf_1
Xwire1552 net1553 VGND VGND VPWR VPWR net1552 sky130_fd_sc_hd__buf_1
Xwire1563 _05909_ VGND VGND VPWR VPWR net1563 sky130_fd_sc_hd__clkbuf_2
Xwire1574 _05577_ VGND VGND VPWR VPWR net1574 sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_85_clk clknet_4_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_85_clk sky130_fd_sc_hd__clkbuf_16
Xwire1585 _05387_ VGND VGND VPWR VPWR net1585 sky130_fd_sc_hd__buf_1
X_15702_ net1535 _07772_ VGND VGND VPWR VPWR _07773_ sky130_fd_sc_hd__xnor2_1
Xwire1596 _05132_ VGND VGND VPWR VPWR net1596 sky130_fd_sc_hd__buf_1
X_12914_ net2310 net1955 VGND VGND VPWR VPWR _05187_ sky130_fd_sc_hd__and2_1
X_19470_ net960 net1420 VGND VGND VPWR VPWR _11307_ sky130_fd_sc_hd__nand2_1
X_13894_ _06125_ _06135_ VGND VGND VPWR VPWR _06160_ sky130_fd_sc_hd__nand2_1
X_16682_ _08712_ _08713_ VGND VGND VPWR VPWR _08714_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_186_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18421_ net6825 net6773 net6798 _10270_ VGND VGND VPWR VPWR _10271_ sky130_fd_sc_hd__a31o_1
X_12845_ net1006 net1005 VGND VGND VPWR VPWR _05118_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15633_ net1857 _07608_ VGND VGND VPWR VPWR _07705_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18352_ net716 net715 _10196_ _10198_ _10202_ VGND VGND VPWR VPWR _10203_ sky130_fd_sc_hd__o32a_1
XFILLER_0_96_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12776_ _04908_ _04914_ _05048_ VGND VGND VPWR VPWR _05049_ sky130_fd_sc_hd__o21ai_1
X_15564_ _07569_ _07635_ VGND VGND VPWR VPWR _07637_ sky130_fd_sc_hd__nor2_1
Xmax_length6270 net6271 VGND VGND VPWR VPWR net6270 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17303_ _09205_ net7630 VGND VGND VPWR VPWR _09217_ sky130_fd_sc_hd__nand2_1
Xmax_length6281 net6275 VGND VGND VPWR VPWR net6281 sky130_fd_sc_hd__clkbuf_1
X_14515_ net5262 _06693_ VGND VGND VPWR VPWR _06696_ sky130_fd_sc_hd__nand2_1
Xmax_length6292 net6293 VGND VGND VPWR VPWR net6292 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_126_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15495_ net1274 net1875 _07566_ _07567_ VGND VGND VPWR VPWR _07568_ sky130_fd_sc_hd__a22o_1
X_18283_ _10057_ _10071_ VGND VGND VPWR VPWR _10134_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17234_ _09170_ _09181_ VGND VGND VPWR VPWR _09182_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14446_ _06638_ matmul0.b_in\[13\] net994 VGND VGND VPWR VPWR _06639_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14377_ net7217 net1296 net2893 net5328 _06585_ VGND VGND VPWR VPWR _06586_ sky130_fd_sc_hd__a221o_1
X_17165_ _09102_ net527 _09117_ VGND VGND VPWR VPWR _09118_ sky130_fd_sc_hd__o21ai_1
Xwire860 _01416_ VGND VGND VPWR VPWR net860 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_107_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire871 _11240_ VGND VGND VPWR VPWR net871 sky130_fd_sc_hd__clkbuf_1
Xwire882 _08386_ VGND VGND VPWR VPWR net882 sky130_fd_sc_hd__dlymetal6s2s_1
X_13328_ _05599_ _05600_ VGND VGND VPWR VPWR _05601_ sky130_fd_sc_hd__and2_1
Xwire893 net894 VGND VGND VPWR VPWR net893 sky130_fd_sc_hd__buf_1
XFILLER_0_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16116_ net1512 _08181_ VGND VGND VPWR VPWR _08182_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17096_ net2595 net3363 _08971_ VGND VGND VPWR VPWR _09053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13259_ svm0.vC\[14\] net2992 VGND VGND VPWR VPWR _05532_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16047_ net2646 net2633 VGND VGND VPWR VPWR _08114_ sky130_fd_sc_hd__nor2_2
XFILLER_0_0_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19806_ net6215 net6157 VGND VGND VPWR VPWR _11640_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17998_ net7083 net7038 VGND VGND VPWR VPWR _09849_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_193_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19737_ net3879 net6026 VGND VGND VPWR VPWR _11572_ sky130_fd_sc_hd__nand2_1
X_16949_ net7125 _08910_ _08912_ VGND VGND VPWR VPWR _00325_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_76_clk clknet_4_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_76_clk sky130_fd_sc_hd__clkbuf_16
X_19668_ _11409_ _11503_ _11501_ VGND VGND VPWR VPWR _11504_ sky130_fd_sc_hd__nor3_1
XFILLER_0_35_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18619_ _10431_ _10465_ VGND VGND VPWR VPWR _10466_ sky130_fd_sc_hd__nor2_1
X_19599_ net6063 net6027 VGND VGND VPWR VPWR _11436_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21630_ net4357 _01640_ _01641_ VGND VGND VPWR VPWR _01642_ sky130_fd_sc_hd__and3_1
XFILLER_0_158_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21561_ net5782 net5501 VGND VGND VPWR VPWR _01573_ sky130_fd_sc_hd__nand2_1
Xwire7209 net7211 VGND VGND VPWR VPWR net7209 sky130_fd_sc_hd__buf_1
X_23300_ _03152_ _03169_ _03168_ _03149_ VGND VGND VPWR VPWR _03170_ sky130_fd_sc_hd__o2bb2a_1
X_20512_ _12295_ net3846 _12297_ net3845 net4060 net3334 VGND VGND VPWR VPWR _12299_
+ sky130_fd_sc_hd__mux4_1
X_24280_ _04060_ _04065_ _04058_ VGND VGND VPWR VPWR _04140_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21492_ net1728 _01390_ _01504_ VGND VGND VPWR VPWR _01505_ sky130_fd_sc_hd__a21o_1
Xwire6508 net6509 VGND VGND VPWR VPWR net6508 sky130_fd_sc_hd__buf_1
Xwire6519 net6520 VGND VGND VPWR VPWR net6519 sky130_fd_sc_hd__buf_1
XFILLER_0_160_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23231_ _03011_ _03012_ _03010_ VGND VGND VPWR VPWR _03101_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_127_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20443_ _12226_ _12236_ _08857_ VGND VGND VPWR VPWR _12237_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5807 net5808 VGND VGND VPWR VPWR net5807 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire5818 net5816 VGND VGND VPWR VPWR net5818 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5829 pid_d.mult0.b\[6\] VGND VGND VPWR VPWR net5829 sky130_fd_sc_hd__buf_1
X_23162_ _03028_ _03029_ _03031_ VGND VGND VPWR VPWR _03032_ sky130_fd_sc_hd__o21ai_2
X_20374_ net950 _12172_ VGND VGND VPWR VPWR _12173_ sky130_fd_sc_hd__xnor2_1
Xmax_length1549 net1550 VGND VGND VPWR VPWR net1549 sky130_fd_sc_hd__clkbuf_1
X_22113_ net2062 net945 VGND VGND VPWR VPWR _02119_ sky130_fd_sc_hd__and2_1
X_23093_ _02946_ _02962_ VGND VGND VPWR VPWR _02963_ sky130_fd_sc_hd__xnor2_2
X_22044_ _02036_ _02050_ VGND VGND VPWR VPWR _02051_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_167_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25803_ clknet_leaf_30_clk _00676_ net8675 VGND VGND VPWR VPWR pid_q.curr_int\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23995_ net7526 _03775_ net333 net7466 net854 VGND VGND VPWR VPWR _03859_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_67_clk clknet_4_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_67_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_173_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_170_Right_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25734_ clknet_leaf_12_clk _00607_ net8605 VGND VGND VPWR VPWR pid_d.ki\[8\] sky130_fd_sc_hd__dfrtp_1
X_22946_ net551 net549 _02324_ VGND VGND VPWR VPWR _02834_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_97_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25665_ clknet_leaf_121_clk _00538_ net8396 VGND VGND VPWR VPWR pid_d.prev_error\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_22877_ _02770_ _02771_ VGND VGND VPWR VPWR _02773_ sky130_fd_sc_hd__or2_1
X_12630_ net7881 net1356 VGND VGND VPWR VPWR _04903_ sky130_fd_sc_hd__nand2_1
X_24616_ net2018 _04470_ VGND VGND VPWR VPWR _04471_ sky130_fd_sc_hd__nand2_1
X_21828_ net5750 net5479 VGND VGND VPWR VPWR _01837_ sky130_fd_sc_hd__nand2_2
X_25596_ clknet_leaf_106_clk _00469_ net8355 VGND VGND VPWR VPWR cordic0.slte0.opB\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8338 net8538 VGND VGND VPWR VPWR net8338 sky130_fd_sc_hd__buf_1
Xwire8400 net8398 VGND VGND VPWR VPWR net8400 sky130_fd_sc_hd__buf_1
X_24547_ net1649 _04354_ VGND VGND VPWR VPWR _04403_ sky130_fd_sc_hd__and2_1
Xwire8411 net8412 VGND VGND VPWR VPWR net8411 sky130_fd_sc_hd__clkbuf_1
X_21759_ _01666_ _01668_ VGND VGND VPWR VPWR _01769_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8422 net8420 VGND VGND VPWR VPWR net8422 sky130_fd_sc_hd__clkbuf_2
Xwire8444 net8441 VGND VGND VPWR VPWR net8444 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire7710 net7705 VGND VGND VPWR VPWR net7710 sky130_fd_sc_hd__buf_1
X_14300_ net1549 VGND VGND VPWR VPWR _06522_ sky130_fd_sc_hd__buf_1
X_15280_ net3486 net3441 VGND VGND VPWR VPWR _07354_ sky130_fd_sc_hd__nor2_1
Xfanout6914 cordic0.vec\[1\]\[10\] VGND VGND VPWR VPWR net6914 sky130_fd_sc_hd__clkbuf_2
Xwire7721 net7717 VGND VGND VPWR VPWR net7721 sky130_fd_sc_hd__buf_1
X_24478_ net5175 pid_q.prev_int\[12\] VGND VGND VPWR VPWR _04335_ sky130_fd_sc_hd__and2_1
Xfanout6936 net6939 VGND VGND VPWR VPWR net6936 sky130_fd_sc_hd__buf_1
XFILLER_0_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7743 net7741 VGND VGND VPWR VPWR net7743 sky130_fd_sc_hd__buf_1
XFILLER_0_18_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14231_ _06481_ _06488_ VGND VGND VPWR VPWR _06489_ sky130_fd_sc_hd__xnor2_1
Xwire7754 svm0.periodTop\[8\] VGND VGND VPWR VPWR net7754 sky130_fd_sc_hd__buf_1
X_23429_ _03262_ _03298_ VGND VGND VPWR VPWR _03299_ sky130_fd_sc_hd__xnor2_1
Xwire7765 net7766 VGND VGND VPWR VPWR net7765 sky130_fd_sc_hd__buf_1
XFILLER_0_150_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3452 _07230_ VGND VGND VPWR VPWR net3452 sky130_fd_sc_hd__clkbuf_1
Xwire156 _06479_ VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__buf_1
XFILLER_0_34_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3463 _07189_ VGND VGND VPWR VPWR net3463 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire167 net168 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__buf_1
Xwire7787 net7788 VGND VGND VPWR VPWR net7787 sky130_fd_sc_hd__buf_1
Xwire178 _02618_ VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_1
Xmax_length3474 net3475 VGND VGND VPWR VPWR net3474 sky130_fd_sc_hd__buf_1
Xwire189 net190 VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__buf_1
Xwire7798 net7791 VGND VGND VPWR VPWR net7798 sky130_fd_sc_hd__clkbuf_1
X_14162_ net217 _06422_ VGND VGND VPWR VPWR _06423_ sky130_fd_sc_hd__nand2_1
Xmax_length3496 net3501 VGND VGND VPWR VPWR net3496 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13113_ _05384_ _05385_ VGND VGND VPWR VPWR _05386_ sky130_fd_sc_hd__xor2_1
XFILLER_0_42_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2795 net2796 VGND VGND VPWR VPWR net2795 sky130_fd_sc_hd__buf_1
X_14093_ _06323_ _06355_ VGND VGND VPWR VPWR _06356_ sky130_fd_sc_hd__xnor2_1
X_18970_ net2530 net3214 VGND VGND VPWR VPWR _10807_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13044_ _05306_ _05310_ _05316_ VGND VGND VPWR VPWR _05317_ sky130_fd_sc_hd__a21o_1
X_17921_ _09665_ _09669_ net3248 VGND VGND VPWR VPWR _09772_ sky130_fd_sc_hd__o21a_1
X_17852_ net7130 net7146 VGND VGND VPWR VPWR _09703_ sky130_fd_sc_hd__and2b_1
Xwire2061 _01798_ VGND VGND VPWR VPWR net2061 sky130_fd_sc_hd__clkbuf_1
X_16803_ _08791_ VGND VGND VPWR VPWR _00300_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2083 _12300_ VGND VGND VPWR VPWR net2083 sky130_fd_sc_hd__clkbuf_1
X_17783_ net7023 net7030 VGND VGND VPWR VPWR _09634_ sky130_fd_sc_hd__and2_1
XFILLER_0_191_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_58_clk clknet_4_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_16
X_14995_ net1898 _07060_ net1896 VGND VGND VPWR VPWR _07069_ sky130_fd_sc_hd__o21bai_1
Xwire2094 _11802_ VGND VGND VPWR VPWR net2094 sky130_fd_sc_hd__clkbuf_1
Xwire1360 net1361 VGND VGND VPWR VPWR net1360 sky130_fd_sc_hd__buf_1
Xwire1371 _04530_ VGND VGND VPWR VPWR net1371 sky130_fd_sc_hd__buf_1
X_19522_ _11291_ VGND VGND VPWR VPWR _11359_ sky130_fd_sc_hd__inv_2
X_16734_ _08755_ VGND VGND VPWR VPWR _00267_ sky130_fd_sc_hd__clkbuf_1
X_13946_ _06137_ _06140_ net530 VGND VGND VPWR VPWR _06212_ sky130_fd_sc_hd__o21ai_1
Xwire1382 net1383 VGND VGND VPWR VPWR net1382 sky130_fd_sc_hd__clkbuf_1
Xwire1393 _00858_ VGND VGND VPWR VPWR net1393 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_72_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19453_ net6119 net6086 VGND VGND VPWR VPWR _11290_ sky130_fd_sc_hd__nand2_1
XFILLER_0_159_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16665_ _08698_ _08694_ matmul0.matmul_stage_inst.mult2\[6\] VGND VGND VPWR VPWR
+ _08699_ sky130_fd_sc_hd__o21ba_1
X_13877_ _06081_ _06143_ VGND VGND VPWR VPWR _06144_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18404_ _10252_ _10254_ VGND VGND VPWR VPWR _10255_ sky130_fd_sc_hd__xnor2_1
X_15616_ net4074 net4069 net4075 VGND VGND VPWR VPWR _07688_ sky130_fd_sc_hd__a21o_1
XFILLER_0_186_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12828_ net1336 _05100_ VGND VGND VPWR VPWR _05101_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_22_Left_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19384_ net2509 _11157_ VGND VGND VPWR VPWR _11221_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16596_ _08646_ VGND VGND VPWR VPWR _08647_ sky130_fd_sc_hd__clkbuf_1
X_18335_ _10157_ _10185_ VGND VGND VPWR VPWR _10186_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_167_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15547_ net3502 net2820 _07526_ _07016_ net3412 VGND VGND VPWR VPWR _07620_ sky130_fd_sc_hd__a32o_1
X_12759_ _05002_ _05031_ VGND VGND VPWR VPWR _05032_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18266_ net3233 _10048_ VGND VGND VPWR VPWR _10117_ sky130_fd_sc_hd__nand2_1
X_15478_ _07402_ net1274 _07550_ _07551_ VGND VGND VPWR VPWR _07552_ sky130_fd_sc_hd__o31a_1
XFILLER_0_112_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17217_ _09163_ _09165_ VGND VGND VPWR VPWR _09166_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14429_ matmul0.beta_pass\[9\] net1293 net2889 net4425 _06625_ VGND VGND VPWR VPWR
+ _06626_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18197_ net3997 net3952 net6996 VGND VGND VPWR VPWR _10048_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_13_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17148_ net1801 _09101_ VGND VGND VPWR VPWR _09102_ sky130_fd_sc_hd__xnor2_2
Xwire690 net691 VGND VGND VPWR VPWR net690 sky130_fd_sc_hd__buf_1
XFILLER_0_188_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_31_Left_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17079_ net1805 _08975_ net2172 net1802 VGND VGND VPWR VPWR _09037_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20090_ _11873_ VGND VGND VPWR VPWR _11919_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length8408 net8405 VGND VGND VPWR VPWR net8408 sky130_fd_sc_hd__clkbuf_1
X_22800_ pid_d.kp\[12\] _02686_ _02694_ VGND VGND VPWR VPWR _02708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23780_ net4810 _03499_ net3049 VGND VGND VPWR VPWR _03646_ sky130_fd_sc_hd__a21oi_1
X_20992_ _00952_ _00955_ net3111 VGND VGND VPWR VPWR _01008_ sky130_fd_sc_hd__a21o_1
X_22731_ _02665_ VGND VGND VPWR VPWR _00600_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_40_Left_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25450_ clknet_leaf_112_clk _00333_ net8341 VGND VGND VPWR VPWR cordic0.vec\[1\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22662_ pid_d.mult0.b\[14\] net3775 VGND VGND VPWR VPWR _02616_ sky130_fd_sc_hd__or2_1
X_24401_ pid_q.prev_int\[11\] _04189_ net5177 VGND VGND VPWR VPWR _04259_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21613_ _01619_ _01624_ VGND VGND VPWR VPWR _01625_ sky130_fd_sc_hd__nand2_1
X_25381_ clknet_leaf_74_clk _00264_ net8466 VGND VGND VPWR VPWR matmul0.b\[0\] sky130_fd_sc_hd__dfrtp_1
X_22593_ net7287 _02566_ VGND VGND VPWR VPWR _02570_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24332_ _04189_ _04190_ VGND VGND VPWR VPWR _04191_ sky130_fd_sc_hd__xnor2_1
Xwire7006 net7007 VGND VGND VPWR VPWR net7006 sky130_fd_sc_hd__buf_1
XFILLER_0_35_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21544_ _01448_ _01450_ _01555_ VGND VGND VPWR VPWR _01556_ sky130_fd_sc_hd__a21oi_2
Xwire7017 net7015 VGND VGND VPWR VPWR net7017 sky130_fd_sc_hd__buf_1
Xwire7028 net7029 VGND VGND VPWR VPWR net7028 sky130_fd_sc_hd__buf_1
XFILLER_0_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24263_ net1159 _04086_ _04122_ VGND VGND VPWR VPWR _04123_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6327 net6328 VGND VGND VPWR VPWR net6327 sky130_fd_sc_hd__buf_1
X_21475_ _01373_ _01375_ _01374_ VGND VGND VPWR VPWR _01488_ sky130_fd_sc_hd__o21a_1
XFILLER_0_172_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6338 net6340 VGND VGND VPWR VPWR net6338 sky130_fd_sc_hd__buf_1
Xwire5604 net5605 VGND VGND VPWR VPWR net5604 sky130_fd_sc_hd__clkbuf_1
Xwire6349 net6350 VGND VGND VPWR VPWR net6349 sky130_fd_sc_hd__clkbuf_1
X_23214_ net5065 _03080_ VGND VGND VPWR VPWR _03084_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5615 net5616 VGND VGND VPWR VPWR net5615 sky130_fd_sc_hd__buf_1
XFILLER_0_161_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length1313 _05730_ VGND VGND VPWR VPWR net1313 sky130_fd_sc_hd__buf_1
XFILLER_0_133_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20426_ net1832 _12221_ net8045 VGND VGND VPWR VPWR _12222_ sky130_fd_sc_hd__o21ai_1
X_24194_ net4580 net4853 VGND VGND VPWR VPWR _04055_ sky130_fd_sc_hd__nand2_1
Xwire5626 net5625 VGND VGND VPWR VPWR net5626 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_30_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5637 net5638 VGND VGND VPWR VPWR net5637 sky130_fd_sc_hd__buf_1
Xwire5648 net5649 VGND VGND VPWR VPWR net5648 sky130_fd_sc_hd__clkbuf_1
Xwire4914 net4915 VGND VGND VPWR VPWR net4914 sky130_fd_sc_hd__clkbuf_1
Xwire5659 net5660 VGND VGND VPWR VPWR net5659 sky130_fd_sc_hd__clkbuf_1
X_23145_ net5084 net4716 VGND VGND VPWR VPWR _03015_ sky130_fd_sc_hd__nand2_2
Xwire4925 net4923 VGND VGND VPWR VPWR net4925 sky130_fd_sc_hd__clkbuf_1
Xwire4936 net4939 VGND VGND VPWR VPWR net4936 sky130_fd_sc_hd__clkbuf_1
X_20357_ net6515 _12157_ _12096_ VGND VGND VPWR VPWR _12158_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4947 net4945 VGND VGND VPWR VPWR net4947 sky130_fd_sc_hd__clkbuf_1
Xwire4958 net4959 VGND VGND VPWR VPWR net4958 sky130_fd_sc_hd__clkbuf_1
Xwire4969 net4973 VGND VGND VPWR VPWR net4969 sky130_fd_sc_hd__buf_1
X_23076_ net2432 _02945_ VGND VGND VPWR VPWR _02946_ sky130_fd_sc_hd__xnor2_2
X_20288_ net3314 _12091_ _12092_ _12093_ net6479 VGND VGND VPWR VPWR _12094_ sky130_fd_sc_hd__o221a_1
X_22027_ _02030_ _02033_ VGND VGND VPWR VPWR _02034_ sky130_fd_sc_hd__xnor2_2
Xhold20 matmul0.matmul_stage_inst.b\[15\] VGND VGND VPWR VPWR net8973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 matmul0.matmul_stage_inst.a\[14\] VGND VGND VPWR VPWR net8984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 svm0.vC\[13\] VGND VGND VPWR VPWR net8995 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 cordic0.cos\[10\] VGND VGND VPWR VPWR net9006 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold64 matmul0.matmul_stage_inst.c\[4\] VGND VGND VPWR VPWR net9017 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 pid_d.curr_error\[3\] VGND VGND VPWR VPWR net9028 sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ net3677 _05947_ VGND VGND VPWR VPWR _06068_ sky130_fd_sc_hd__nor2_1
Xhold86 matmul0.matmul_stage_inst.b\[9\] VGND VGND VPWR VPWR net9039 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 pid_d.curr_error\[2\] VGND VGND VPWR VPWR net9050 sky130_fd_sc_hd__dlygate4sd3_1
X_14780_ net4223 _06858_ VGND VGND VPWR VPWR _06904_ sky130_fd_sc_hd__and2_1
X_23978_ _03839_ _03841_ VGND VGND VPWR VPWR _03842_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13731_ _05927_ _05929_ _05996_ _05999_ VGND VGND VPWR VPWR _06000_ sky130_fd_sc_hd__a211o_1
X_25717_ clknet_leaf_9_clk _00590_ net8555 VGND VGND VPWR VPWR pid_d.mult0.a\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_22929_ _02819_ VGND VGND VPWR VPWR _00644_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16450_ net2634 net2641 VGND VGND VPWR VPWR _08511_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13662_ _05930_ _05931_ VGND VGND VPWR VPWR _05932_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25648_ clknet_leaf_122_clk _00521_ net8407 VGND VGND VPWR VPWR pid_d.curr_int\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15401_ _07405_ _07408_ _07474_ _07072_ VGND VGND VPWR VPWR _07475_ sky130_fd_sc_hd__o2bb2a_1
X_12613_ net4315 VGND VGND VPWR VPWR _04887_ sky130_fd_sc_hd__inv_2
X_13593_ _05840_ net783 _05841_ VGND VGND VPWR VPWR _05863_ sky130_fd_sc_hd__o21ai_1
X_16381_ net1250 _08442_ net2815 VGND VGND VPWR VPWR _08443_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_137_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25579_ clknet_leaf_98_clk _00452_ net8384 VGND VGND VPWR VPWR cordic0.sin\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_18120_ _09960_ _09970_ VGND VGND VPWR VPWR _09971_ sky130_fd_sc_hd__xor2_1
Xwire8230 net8231 VGND VGND VPWR VPWR net8230 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15332_ _07124_ net1117 VGND VGND VPWR VPWR _07406_ sky130_fd_sc_hd__or2_1
Xwire8241 net8242 VGND VGND VPWR VPWR net8241 sky130_fd_sc_hd__clkbuf_1
Xwire8252 net27 VGND VGND VPWR VPWR net8252 sky130_fd_sc_hd__clkbuf_1
Xwire8263 net8264 VGND VGND VPWR VPWR net8263 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8274 net8275 VGND VGND VPWR VPWR net8274 sky130_fd_sc_hd__clkbuf_1
Xwire8285 net8286 VGND VGND VPWR VPWR net8285 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18051_ net7078 net7112 VGND VGND VPWR VPWR _09902_ sky130_fd_sc_hd__xnor2_2
Xwire7540 net7541 VGND VGND VPWR VPWR net7540 sky130_fd_sc_hd__clkbuf_1
Xwire8296 net8297 VGND VGND VPWR VPWR net8296 sky130_fd_sc_hd__clkbuf_1
X_15263_ _07259_ _07257_ _07235_ _07255_ VGND VGND VPWR VPWR _07337_ sky130_fd_sc_hd__o211a_1
Xfanout6755 net6767 VGND VGND VPWR VPWR net6755 sky130_fd_sc_hd__buf_1
XFILLER_0_81_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7551 net7552 VGND VGND VPWR VPWR net7551 sky130_fd_sc_hd__clkbuf_1
Xwire7562 net7563 VGND VGND VPWR VPWR net7562 sky130_fd_sc_hd__clkbuf_1
Xwire7573 matmul0.b_in\[3\] VGND VGND VPWR VPWR net7573 sky130_fd_sc_hd__clkbuf_1
Xwire7584 matmul0.a_in\[14\] VGND VGND VPWR VPWR net7584 sky130_fd_sc_hd__buf_1
X_17002_ net1833 _08963_ net8042 VGND VGND VPWR VPWR _08964_ sky130_fd_sc_hd__o21ai_1
Xfanout6777 net6782 VGND VGND VPWR VPWR net6777 sky130_fd_sc_hd__clkbuf_1
X_14214_ net1121 _06471_ net1304 net7629 VGND VGND VPWR VPWR _06473_ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout6788 net6806 VGND VGND VPWR VPWR net6788 sky130_fd_sc_hd__buf_1
Xmax_length3282 net3283 VGND VGND VPWR VPWR net3282 sky130_fd_sc_hd__clkbuf_2
X_15194_ net3554 VGND VGND VPWR VPWR _07268_ sky130_fd_sc_hd__clkbuf_1
Xwire7595 net7596 VGND VGND VPWR VPWR net7595 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length2570 net2571 VGND VGND VPWR VPWR net2570 sky130_fd_sc_hd__buf_1
X_14145_ net7647 net1120 VGND VGND VPWR VPWR _06406_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length2592 net2593 VGND VGND VPWR VPWR net2592 sky130_fd_sc_hd__buf_1
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14076_ net7646 _06336_ _06337_ net7633 _06338_ VGND VGND VPWR VPWR _06339_ sky130_fd_sc_hd__o221a_1
X_18953_ net6085 VGND VGND VPWR VPWR _10790_ sky130_fd_sc_hd__inv_2
X_13027_ _05160_ _05161_ VGND VGND VPWR VPWR _05300_ sky130_fd_sc_hd__nand2_1
X_17904_ _09753_ _09754_ VGND VGND VPWR VPWR _09755_ sky130_fd_sc_hd__nand2b_1
X_18884_ _10723_ net873 VGND VGND VPWR VPWR _10726_ sky130_fd_sc_hd__xnor2_1
X_17835_ net7019 _09602_ _09684_ _09051_ _09685_ VGND VGND VPWR VPWR _09686_ sky130_fd_sc_hd__o221a_2
X_17766_ net7118 VGND VGND VPWR VPWR _09617_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14978_ _07050_ _07051_ VGND VGND VPWR VPWR _07052_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1190 _11638_ VGND VGND VPWR VPWR net1190 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19505_ net1751 _11341_ VGND VGND VPWR VPWR _11342_ sky130_fd_sc_hd__xnor2_2
X_16717_ _08742_ _08743_ VGND VGND VPWR VPWR _08744_ sky130_fd_sc_hd__xnor2_1
X_13929_ _06193_ _06194_ VGND VGND VPWR VPWR _06195_ sky130_fd_sc_hd__xnor2_1
X_17697_ _09204_ _09573_ VGND VGND VPWR VPWR _00413_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19436_ net3870 _10971_ _11272_ VGND VGND VPWR VPWR _11273_ sky130_fd_sc_hd__o21a_1
X_16648_ net7328 net1838 net6551 VGND VGND VPWR VPWR _08685_ sky130_fd_sc_hd__mux2_1
XFILLER_0_187_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19367_ net1753 _11089_ VGND VGND VPWR VPWR _11204_ sky130_fd_sc_hd__xor2_1
X_16579_ matmul0.matmul_stage_inst.mult2\[0\] net494 net2620 VGND VGND VPWR VPWR _08637_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18318_ net6842 net6789 VGND VGND VPWR VPWR _10169_ sky130_fd_sc_hd__xnor2_2
Xfanout8680 net8685 VGND VGND VPWR VPWR net8680 sky130_fd_sc_hd__buf_1
XFILLER_0_128_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19298_ net2512 _11134_ VGND VGND VPWR VPWR _11135_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18249_ _10095_ _10096_ _10098_ net2544 VGND VGND VPWR VPWR _10100_ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21260_ net1730 _01274_ VGND VGND VPWR VPWR _01275_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_163_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20211_ net8120 net8119 VGND VGND VPWR VPWR _12034_ sky130_fd_sc_hd__nor2_1
X_21191_ _01142_ _01140_ VGND VGND VPWR VPWR _01207_ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3509 net3510 VGND VGND VPWR VPWR net3509 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20142_ _11968_ _11949_ net2493 VGND VGND VPWR VPWR _11969_ sky130_fd_sc_hd__a21o_1
Xwire2819 net2820 VGND VGND VPWR VPWR net2819 sky130_fd_sc_hd__buf_1
XFILLER_0_148_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24950_ _04727_ VGND VGND VPWR VPWR _00757_ sky130_fd_sc_hd__clkbuf_1
X_20073_ net1404 _11898_ _11901_ net6002 VGND VGND VPWR VPWR _11902_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23901_ _03764_ _03765_ VGND VGND VPWR VPWR _03766_ sky130_fd_sc_hd__nand2_1
X_24881_ _04678_ net4602 net1996 VGND VGND VPWR VPWR _04679_ sky130_fd_sc_hd__mux2_1
X_23832_ _03695_ _03696_ VGND VGND VPWR VPWR _03697_ sky130_fd_sc_hd__xnor2_1
X_23763_ _03620_ _03628_ VGND VGND VPWR VPWR _03629_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_196_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20975_ net5631 net5821 _00989_ _00990_ VGND VGND VPWR VPWR _00991_ sky130_fd_sc_hd__a31o_1
XFILLER_0_164_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25502_ clknet_leaf_41_clk _00382_ net8772 VGND VGND VPWR VPWR svm0.delta\[7\] sky130_fd_sc_hd__dfrtp_1
X_22714_ net5373 net3705 _04886_ net5372 VGND VGND VPWR VPWR _02651_ sky130_fd_sc_hd__a22o_1
X_23694_ _03451_ _03461_ _03560_ VGND VGND VPWR VPWR _03561_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25433_ clknet_leaf_97_clk _00316_ net8400 VGND VGND VPWR VPWR matmul0.sin\[6\] sky130_fd_sc_hd__dfrtp_1
X_22645_ net5840 net3082 _02607_ net946 net8893 VGND VGND VPWR VPWR _00572_ sky130_fd_sc_hd__o221a_1
XFILLER_0_36_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25364_ clknet_leaf_72_clk _00247_ net8477 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult2\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout6007 net6011 VGND VGND VPWR VPWR net6007 sky130_fd_sc_hd__buf_1
X_22576_ net9028 net2043 net3093 net2458 VGND VGND VPWR VPWR _00554_ sky130_fd_sc_hd__a22o_1
Xfanout6018 net6035 VGND VGND VPWR VPWR net6018 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24315_ pid_q.curr_int\[10\] pid_q.prev_int\[10\] VGND VGND VPWR VPWR _04175_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6102 net6103 VGND VGND VPWR VPWR net6102 sky130_fd_sc_hd__buf_1
X_21527_ net4384 _01440_ net416 net4320 net1723 VGND VGND VPWR VPWR _01540_ sky130_fd_sc_hd__a221o_1
XFILLER_0_173_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25295_ clknet_leaf_89_clk _00178_ net8420 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.d\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire6124 net6125 VGND VGND VPWR VPWR net6124 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24246_ _04105_ _04106_ VGND VGND VPWR VPWR _04107_ sky130_fd_sc_hd__or2_1
Xwire5401 net5402 VGND VGND VPWR VPWR net5401 sky130_fd_sc_hd__buf_1
Xwire5412 net5409 VGND VGND VPWR VPWR net5412 sky130_fd_sc_hd__buf_1
X_21458_ _01343_ _01345_ _01344_ VGND VGND VPWR VPWR _01471_ sky130_fd_sc_hd__o21a_1
Xwire6157 net6156 VGND VGND VPWR VPWR net6157 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_16_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5434 net5435 VGND VGND VPWR VPWR net5434 sky130_fd_sc_hd__buf_1
XFILLER_0_160_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6179 net6177 VGND VGND VPWR VPWR net6179 sky130_fd_sc_hd__buf_1
XFILLER_0_120_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20409_ net811 _12197_ VGND VGND VPWR VPWR _12206_ sky130_fd_sc_hd__and2b_1
Xwire5445 net5446 VGND VGND VPWR VPWR net5445 sky130_fd_sc_hd__clkbuf_1
Xwire4711 pid_q.mult0.a\[4\] VGND VGND VPWR VPWR net4711 sky130_fd_sc_hd__clkbuf_1
X_24177_ pid_q.curr_int\[8\] VGND VGND VPWR VPWR _04038_ sky130_fd_sc_hd__inv_2
Xwire5456 net5457 VGND VGND VPWR VPWR net5456 sky130_fd_sc_hd__buf_1
Xmax_length1154 _05026_ VGND VGND VPWR VPWR net1154 sky130_fd_sc_hd__clkbuf_1
Xwire5467 net5468 VGND VGND VPWR VPWR net5467 sky130_fd_sc_hd__clkbuf_1
X_21389_ net5651 _01402_ VGND VGND VPWR VPWR _01403_ sky130_fd_sc_hd__xnor2_2
Xwire4733 net4724 VGND VGND VPWR VPWR net4733 sky130_fd_sc_hd__buf_1
Xwire5489 pid_d.mult0.a\[10\] VGND VGND VPWR VPWR net5489 sky130_fd_sc_hd__buf_1
XFILLER_0_120_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length1176 _01642_ VGND VGND VPWR VPWR net1176 sky130_fd_sc_hd__clkbuf_1
Xwire4755 net4753 VGND VGND VPWR VPWR net4755 sky130_fd_sc_hd__buf_1
X_23128_ _02996_ _02997_ VGND VGND VPWR VPWR _02998_ sky130_fd_sc_hd__nand2_1
Xwire4766 net4767 VGND VGND VPWR VPWR net4766 sky130_fd_sc_hd__clkbuf_1
Xwire4777 net4778 VGND VGND VPWR VPWR net4777 sky130_fd_sc_hd__buf_1
Xwire4788 net4789 VGND VGND VPWR VPWR net4788 sky130_fd_sc_hd__buf_1
Xwire4799 net4800 VGND VGND VPWR VPWR net4799 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23059_ _02924_ _02927_ _02928_ VGND VGND VPWR VPWR _02929_ sky130_fd_sc_hd__mux2_1
X_15950_ net984 _08017_ _07959_ VGND VGND VPWR VPWR _08018_ sky130_fd_sc_hd__o21ai_2
Xinput110 pid_d_data[7] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_1
Xinput121 pid_q_addr[1] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_1
Xinput132 pid_q_data[11] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_1
X_14901_ net6542 net6586 net7398 VGND VGND VPWR VPWR _06975_ sky130_fd_sc_hd__o21a_1
Xinput143 pid_q_data[7] VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_1
X_15881_ net2700 _07929_ net3396 _07842_ VGND VGND VPWR VPWR _07950_ sky130_fd_sc_hd__o211a_1
X_17620_ net4018 svm0.tB\[3\] _09500_ VGND VGND VPWR VPWR _09501_ sky130_fd_sc_hd__a21oi_1
X_14832_ matmul0.a\[5\] matmul0.matmul_stage_inst.e\[5\] net3610 VGND VGND VPWR VPWR
+ _06933_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17551_ net4006 svm0.tC\[7\] svm0.tC\[5\] _09230_ _09432_ VGND VGND VPWR VPWR _09433_
+ sky130_fd_sc_hd__o221a_1
Xmax_length8761 net8762 VGND VGND VPWR VPWR net8761 sky130_fd_sc_hd__buf_1
XFILLER_0_187_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14763_ net7152 _06842_ net3615 VGND VGND VPWR VPWR _06892_ sky130_fd_sc_hd__o21a_1
X_16502_ net2750 _08560_ _08561_ net2783 net2638 VGND VGND VPWR VPWR _08562_ sky130_fd_sc_hd__o221a_1
X_13714_ _05979_ net727 VGND VGND VPWR VPWR _05983_ sky130_fd_sc_hd__xnor2_1
X_17482_ svm0.delta\[7\] _09372_ VGND VGND VPWR VPWR _09373_ sky130_fd_sc_hd__xnor2_1
X_14694_ net7153 _06840_ VGND VGND VPWR VPWR _06841_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19221_ net6240 net2519 _11057_ VGND VGND VPWR VPWR _11058_ sky130_fd_sc_hd__o21a_1
X_16433_ net303 _08482_ VGND VGND VPWR VPWR _08494_ sky130_fd_sc_hd__nand2_1
X_13645_ _05821_ _05831_ _05830_ VGND VGND VPWR VPWR _05915_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19152_ net6290 net6334 VGND VGND VPWR VPWR _10989_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16364_ _08424_ net773 VGND VGND VPWR VPWR _08427_ sky130_fd_sc_hd__or2_2
X_13576_ net577 _05846_ VGND VGND VPWR VPWR _05847_ sky130_fd_sc_hd__xnor2_1
X_18103_ net2549 _09952_ _09953_ VGND VGND VPWR VPWR _09954_ sky130_fd_sc_hd__a21o_1
Xwire8060 net8061 VGND VGND VPWR VPWR net8060 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8071 net8072 VGND VGND VPWR VPWR net8071 sky130_fd_sc_hd__clkbuf_1
X_15315_ net3461 net3555 VGND VGND VPWR VPWR _07389_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8082 net8083 VGND VGND VPWR VPWR net8082 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19083_ net3211 _10829_ net3192 VGND VGND VPWR VPWR _10920_ sky130_fd_sc_hd__mux2_1
X_16295_ _08308_ _08358_ VGND VGND VPWR VPWR _08359_ sky130_fd_sc_hd__xnor2_2
Xwire8093 net8094 VGND VGND VPWR VPWR net8093 sky130_fd_sc_hd__clkbuf_1
X_18034_ _09862_ _09851_ VGND VGND VPWR VPWR _09885_ sky130_fd_sc_hd__xnor2_2
Xwire7370 net7371 VGND VGND VPWR VPWR net7370 sky130_fd_sc_hd__clkbuf_1
X_15246_ net3594 net3592 net4127 net4125 VGND VGND VPWR VPWR _07320_ sky130_fd_sc_hd__o22a_1
Xwire7381 matmul0.matmul_stage_inst.f\[12\] VGND VGND VPWR VPWR net7381 sky130_fd_sc_hd__clkbuf_1
Xfanout5840 pid_d.mult0.b\[5\] VGND VGND VPWR VPWR net5840 sky130_fd_sc_hd__buf_1
XFILLER_0_169_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7392 net7393 VGND VGND VPWR VPWR net7392 sky130_fd_sc_hd__clkbuf_1
Xwire6680 net6681 VGND VGND VPWR VPWR net6680 sky130_fd_sc_hd__clkbuf_1
Xwire6691 net6692 VGND VGND VPWR VPWR net6691 sky130_fd_sc_hd__buf_1
XFILLER_0_2_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15177_ net1883 _07250_ VGND VGND VPWR VPWR _07251_ sky130_fd_sc_hd__nand2_1
Xfanout5895 pid_d.mult0.b\[3\] VGND VGND VPWR VPWR net5895 sky130_fd_sc_hd__buf_1
XFILLER_0_111_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14128_ net1597 net1125 _06174_ _06221_ VGND VGND VPWR VPWR _06390_ sky130_fd_sc_hd__or4b_1
Xwire5990 net5988 VGND VGND VPWR VPWR net5990 sky130_fd_sc_hd__buf_1
X_19985_ _11814_ _11815_ VGND VGND VPWR VPWR _11816_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_105_Left_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14059_ _06290_ _06309_ _06246_ VGND VGND VPWR VPWR _06322_ sky130_fd_sc_hd__a21bo_1
X_18936_ net6863 net6878 net6813 net6779 VGND VGND VPWR VPWR _10775_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18867_ net6832 net3224 VGND VGND VPWR VPWR _10709_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17818_ net3260 _09667_ _09668_ VGND VGND VPWR VPWR _09669_ sky130_fd_sc_hd__a21o_1
X_18798_ net2588 _10218_ _10546_ VGND VGND VPWR VPWR _10642_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17749_ _09599_ VGND VGND VPWR VPWR _09600_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20760_ _12509_ _12510_ VGND VGND VPWR VPWR _12531_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_114_Left_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19419_ net6317 _10797_ VGND VGND VPWR VPWR _11256_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20691_ _12463_ _12465_ VGND VGND VPWR VPWR _12466_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_92_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22430_ net5723 net5749 net5389 net5711 VGND VGND VPWR VPWR _02432_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22361_ _02360_ _02363_ VGND VGND VPWR VPWR _02364_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24100_ net5149 net4483 net3749 _03886_ VGND VGND VPWR VPWR _03962_ sky130_fd_sc_hd__and4_1
X_21312_ _00877_ _00933_ _01326_ VGND VGND VPWR VPWR _01327_ sky130_fd_sc_hd__o21ai_1
X_25080_ _04824_ _04825_ VGND VGND VPWR VPWR _04826_ sky130_fd_sc_hd__or2_1
X_22292_ _02290_ _02295_ VGND VGND VPWR VPWR _02296_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24031_ net4552 net4911 VGND VGND VPWR VPWR _03894_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4007 _09376_ VGND VGND VPWR VPWR net4007 sky130_fd_sc_hd__buf_1
XFILLER_0_103_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21243_ net5844 net5495 VGND VGND VPWR VPWR _01258_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4029 net4030 VGND VGND VPWR VPWR net4029 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_123_Left_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire3306 net3312 VGND VGND VPWR VPWR net3306 sky130_fd_sc_hd__clkbuf_1
X_21174_ net3839 _01189_ VGND VGND VPWR VPWR _01190_ sky130_fd_sc_hd__xnor2_1
Xwire3317 net3318 VGND VGND VPWR VPWR net3317 sky130_fd_sc_hd__buf_1
Xwire3328 net3329 VGND VGND VPWR VPWR net3328 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_102_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3339 net3340 VGND VGND VPWR VPWR net3339 sky130_fd_sc_hd__buf_1
Xwire2605 _08950_ VGND VGND VPWR VPWR net2605 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20125_ net5999 _11900_ _11952_ _11897_ VGND VGND VPWR VPWR _11953_ sky130_fd_sc_hd__a2bb2o_1
Xwire2616 net2617 VGND VGND VPWR VPWR net2616 sky130_fd_sc_hd__buf_1
Xwire2638 net2639 VGND VGND VPWR VPWR net2638 sky130_fd_sc_hd__buf_1
Xwire1904 net1905 VGND VGND VPWR VPWR net1904 sky130_fd_sc_hd__clkbuf_1
Xwire2649 net2650 VGND VGND VPWR VPWR net2649 sky130_fd_sc_hd__buf_1
Xwire1915 net1916 VGND VGND VPWR VPWR net1915 sky130_fd_sc_hd__buf_1
X_24933_ net8868 net143 VGND VGND VPWR VPWR _04716_ sky130_fd_sc_hd__and2b_1
Xwire1926 net1927 VGND VGND VPWR VPWR net1926 sky130_fd_sc_hd__dlymetal6s2s_1
X_20056_ _11880_ _11884_ net6058 VGND VGND VPWR VPWR _11885_ sky130_fd_sc_hd__o21a_1
Xwire1937 _05642_ VGND VGND VPWR VPWR net1937 sky130_fd_sc_hd__buf_1
Xwire1948 _05287_ VGND VGND VPWR VPWR net1948 sky130_fd_sc_hd__buf_1
XFILLER_0_175_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1959 _05056_ VGND VGND VPWR VPWR net1959 sky130_fd_sc_hd__buf_1
X_24864_ pid_q.ki\[3\] net2398 net3008 pid_q.kp\[3\] VGND VGND VPWR VPWR _04667_ sky130_fd_sc_hd__a22o_1
X_23815_ _03652_ _03654_ VGND VGND VPWR VPWR _03680_ sky130_fd_sc_hd__or2_1
XFILLER_0_169_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24795_ _04614_ _04613_ VGND VGND VPWR VPWR _04620_ sky130_fd_sc_hd__nand2_1
Xmax_length6611 net6612 VGND VGND VPWR VPWR net6611 sky130_fd_sc_hd__buf_1
XFILLER_0_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23746_ net1662 _03610_ VGND VGND VPWR VPWR _03612_ sky130_fd_sc_hd__nand2_1
X_20958_ net5635 net5793 _00959_ _00973_ VGND VGND VPWR VPWR _00974_ sky130_fd_sc_hd__a31o_1
XFILLER_0_36_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length5910 net5911 VGND VGND VPWR VPWR net5910 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length5932 net5933 VGND VGND VPWR VPWR net5932 sky130_fd_sc_hd__clkbuf_1
X_23677_ _03441_ _03443_ _03439_ VGND VGND VPWR VPWR _03544_ sky130_fd_sc_hd__o21a_1
X_20889_ _00901_ _00902_ _00904_ VGND VGND VPWR VPWR _00905_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_193_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13430_ _05701_ _05702_ VGND VGND VPWR VPWR _05703_ sky130_fd_sc_hd__xnor2_1
X_25416_ clknet_leaf_89_clk _00299_ net8422 VGND VGND VPWR VPWR matmul0.cos\[3\] sky130_fd_sc_hd__dfrtp_1
X_22628_ _02597_ VGND VGND VPWR VPWR _00565_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length5987 pid_d.curr_int\[0\] VGND VGND VPWR VPWR net5987 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_192_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13361_ net731 _05633_ VGND VGND VPWR VPWR _05634_ sky130_fd_sc_hd__xor2_1
X_22559_ _04873_ _02542_ VGND VGND VPWR VPWR _02543_ sky130_fd_sc_hd__or2_1
X_25347_ clknet_leaf_72_clk _00230_ net8477 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout5103 pid_q.mult0.b\[2\] VGND VGND VPWR VPWR net5103 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length832 _06652_ VGND VGND VPWR VPWR net832 sky130_fd_sc_hd__clkbuf_2
X_15100_ net4190 net4184 net3583 net3581 VGND VGND VPWR VPWR _07174_ sky130_fd_sc_hd__o22a_1
X_13292_ _05482_ _05564_ VGND VGND VPWR VPWR _05565_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16080_ _08140_ _08146_ VGND VGND VPWR VPWR _08147_ sky130_fd_sc_hd__xnor2_2
X_25278_ clknet_leaf_70_clk _00161_ net8447 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.c\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire5220 net5221 VGND VGND VPWR VPWR net5220 sky130_fd_sc_hd__buf_1
Xwire5231 net5232 VGND VGND VPWR VPWR net5231 sky130_fd_sc_hd__clkbuf_1
X_15031_ _07084_ _07104_ VGND VGND VPWR VPWR _07105_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24229_ net4590 net4604 net3053 VGND VGND VPWR VPWR _04090_ sky130_fd_sc_hd__and3_1
Xmax_length898 _06606_ VGND VGND VPWR VPWR net898 sky130_fd_sc_hd__buf_1
Xwire5242 matmul0.beta_pass\[9\] VGND VGND VPWR VPWR net5242 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5264 matmul0.beta_pass\[6\] VGND VGND VPWR VPWR net5264 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5275 net5277 VGND VGND VPWR VPWR net5275 sky130_fd_sc_hd__clkbuf_1
Xwire4541 net4542 VGND VGND VPWR VPWR net4541 sky130_fd_sc_hd__clkbuf_1
Xwire5286 net5287 VGND VGND VPWR VPWR net5286 sky130_fd_sc_hd__buf_1
Xwire4552 net4553 VGND VGND VPWR VPWR net4552 sky130_fd_sc_hd__clkbuf_1
Xwire5297 net5298 VGND VGND VPWR VPWR net5297 sky130_fd_sc_hd__buf_1
Xwire4563 net4564 VGND VGND VPWR VPWR net4563 sky130_fd_sc_hd__buf_1
XFILLER_0_43_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4574 net4570 VGND VGND VPWR VPWR net4574 sky130_fd_sc_hd__buf_1
XFILLER_0_102_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3840 net3841 VGND VGND VPWR VPWR net3840 sky130_fd_sc_hd__buf_1
Xwire4585 net4586 VGND VGND VPWR VPWR net4585 sky130_fd_sc_hd__clkbuf_1
X_19770_ _11601_ _11604_ VGND VGND VPWR VPWR _11605_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4596 net4599 VGND VGND VPWR VPWR net4596 sky130_fd_sc_hd__clkbuf_1
Xwire3851 _12267_ VGND VGND VPWR VPWR net3851 sky130_fd_sc_hd__clkbuf_1
X_16982_ net6520 net4052 net6460 VGND VGND VPWR VPWR _08944_ sky130_fd_sc_hd__a21o_1
Xwire3862 net3863 VGND VGND VPWR VPWR net3862 sky130_fd_sc_hd__buf_1
Xwire3884 _10943_ VGND VGND VPWR VPWR net3884 sky130_fd_sc_hd__clkbuf_1
X_18721_ net421 _10566_ VGND VGND VPWR VPWR _10567_ sky130_fd_sc_hd__xor2_1
Xwire3895 _10878_ VGND VGND VPWR VPWR net3895 sky130_fd_sc_hd__buf_1
XFILLER_0_3_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15933_ _07999_ _08001_ VGND VGND VPWR VPWR _08002_ sky130_fd_sc_hd__xnor2_1
X_18652_ _10493_ _10498_ VGND VGND VPWR VPWR _10499_ sky130_fd_sc_hd__xnor2_1
X_15864_ _07932_ VGND VGND VPWR VPWR _07933_ sky130_fd_sc_hd__clkbuf_1
X_17603_ net4015 svm0.tB\[10\] VGND VGND VPWR VPWR _09484_ sky130_fd_sc_hd__nor2_1
X_14815_ net9044 net2877 net2854 _06924_ VGND VGND VPWR VPWR _00179_ sky130_fd_sc_hd__o22a_1
XFILLER_0_189_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18583_ net7000 net6895 VGND VGND VPWR VPWR _10431_ sky130_fd_sc_hd__xnor2_2
X_15795_ net3458 _07864_ VGND VGND VPWR VPWR _07865_ sky130_fd_sc_hd__nor2_1
XFILLER_0_192_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length8580 net8575 VGND VGND VPWR VPWR net8580 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_98_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17534_ svm0.delta\[15\] _09416_ VGND VGND VPWR VPWR _09417_ sky130_fd_sc_hd__xnor2_1
X_14746_ _06835_ _06878_ net7448 VGND VGND VPWR VPWR _06879_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17465_ svm0.counter\[4\] VGND VGND VPWR VPWR _09358_ sky130_fd_sc_hd__inv_2
XFILLER_0_168_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14677_ net4223 _06827_ VGND VGND VPWR VPWR _06828_ sky130_fd_sc_hd__or2_1
X_19204_ net3183 _11029_ VGND VGND VPWR VPWR _11041_ sky130_fd_sc_hd__and2_1
X_16416_ _08421_ _08413_ _08477_ VGND VGND VPWR VPWR _08478_ sky130_fd_sc_hd__a21o_1
X_13628_ net7686 net2331 net2326 VGND VGND VPWR VPWR _05898_ sky130_fd_sc_hd__and3_1
X_17396_ _09299_ net614 _09300_ _09302_ VGND VGND VPWR VPWR _00382_ sky130_fd_sc_hd__a31o_1
XFILLER_0_27_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout7050 net7055 VGND VGND VPWR VPWR net7050 sky130_fd_sc_hd__buf_1
X_19135_ net6175 net6151 VGND VGND VPWR VPWR _10972_ sky130_fd_sc_hd__and2b_1
XFILLER_0_13_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16347_ net1250 _08409_ VGND VGND VPWR VPWR _08410_ sky130_fd_sc_hd__xnor2_1
X_13559_ _05822_ _05829_ VGND VGND VPWR VPWR _05830_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19066_ _10877_ _10883_ VGND VGND VPWR VPWR _10903_ sky130_fd_sc_hd__xor2_1
XFILLER_0_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16278_ net2840 net2644 _08341_ VGND VGND VPWR VPWR _08342_ sky130_fd_sc_hd__a21o_1
X_18017_ net2551 _09866_ _09867_ VGND VGND VPWR VPWR _09868_ sky130_fd_sc_hd__a21oi_1
X_15229_ net4169 net4164 net4127 net4124 VGND VGND VPWR VPWR _07303_ sky130_fd_sc_hd__o22a_1
XFILLER_0_1_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout4980 net5005 VGND VGND VPWR VPWR net4980 sky130_fd_sc_hd__buf_1
X_19968_ _10788_ _11798_ net6081 VGND VGND VPWR VPWR _11799_ sky130_fd_sc_hd__mux2_1
X_18919_ _10752_ _10753_ _10756_ _10758_ VGND VGND VPWR VPWR _10759_ sky130_fd_sc_hd__o211a_1
X_19899_ _11667_ net708 _11715_ VGND VGND VPWR VPWR _11731_ sky130_fd_sc_hd__nand3_1
X_21930_ _01932_ _01937_ VGND VGND VPWR VPWR _01938_ sky130_fd_sc_hd__xor2_1
XFILLER_0_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21861_ net5394 _01782_ _01869_ net5857 VGND VGND VPWR VPWR _01870_ sky130_fd_sc_hd__o22a_1
XFILLER_0_145_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23600_ _03463_ _03467_ VGND VGND VPWR VPWR _03468_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20812_ net5810 net5524 VGND VGND VPWR VPWR _00828_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24580_ _04433_ _04434_ _04430_ VGND VGND VPWR VPWR _04436_ sky130_fd_sc_hd__a21o_1
X_21792_ _01744_ _01801_ VGND VGND VPWR VPWR _01802_ sky130_fd_sc_hd__xnor2_2
Xmax_length5206 net5207 VGND VGND VPWR VPWR net5206 sky130_fd_sc_hd__buf_1
X_23531_ _03330_ _03331_ _03398_ VGND VGND VPWR VPWR _03399_ sky130_fd_sc_hd__a21bo_1
X_20743_ net5914 net5473 VGND VGND VPWR VPWR _12514_ sky130_fd_sc_hd__nand2_2
Xmax_length4505 net4506 VGND VGND VPWR VPWR net4505 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8818 net8819 VGND VGND VPWR VPWR net8818 sky130_fd_sc_hd__clkbuf_1
Xwire8829 net8830 VGND VGND VPWR VPWR net8829 sky130_fd_sc_hd__clkbuf_1
X_23462_ net4532 net5128 VGND VGND VPWR VPWR _03331_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20674_ _12448_ _12449_ _12450_ net6091 VGND VGND VPWR VPWR _00513_ sky130_fd_sc_hd__o22a_1
XFILLER_0_174_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire508 _04653_ VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22413_ _02383_ _02413_ _02414_ VGND VGND VPWR VPWR _02415_ sky130_fd_sc_hd__a21o_1
Xwire519 _02512_ VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__clkbuf_1
X_25201_ clknet_leaf_82_clk _00090_ net8496 VGND VGND VPWR VPWR matmul0.b_in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_23393_ _03216_ _03227_ net1674 VGND VGND VPWR VPWR _03263_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25132_ clknet_leaf_52_clk _00021_ net8803 VGND VGND VPWR VPWR svm0.tC\[4\] sky130_fd_sc_hd__dfrtp_1
X_22344_ _02291_ _02292_ _02346_ VGND VGND VPWR VPWR _02347_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_115_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25063_ net3732 _04806_ _04810_ VGND VGND VPWR VPWR _04811_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22275_ _02242_ _02243_ _02278_ VGND VGND VPWR VPWR _02279_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24014_ _03807_ _03809_ _03808_ VGND VGND VPWR VPWR _03877_ sky130_fd_sc_hd__o21ai_1
Xhold150 pid_q.target\[8\] VGND VGND VPWR VPWR net9103 sky130_fd_sc_hd__dlygate4sd3_1
X_21226_ _00935_ _01241_ VGND VGND VPWR VPWR _01242_ sky130_fd_sc_hd__xor2_1
Xwire3103 net3104 VGND VGND VPWR VPWR net3103 sky130_fd_sc_hd__clkbuf_2
Xwire3114 net3116 VGND VGND VPWR VPWR net3114 sky130_fd_sc_hd__clkbuf_1
Xhold161 pid_d.prev_error\[7\] VGND VGND VPWR VPWR net9114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 pid_q.prev_int\[13\] VGND VGND VPWR VPWR net9125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 svm0.tA\[5\] VGND VGND VPWR VPWR net9136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 svm0.tC\[3\] VGND VGND VPWR VPWR net9147 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3136 _11447_ VGND VGND VPWR VPWR net3136 sky130_fd_sc_hd__clkbuf_2
Xwire2402 net2403 VGND VGND VPWR VPWR net2402 sky130_fd_sc_hd__clkbuf_1
X_21157_ net5611 net5948 net5928 net5629 VGND VGND VPWR VPWR _01173_ sky130_fd_sc_hd__a22o_1
Xwire3147 net3148 VGND VGND VPWR VPWR net3147 sky130_fd_sc_hd__buf_1
Xwire2413 _03501_ VGND VGND VPWR VPWR net2413 sky130_fd_sc_hd__buf_1
Xwire3158 net3159 VGND VGND VPWR VPWR net3158 sky130_fd_sc_hd__clkbuf_2
Xwire2424 net2425 VGND VGND VPWR VPWR net2424 sky130_fd_sc_hd__clkbuf_2
Xwire3169 net3170 VGND VGND VPWR VPWR net3169 sky130_fd_sc_hd__buf_1
Xwire2435 net2436 VGND VGND VPWR VPWR net2435 sky130_fd_sc_hd__clkbuf_1
X_20108_ net6001 _11890_ net6063 net3140 VGND VGND VPWR VPWR _11936_ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2446 _02624_ VGND VGND VPWR VPWR net2446 sky130_fd_sc_hd__buf_1
Xwire1701 _02522_ VGND VGND VPWR VPWR net1701 sky130_fd_sc_hd__buf_1
Xwire1712 _02059_ VGND VGND VPWR VPWR net1712 sky130_fd_sc_hd__buf_1
X_21088_ net5642 net5793 _01100_ _01102_ _01103_ VGND VGND VPWR VPWR _01104_ sky130_fd_sc_hd__a311o_1
Xwire2457 net2458 VGND VGND VPWR VPWR net2457 sky130_fd_sc_hd__clkbuf_1
Xwire2468 net2469 VGND VGND VPWR VPWR net2468 sky130_fd_sc_hd__buf_1
Xwire1723 _01539_ VGND VGND VPWR VPWR net1723 sky130_fd_sc_hd__clkbuf_1
Xwire2479 _01306_ VGND VGND VPWR VPWR net2479 sky130_fd_sc_hd__buf_1
Xwire1734 _00958_ VGND VGND VPWR VPWR net1734 sky130_fd_sc_hd__clkbuf_2
Xwire1745 net1746 VGND VGND VPWR VPWR net1745 sky130_fd_sc_hd__clkbuf_2
X_24916_ pid_q.ki\[1\] _04704_ _04702_ VGND VGND VPWR VPWR _04705_ sky130_fd_sc_hd__mux2_1
X_12930_ _05199_ _05202_ VGND VGND VPWR VPWR _05203_ sky130_fd_sc_hd__xnor2_2
X_20039_ _11806_ _11868_ VGND VGND VPWR VPWR _11869_ sky130_fd_sc_hd__xnor2_1
Xwire1756 _10932_ VGND VGND VPWR VPWR net1756 sky130_fd_sc_hd__buf_1
X_25896_ clknet_leaf_15_clk _00769_ net8622 VGND VGND VPWR VPWR pid_q.kp\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1778 _09981_ VGND VGND VPWR VPWR net1778 sky130_fd_sc_hd__clkbuf_1
Xwire1789 net1790 VGND VGND VPWR VPWR net1789 sky130_fd_sc_hd__buf_1
X_24847_ net4841 net2007 _04540_ net258 VGND VGND VPWR VPWR _00725_ sky130_fd_sc_hd__a22o_1
X_12861_ net2334 net2329 VGND VGND VPWR VPWR _05134_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length7120 net7121 VGND VGND VPWR VPWR net7120 sky130_fd_sc_hd__buf_1
X_14600_ net9084 net892 _06773_ net2887 VGND VGND VPWR VPWR _00115_ sky130_fd_sc_hd__a22o_1
X_15580_ net2833 net3489 net2677 _07580_ VGND VGND VPWR VPWR _07652_ sky130_fd_sc_hd__a31o_1
X_24778_ net7980 _04598_ VGND VGND VPWR VPWR _04605_ sky130_fd_sc_hd__nand2_1
X_12792_ net1959 _04965_ _05064_ net7935 _05060_ VGND VGND VPWR VPWR _05065_ sky130_fd_sc_hd__o221a_1
XFILLER_0_157_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14531_ _06709_ VGND VGND VPWR VPWR _06710_ sky130_fd_sc_hd__clkbuf_2
X_23729_ _03512_ _03514_ _03594_ VGND VGND VPWR VPWR _03595_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_194_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17250_ net2164 net221 net1799 net9090 VGND VGND VPWR VPWR _00348_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14462_ _06513_ _06541_ VGND VGND VPWR VPWR _06650_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16201_ _08261_ _08265_ VGND VGND VPWR VPWR _08266_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_181_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13413_ net2949 net1941 VGND VGND VPWR VPWR _05686_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17181_ net6850 _09131_ _09132_ VGND VGND VPWR VPWR _00337_ sky130_fd_sc_hd__a21bo_1
X_14393_ net5306 net1297 net2894 net4467 _06597_ VGND VGND VPWR VPWR _06598_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16132_ _08196_ _08197_ VGND VGND VPWR VPWR _08198_ sky130_fd_sc_hd__and2_1
X_13344_ net2294 VGND VGND VPWR VPWR _05617_ sky130_fd_sc_hd__buf_1
XFILLER_0_134_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16063_ _08127_ net1092 VGND VGND VPWR VPWR _08130_ sky130_fd_sc_hd__xor2_1
X_13275_ _05545_ _05546_ _05538_ VGND VGND VPWR VPWR _05548_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_51_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5050 net5056 VGND VGND VPWR VPWR net5050 sky130_fd_sc_hd__clkbuf_1
X_15014_ net6629 matmul0.matmul_stage_inst.d\[1\] net7418 net6534 VGND VGND VPWR VPWR
+ _07088_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_184_Right_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5094 net5096 VGND VGND VPWR VPWR net5094 sky130_fd_sc_hd__clkbuf_1
Xwire4360 net4359 VGND VGND VPWR VPWR net4360 sky130_fd_sc_hd__buf_1
Xwire4371 net4372 VGND VGND VPWR VPWR net4371 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19822_ _11574_ net958 net956 VGND VGND VPWR VPWR _11656_ sky130_fd_sc_hd__o21ai_2
Xwire4382 net4379 VGND VGND VPWR VPWR net4382 sky130_fd_sc_hd__buf_1
XFILLER_0_120_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4393 pid_q.out\[15\] VGND VGND VPWR VPWR net4393 sky130_fd_sc_hd__buf_1
Xwire3670 net3671 VGND VGND VPWR VPWR net3670 sky130_fd_sc_hd__buf_1
Xwire3681 _05615_ VGND VGND VPWR VPWR net3681 sky130_fd_sc_hd__clkbuf_1
X_16965_ net6195 net6167 net6504 VGND VGND VPWR VPWR _08928_ sky130_fd_sc_hd__mux2_1
X_19753_ net6046 net4045 VGND VGND VPWR VPWR _11588_ sky130_fd_sc_hd__nand2_2
XFILLER_0_194_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3692 _05022_ VGND VGND VPWR VPWR net3692 sky130_fd_sc_hd__clkbuf_1
Xwire2980 _04929_ VGND VGND VPWR VPWR net2980 sky130_fd_sc_hd__clkbuf_1
X_15916_ net884 _07983_ VGND VGND VPWR VPWR _07985_ sky130_fd_sc_hd__nand2_1
X_18704_ _10545_ _10548_ VGND VGND VPWR VPWR _10550_ sky130_fd_sc_hd__nand2_1
X_19684_ _11046_ net6257 VGND VGND VPWR VPWR _11520_ sky130_fd_sc_hd__nor2_1
Xwire2991 _04890_ VGND VGND VPWR VPWR net2991 sky130_fd_sc_hd__buf_1
X_16896_ net6369 _08858_ _08859_ VGND VGND VPWR VPWR _08860_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_188_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18635_ net6813 net6779 net6795 VGND VGND VPWR VPWR _10482_ sky130_fd_sc_hd__o21ai_1
X_15847_ _07819_ _07915_ VGND VGND VPWR VPWR _07917_ sky130_fd_sc_hd__nor2_1
XFILLER_0_189_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18566_ net1071 _10380_ net961 VGND VGND VPWR VPWR _10414_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15778_ net2650 _07761_ VGND VGND VPWR VPWR _07848_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17517_ net6697 _09272_ VGND VGND VPWR VPWR _09403_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14729_ net8980 net2872 _06865_ VGND VGND VPWR VPWR _00152_ sky130_fd_sc_hd__a21o_1
X_18497_ net874 _10345_ VGND VGND VPWR VPWR _10346_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17448_ net6743 _09343_ VGND VGND VPWR VPWR _09344_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17379_ net2572 _09288_ VGND VGND VPWR VPWR _09289_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19118_ net6245 net3896 VGND VGND VPWR VPWR _10955_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20390_ cordic0.slte0.opA\[8\] net1399 VGND VGND VPWR VPWR _12189_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19049_ _10877_ _10883_ _10885_ VGND VGND VPWR VPWR _10886_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22060_ net1038 _02066_ VGND VGND VPWR VPWR _02067_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_151_Right_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21011_ net862 _01025_ _01026_ VGND VGND VPWR VPWR _01027_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_49_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1008 _04948_ VGND VGND VPWR VPWR net1008 sky130_fd_sc_hd__buf_2
Xwire1019 _03511_ VGND VGND VPWR VPWR net1019 sky130_fd_sc_hd__buf_1
XFILLER_0_156_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25750_ clknet_leaf_12_clk _00623_ net8605 VGND VGND VPWR VPWR pid_d.kp\[8\] sky130_fd_sc_hd__dfrtp_1
X_22962_ matmul0.beta_pass\[0\] net4063 net6572 VGND VGND VPWR VPWR _02849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24701_ net1621 _04537_ VGND VGND VPWR VPWR _04538_ sky130_fd_sc_hd__nand2_1
X_21913_ _01919_ _01920_ VGND VGND VPWR VPWR _01921_ sky130_fd_sc_hd__xnor2_1
X_25681_ clknet_leaf_0_clk _00554_ net8409 VGND VGND VPWR VPWR pid_d.curr_error\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_22893_ _02017_ _02779_ _02786_ VGND VGND VPWR VPWR _02787_ sky130_fd_sc_hd__a21o_1
X_24632_ _04477_ _04486_ VGND VGND VPWR VPWR _04487_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_179_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21844_ _01764_ _01765_ _01763_ VGND VGND VPWR VPWR _01853_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_194_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24563_ _04343_ _04345_ VGND VGND VPWR VPWR _04419_ sky130_fd_sc_hd__nor2_1
X_21775_ _01781_ _01784_ VGND VGND VPWR VPWR _01785_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8604 net8602 VGND VGND VPWR VPWR net8604 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_19_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23514_ _03318_ _03382_ VGND VGND VPWR VPWR _03383_ sky130_fd_sc_hd__xnor2_1
X_20726_ net2284 _12497_ net4246 net5994 VGND VGND VPWR VPWR _12498_ sky130_fd_sc_hd__a2bb2o_1
Xwire8626 net8623 VGND VGND VPWR VPWR net8626 sky130_fd_sc_hd__buf_1
XFILLER_0_33_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8637 net8638 VGND VGND VPWR VPWR net8637 sky130_fd_sc_hd__clkbuf_1
X_24494_ net4919 _04350_ net4491 VGND VGND VPWR VPWR _04351_ sky130_fd_sc_hd__o21ai_1
Xwire7903 net7904 VGND VGND VPWR VPWR net7903 sky130_fd_sc_hd__clkbuf_1
Xwire8648 net8645 VGND VGND VPWR VPWR net8648 sky130_fd_sc_hd__buf_1
XFILLER_0_19_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4335 net4336 VGND VGND VPWR VPWR net4335 sky130_fd_sc_hd__buf_1
XFILLER_0_163_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8659 net8660 VGND VGND VPWR VPWR net8659 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_52_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length3612 _06928_ VGND VGND VPWR VPWR net3612 sky130_fd_sc_hd__buf_1
Xwire305 net306 VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__clkbuf_1
Xwire7925 net7918 VGND VGND VPWR VPWR net7925 sky130_fd_sc_hd__buf_1
X_23445_ pid_q.curr_int\[0\] net3061 net2028 _03314_ VGND VGND VPWR VPWR _00665_ sky130_fd_sc_hd__a22o_1
X_20657_ _12431_ _12434_ VGND VGND VPWR VPWR _12435_ sky130_fd_sc_hd__and2_1
Xwire316 net317 VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire327 _04655_ VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__clkbuf_1
Xwire7936 net7937 VGND VGND VPWR VPWR net7936 sky130_fd_sc_hd__buf_1
Xmax_length3623 _06823_ VGND VGND VPWR VPWR net3623 sky130_fd_sc_hd__clkbuf_1
Xwire7947 net7948 VGND VGND VPWR VPWR net7947 sky130_fd_sc_hd__buf_1
Xwire338 net339 VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__clkbuf_1
Xwire7958 net7959 VGND VGND VPWR VPWR net7958 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire349 _02007_ VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__clkbuf_1
Xmax_length2922 net2923 VGND VGND VPWR VPWR net2922 sky130_fd_sc_hd__clkbuf_1
X_23376_ _03186_ _03187_ _03188_ VGND VGND VPWR VPWR _03246_ sky130_fd_sc_hd__o21a_1
Xwire7969 net7970 VGND VGND VPWR VPWR net7969 sky130_fd_sc_hd__clkbuf_1
Xmax_length3667 net3668 VGND VGND VPWR VPWR net3667 sky130_fd_sc_hd__buf_1
X_20588_ _12369_ _12362_ VGND VGND VPWR VPWR _12371_ sky130_fd_sc_hd__or2b_1
X_25115_ pid_d.prev_int\[3\] net2392 net1992 pid_d.curr_int\[3\] VGND VGND VPWR VPWR
+ _00796_ sky130_fd_sc_hd__a22o_1
X_22327_ pid_d.curr_int\[13\] pid_d.prev_int\[13\] VGND VGND VPWR VPWR _02330_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13060_ _05151_ _05328_ _05144_ _05332_ VGND VGND VPWR VPWR _05333_ sky130_fd_sc_hd__a211o_1
X_25046_ _04795_ _04796_ VGND VGND VPWR VPWR _04797_ sky130_fd_sc_hd__nand2_1
X_22258_ pid_d.prev_error\[12\] pid_d.curr_error\[12\] VGND VGND VPWR VPWR _02262_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21209_ _01223_ net1734 VGND VGND VPWR VPWR _01225_ sky130_fd_sc_hd__nor2_1
X_22189_ _02159_ net859 _02160_ _02162_ VGND VGND VPWR VPWR _02194_ sky130_fd_sc_hd__a211o_1
Xwire2210 net2211 VGND VGND VPWR VPWR net2210 sky130_fd_sc_hd__buf_1
Xwire2221 _07810_ VGND VGND VPWR VPWR net2221 sky130_fd_sc_hd__clkbuf_1
Xwire2232 _07394_ VGND VGND VPWR VPWR net2232 sky130_fd_sc_hd__clkbuf_1
Xwire2243 net2244 VGND VGND VPWR VPWR net2243 sky130_fd_sc_hd__clkbuf_1
Xwire2254 net2255 VGND VGND VPWR VPWR net2254 sky130_fd_sc_hd__clkbuf_1
Xwire1520 _08043_ VGND VGND VPWR VPWR net1520 sky130_fd_sc_hd__buf_1
Xwire2265 net2266 VGND VGND VPWR VPWR net2265 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2276 net2277 VGND VGND VPWR VPWR net2276 sky130_fd_sc_hd__clkbuf_1
Xwire1531 net1532 VGND VGND VPWR VPWR net1531 sky130_fd_sc_hd__clkbuf_1
X_16750_ net7562 net9242 net3380 VGND VGND VPWR VPWR _08764_ sky130_fd_sc_hd__mux2_1
X_13962_ _06225_ _06226_ VGND VGND VPWR VPWR _06227_ sky130_fd_sc_hd__nand2_1
Xwire1542 _07359_ VGND VGND VPWR VPWR net1542 sky130_fd_sc_hd__buf_1
Xwire2298 net2299 VGND VGND VPWR VPWR net2298 sky130_fd_sc_hd__buf_1
Xwire1553 _06509_ VGND VGND VPWR VPWR net1553 sky130_fd_sc_hd__buf_1
Xwire1564 net1565 VGND VGND VPWR VPWR net1564 sky130_fd_sc_hd__clkbuf_1
X_15701_ _07768_ net1530 VGND VGND VPWR VPWR _07772_ sky130_fd_sc_hd__xnor2_1
Xwire1575 net1576 VGND VGND VPWR VPWR net1575 sky130_fd_sc_hd__clkbuf_1
X_12913_ _05184_ _05185_ VGND VGND VPWR VPWR _05186_ sky130_fd_sc_hd__and2_1
Xwire1586 net1587 VGND VGND VPWR VPWR net1586 sky130_fd_sc_hd__buf_1
X_16681_ matmul0.matmul_stage_inst.mult2\[9\] matmul0.matmul_stage_inst.mult1\[9\]
+ VGND VGND VPWR VPWR _08713_ sky130_fd_sc_hd__xor2_1
X_25879_ clknet_leaf_14_clk _00752_ net8621 VGND VGND VPWR VPWR pid_q.ki\[7\] sky130_fd_sc_hd__dfrtp_1
X_13893_ _06137_ _06140_ VGND VGND VPWR VPWR _06159_ sky130_fd_sc_hd__nand2_1
Xwire1597 _05132_ VGND VGND VPWR VPWR net1597 sky130_fd_sc_hd__buf_1
X_18420_ _10172_ _10208_ _10209_ VGND VGND VPWR VPWR _10270_ sky130_fd_sc_hd__o21ai_1
X_15632_ net1857 _07608_ VGND VGND VPWR VPWR _07704_ sky130_fd_sc_hd__or2_1
X_12844_ _05114_ _05115_ _05107_ VGND VGND VPWR VPWR _05117_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_152_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18351_ _10192_ _10195_ _10201_ VGND VGND VPWR VPWR _10202_ sky130_fd_sc_hd__o21a_1
XFILLER_0_174_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15563_ _07569_ _07635_ VGND VGND VPWR VPWR _07636_ sky130_fd_sc_hd__and2_1
X_12775_ net7881 net1356 _04908_ _04914_ VGND VGND VPWR VPWR _05048_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17302_ _09205_ net7630 _09214_ net7607 net4031 VGND VGND VPWR VPWR _09216_ sky130_fd_sc_hd__o311a_1
X_14514_ net5262 _06693_ _06694_ VGND VGND VPWR VPWR _06695_ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18282_ _10057_ _10071_ VGND VGND VPWR VPWR _10133_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15494_ _07543_ _07544_ VGND VGND VPWR VPWR _07567_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17233_ _09163_ _09171_ _09174_ _09175_ _09180_ VGND VGND VPWR VPWR _09181_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_153_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14445_ net5202 _06608_ net3647 net4402 _06637_ VGND VGND VPWR VPWR _06638_ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17164_ _09102_ net527 net6901 VGND VGND VPWR VPWR _09117_ sky130_fd_sc_hd__a21o_1
Xwire850 _05183_ VGND VGND VPWR VPWR net850 sky130_fd_sc_hd__clkbuf_2
X_14376_ net8290 net3637 VGND VGND VPWR VPWR _06585_ sky130_fd_sc_hd__and2_1
XFILLER_0_141_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire861 _01230_ VGND VGND VPWR VPWR net861 sky130_fd_sc_hd__buf_1
Xwire872 _11022_ VGND VGND VPWR VPWR net872 sky130_fd_sc_hd__buf_1
Xwire883 _08060_ VGND VGND VPWR VPWR net883 sky130_fd_sc_hd__clkbuf_1
X_16115_ _08177_ _08180_ VGND VGND VPWR VPWR _08181_ sky130_fd_sc_hd__xnor2_1
X_13327_ net7713 net7687 net1606 net1339 net1946 VGND VGND VPWR VPWR _05600_ sky130_fd_sc_hd__a41o_1
XFILLER_0_51_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire894 _06651_ VGND VGND VPWR VPWR net894 sky130_fd_sc_hd__buf_1
X_17095_ _08820_ _08821_ _09031_ VGND VGND VPWR VPWR _09052_ sky130_fd_sc_hd__mux2_1
X_16046_ net1518 _08047_ _08112_ VGND VGND VPWR VPWR _08113_ sky130_fd_sc_hd__o21a_1
XFILLER_0_177_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13258_ _05529_ _05530_ _05052_ VGND VGND VPWR VPWR _05531_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_122_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13189_ _05456_ _05461_ VGND VGND VPWR VPWR _05462_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19805_ net6215 net6157 VGND VGND VPWR VPWR _11639_ sky130_fd_sc_hd__or2_1
X_17997_ net6940 _09845_ net2555 _09026_ VGND VGND VPWR VPWR _09848_ sky130_fd_sc_hd__a211o_1
XFILLER_0_159_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16948_ net7125 net1818 _08908_ VGND VGND VPWR VPWR _08912_ sky130_fd_sc_hd__or3_1
X_19736_ net6045 net3138 VGND VGND VPWR VPWR _11571_ sky130_fd_sc_hd__nand2_1
X_16879_ _08820_ _08842_ net6525 VGND VGND VPWR VPWR _08843_ sky130_fd_sc_hd__mux2_1
X_19667_ net3881 net6102 VGND VGND VPWR VPWR _11503_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18618_ net6919 _10223_ net3959 VGND VGND VPWR VPWR _10465_ sky130_fd_sc_hd__mux2_1
X_19598_ _10995_ net2106 _11389_ VGND VGND VPWR VPWR _11435_ sky130_fd_sc_hd__or3_1
XFILLER_0_176_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18549_ _10332_ _10339_ _10333_ VGND VGND VPWR VPWR _10398_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_47_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21560_ net5769 net5505 VGND VGND VPWR VPWR _01572_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20511_ net7113 net7088 net7056 net7042 net6514 net6489 VGND VGND VPWR VPWR _12298_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_173_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21491_ net1728 _01390_ _01386_ VGND VGND VPWR VPWR _01504_ sky130_fd_sc_hd__o21a_1
XFILLER_0_172_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23230_ _03098_ _03099_ VGND VGND VPWR VPWR _03100_ sky130_fd_sc_hd__xnor2_2
Xwire6509 net6510 VGND VGND VPWR VPWR net6509 sky130_fd_sc_hd__buf_1
X_20442_ _12228_ VGND VGND VPWR VPWR _12236_ sky130_fd_sc_hd__inv_2
Xmax_length2218 net2219 VGND VGND VPWR VPWR net2218 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire5808 net5802 VGND VGND VPWR VPWR net5808 sky130_fd_sc_hd__clkbuf_1
X_23161_ _03028_ _03029_ _03030_ VGND VGND VPWR VPWR _03031_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20373_ _09006_ _12171_ VGND VGND VPWR VPWR _12172_ sky130_fd_sc_hd__nor2_1
Xmax_length1528 _07902_ VGND VGND VPWR VPWR net1528 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22112_ net802 _02079_ _02117_ VGND VGND VPWR VPWR _02118_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_28_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23092_ _02948_ _02961_ VGND VGND VPWR VPWR _02962_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22043_ _02038_ _02049_ VGND VGND VPWR VPWR _02050_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25802_ clknet_leaf_30_clk _00675_ net8676 VGND VGND VPWR VPWR pid_q.curr_int\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_177_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23994_ net7504 _03856_ _03857_ VGND VGND VPWR VPWR _03858_ sky130_fd_sc_hd__and3_1
X_25733_ clknet_leaf_10_clk _00606_ net8555 VGND VGND VPWR VPWR pid_d.ki\[7\] sky130_fd_sc_hd__dfrtp_1
X_22945_ _02827_ _02833_ net8904 VGND VGND VPWR VPWR _00646_ sky130_fd_sc_hd__o21a_1
XFILLER_0_183_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25664_ clknet_leaf_121_clk _00537_ net8396 VGND VGND VPWR VPWR pid_d.prev_error\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_22876_ _02770_ _02771_ VGND VGND VPWR VPWR _02772_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24615_ net1651 net1649 _04435_ _04469_ VGND VGND VPWR VPWR _04470_ sky130_fd_sc_hd__a31o_1
X_21827_ _01832_ _01835_ VGND VGND VPWR VPWR _01836_ sky130_fd_sc_hd__xnor2_2
X_25595_ clknet_leaf_106_clk _00468_ net8355 VGND VGND VPWR VPWR cordic0.slte0.opB\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout8328 net8339 VGND VGND VPWR VPWR net8328 sky130_fd_sc_hd__clkbuf_1
Xfanout7605 net7613 VGND VGND VPWR VPWR net7605 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24546_ _04395_ _04401_ VGND VGND VPWR VPWR _04402_ sky130_fd_sc_hd__nand2_1
Xwire8412 net8413 VGND VGND VPWR VPWR net8412 sky130_fd_sc_hd__buf_1
X_21758_ _01666_ _01668_ VGND VGND VPWR VPWR _01768_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8434 net8432 VGND VGND VPWR VPWR net8434 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout7649 svm0.periodTop\[13\] VGND VGND VPWR VPWR net7649 sky130_fd_sc_hd__buf_1
XFILLER_0_135_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20709_ net6051 _12475_ VGND VGND VPWR VPWR _12482_ sky130_fd_sc_hd__nand2_1
Xwire8456 net8453 VGND VGND VPWR VPWR net8456 sky130_fd_sc_hd__buf_1
X_24477_ net5175 pid_q.prev_int\[12\] VGND VGND VPWR VPWR _04334_ sky130_fd_sc_hd__or2_1
Xwire8467 net8465 VGND VGND VPWR VPWR net8467 sky130_fd_sc_hd__buf_1
Xwire7733 net7724 VGND VGND VPWR VPWR net7733 sky130_fd_sc_hd__buf_1
X_21689_ _01577_ _01579_ _01699_ VGND VGND VPWR VPWR _01700_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8478 net8475 VGND VGND VPWR VPWR net8478 sky130_fd_sc_hd__buf_1
Xwire7744 net7741 VGND VGND VPWR VPWR net7744 sky130_fd_sc_hd__buf_1
X_14230_ _06482_ _06487_ net7602 VGND VGND VPWR VPWR _06488_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8489 net8488 VGND VGND VPWR VPWR net8489 sky130_fd_sc_hd__buf_1
X_23428_ _03296_ _03297_ VGND VGND VPWR VPWR _03298_ sky130_fd_sc_hd__nor2_1
Xwire7766 net7767 VGND VGND VPWR VPWR net7766 sky130_fd_sc_hd__buf_1
Xwire157 _06431_ VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__buf_1
XFILLER_0_135_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire168 net169 VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_1
Xwire7788 net7789 VGND VGND VPWR VPWR net7788 sky130_fd_sc_hd__buf_1
XFILLER_0_22_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire179 _12027_ VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__buf_1
XFILLER_0_180_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14161_ net403 _06368_ VGND VGND VPWR VPWR _06422_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23359_ net1674 _03228_ VGND VGND VPWR VPWR _03229_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_34_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length2763 _07190_ VGND VGND VPWR VPWR net2763 sky130_fd_sc_hd__clkbuf_1
X_13112_ net7801 net2976 net2974 VGND VGND VPWR VPWR _05385_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14092_ _06352_ _06354_ VGND VGND VPWR VPWR _06355_ sky130_fd_sc_hd__xor2_1
XFILLER_0_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25029_ _03671_ _04774_ _04781_ VGND VGND VPWR VPWR _04782_ sky130_fd_sc_hd__a21o_1
X_13043_ _05311_ _05312_ _05315_ net790 _05204_ VGND VGND VPWR VPWR _05316_ sky130_fd_sc_hd__a32o_1
X_17920_ _09747_ _09760_ _09769_ _09770_ VGND VGND VPWR VPWR _09771_ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17851_ _09622_ net3265 VGND VGND VPWR VPWR _09702_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2040 net2041 VGND VGND VPWR VPWR net2040 sky130_fd_sc_hd__buf_1
Xwire2051 _02307_ VGND VGND VPWR VPWR net2051 sky130_fd_sc_hd__buf_1
X_16802_ cordic0.cos\[4\] net7180 net3369 VGND VGND VPWR VPWR _08791_ sky130_fd_sc_hd__mux2_1
Xwire2062 net2063 VGND VGND VPWR VPWR net2062 sky130_fd_sc_hd__buf_2
Xwire2073 _01155_ VGND VGND VPWR VPWR net2073 sky130_fd_sc_hd__buf_1
X_17782_ net7119 _09632_ VGND VGND VPWR VPWR _09633_ sky130_fd_sc_hd__nand2_1
X_14994_ net3536 net3529 _07065_ _07067_ VGND VGND VPWR VPWR _07068_ sky130_fd_sc_hd__o31a_1
Xwire2084 net2085 VGND VGND VPWR VPWR net2084 sky130_fd_sc_hd__clkbuf_2
Xwire2095 net2096 VGND VGND VPWR VPWR net2095 sky130_fd_sc_hd__buf_1
Xwire1361 net1362 VGND VGND VPWR VPWR net1361 sky130_fd_sc_hd__clkbuf_2
X_19521_ _11286_ _11355_ _11356_ _11357_ _11288_ VGND VGND VPWR VPWR _11358_ sky130_fd_sc_hd__a32o_1
X_16733_ net7573 matmul0.b\[3\] net3702 VGND VGND VPWR VPWR _08755_ sky130_fd_sc_hd__mux2_1
X_13945_ _06162_ _06210_ VGND VGND VPWR VPWR _06211_ sky130_fd_sc_hd__xnor2_1
Xwire1372 net1373 VGND VGND VPWR VPWR net1372 sky130_fd_sc_hd__buf_1
Xwire1383 _03668_ VGND VGND VPWR VPWR net1383 sky130_fd_sc_hd__buf_1
Xwire1394 _12428_ VGND VGND VPWR VPWR net1394 sky130_fd_sc_hd__buf_1
X_19452_ net6025 VGND VGND VPWR VPWR _11289_ sky130_fd_sc_hd__inv_2
X_16664_ matmul0.matmul_stage_inst.mult1\[6\] VGND VGND VPWR VPWR _08698_ sky130_fd_sc_hd__inv_2
X_13876_ net532 _06080_ VGND VGND VPWR VPWR _06143_ sky130_fd_sc_hd__and2_1
XFILLER_0_158_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15615_ net2851 _07686_ VGND VGND VPWR VPWR _07687_ sky130_fd_sc_hd__nand2_1
X_18403_ net1073 _10157_ _10253_ VGND VGND VPWR VPWR _10254_ sky130_fd_sc_hd__a21oi_2
X_12827_ _05040_ _05041_ _05099_ VGND VGND VPWR VPWR _05100_ sky130_fd_sc_hd__o21ai_2
X_19383_ _11207_ _11219_ VGND VGND VPWR VPWR _11220_ sky130_fd_sc_hd__xnor2_1
X_16595_ net6658 VGND VGND VPWR VPWR _08646_ sky130_fd_sc_hd__inv_2
XFILLER_0_174_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18334_ net1211 net1073 VGND VGND VPWR VPWR _10185_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15546_ net3423 net2689 _07618_ VGND VGND VPWR VPWR _07619_ sky130_fd_sc_hd__o21a_1
X_12758_ _05020_ _05025_ _05030_ VGND VGND VPWR VPWR _05031_ sky130_fd_sc_hd__a21o_1
XFILLER_0_189_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8862 net8874 VGND VGND VPWR VPWR net8862 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout8873 net146 VGND VGND VPWR VPWR net8873 sky130_fd_sc_hd__clkbuf_1
X_18265_ _10113_ _10114_ _10093_ VGND VGND VPWR VPWR _10116_ sky130_fd_sc_hd__a21o_1
XFILLER_0_154_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15477_ _07402_ net1274 net1875 _07546_ VGND VGND VPWR VPWR _07551_ sky130_fd_sc_hd__a211o_1
XFILLER_0_84_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12689_ net7303 _04856_ net4278 VGND VGND VPWR VPWR _04962_ sky130_fd_sc_hd__nand3_1
Xfanout8895 net8899 VGND VGND VPWR VPWR net8895 sky130_fd_sc_hd__buf_1
X_17216_ net5998 _08834_ net2583 VGND VGND VPWR VPWR _09165_ sky130_fd_sc_hd__mux2_2
XFILLER_0_86_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14428_ net8123 net3631 VGND VGND VPWR VPWR _06625_ sky130_fd_sc_hd__and2_1
X_18196_ _08984_ net3952 _09609_ VGND VGND VPWR VPWR _10047_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17147_ net1504 net822 VGND VGND VPWR VPWR _09101_ sky130_fd_sc_hd__or2_1
XFILLER_0_188_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire680 _05836_ VGND VGND VPWR VPWR net680 sky130_fd_sc_hd__clkbuf_1
X_14359_ net994 VGND VGND VPWR VPWR _06572_ sky130_fd_sc_hd__buf_1
Xwire691 _04591_ VGND VGND VPWR VPWR net691 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17078_ net2609 _09030_ _09035_ net5990 VGND VGND VPWR VPWR _09036_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16029_ net2722 net3417 VGND VGND VPWR VPWR _08096_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_179_Left_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length8409 net8405 VGND VGND VPWR VPWR net8409 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_46_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19719_ net569 _11544_ _11553_ net3857 VGND VGND VPWR VPWR _11554_ sky130_fd_sc_hd__a22o_1
X_20991_ _00952_ _00955_ net3111 VGND VGND VPWR VPWR _01007_ sky130_fd_sc_hd__nand3_2
X_22730_ pid_d.ki\[1\] _02664_ net1688 VGND VGND VPWR VPWR _02665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22661_ _02395_ net3079 net856 _02615_ net8905 VGND VGND VPWR VPWR _00580_ sky130_fd_sc_hd__o311a_1
XFILLER_0_153_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24400_ net9077 net3757 net2433 _04258_ VGND VGND VPWR VPWR _00676_ sky130_fd_sc_hd__a22o_1
X_21612_ net1179 _01621_ _01623_ VGND VGND VPWR VPWR _01624_ sky130_fd_sc_hd__a21oi_1
X_25380_ clknet_leaf_64_clk _00263_ net8663 VGND VGND VPWR VPWR matmul0.alpha_pass\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_22592_ net7287 _02566_ VGND VGND VPWR VPWR _02569_ sky130_fd_sc_hd__nor2_1
XFILLER_0_168_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24331_ net5177 pid_q.prev_int\[11\] VGND VGND VPWR VPWR _04190_ sky130_fd_sc_hd__xnor2_1
Xwire7007 net7004 VGND VGND VPWR VPWR net7007 sky130_fd_sc_hd__buf_1
XFILLER_0_75_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21543_ _01448_ _01450_ _01449_ VGND VGND VPWR VPWR _01555_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_188_Left_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24262_ net1159 _04086_ _04074_ VGND VGND VPWR VPWR _04122_ sky130_fd_sc_hd__o21a_1
X_21474_ _01483_ _01486_ VGND VGND VPWR VPWR _01487_ sky130_fd_sc_hd__xnor2_2
Xwire6317 net6319 VGND VGND VPWR VPWR net6317 sky130_fd_sc_hd__buf_1
Xwire6328 net6329 VGND VGND VPWR VPWR net6328 sky130_fd_sc_hd__buf_1
Xwire6339 net6340 VGND VGND VPWR VPWR net6339 sky130_fd_sc_hd__buf_1
XFILLER_0_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23213_ _03075_ _03078_ VGND VGND VPWR VPWR _03083_ sky130_fd_sc_hd__and2_1
Xwire5605 net5607 VGND VGND VPWR VPWR net5605 sky130_fd_sc_hd__buf_1
X_20425_ net863 _12220_ VGND VGND VPWR VPWR _12221_ sky130_fd_sc_hd__xnor2_1
Xmax_length1303 _06522_ VGND VGND VPWR VPWR net1303 sky130_fd_sc_hd__clkbuf_1
Xwire5616 net5614 VGND VGND VPWR VPWR net5616 sky130_fd_sc_hd__buf_1
X_24193_ net4590 net4836 VGND VGND VPWR VPWR _04054_ sky130_fd_sc_hd__nand2_1
Xwire5627 net5625 VGND VGND VPWR VPWR net5627 sky130_fd_sc_hd__buf_1
Xwire5638 net5636 VGND VGND VPWR VPWR net5638 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_15_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4904 net4905 VGND VGND VPWR VPWR net4904 sky130_fd_sc_hd__clkbuf_1
Xwire5649 net5645 VGND VGND VPWR VPWR net5649 sky130_fd_sc_hd__buf_1
XFILLER_0_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23144_ _03010_ _03013_ VGND VGND VPWR VPWR _03014_ sky130_fd_sc_hd__xnor2_2
X_20356_ net6472 net4037 _12084_ VGND VGND VPWR VPWR _12157_ sky130_fd_sc_hd__a21o_1
Xwire4926 net4927 VGND VGND VPWR VPWR net4926 sky130_fd_sc_hd__buf_1
Xmax_length1369 net1370 VGND VGND VPWR VPWR net1369 sky130_fd_sc_hd__buf_1
Xwire4937 net4938 VGND VGND VPWR VPWR net4937 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_141_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4948 net4949 VGND VGND VPWR VPWR net4948 sky130_fd_sc_hd__buf_1
XFILLER_0_31_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23075_ _02939_ _02944_ VGND VGND VPWR VPWR _02945_ sky130_fd_sc_hd__xnor2_1
X_20287_ net6516 net6468 VGND VGND VPWR VPWR _12093_ sky130_fd_sc_hd__or2_1
X_22026_ _02031_ _02032_ VGND VGND VPWR VPWR _02033_ sky130_fd_sc_hd__xor2_1
Xhold10 _00408_ VGND VGND VPWR VPWR net8963 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 matmul0.matmul_stage_inst.c\[5\] VGND VGND VPWR VPWR net8974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 pid_q.target\[3\] VGND VGND VPWR VPWR net8985 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 pid_q.curr_int\[2\] VGND VGND VPWR VPWR net8996 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 matmul0.matmul_stage_inst.d\[0\] VGND VGND VPWR VPWR net9007 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 pid_d.curr_int\[9\] VGND VGND VPWR VPWR net9018 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 cordic0.cos\[1\] VGND VGND VPWR VPWR net9029 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 matmul0.matmul_stage_inst.c\[11\] VGND VGND VPWR VPWR net9040 sky130_fd_sc_hd__dlygate4sd3_1
X_23977_ _03737_ _03743_ _03840_ VGND VGND VPWR VPWR _03841_ sky130_fd_sc_hd__a21o_1
Xhold98 svm0.vC\[3\] VGND VGND VPWR VPWR net9051 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13730_ _05927_ _05929_ _05919_ VGND VGND VPWR VPWR _05999_ sky130_fd_sc_hd__o21ba_1
X_25716_ clknet_leaf_9_clk _00589_ net8559 VGND VGND VPWR VPWR pid_d.mult0.a\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_22928_ net8907 _02818_ VGND VGND VPWR VPWR _02819_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13661_ _05927_ _05929_ VGND VGND VPWR VPWR _05931_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25647_ clknet_leaf_122_clk _00520_ net8403 VGND VGND VPWR VPWR pid_d.curr_int\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_196_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22859_ net5364 _02756_ net3066 VGND VGND VPWR VPWR _02757_ sky130_fd_sc_hd__mux2_1
X_15400_ _07405_ _07406_ _07473_ net1280 VGND VGND VPWR VPWR _07474_ sky130_fd_sc_hd__a22oi_1
X_12612_ net3696 VGND VGND VPWR VPWR _00003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16380_ net2707 net2648 VGND VGND VPWR VPWR _08442_ sky130_fd_sc_hd__nor2_1
X_13592_ net367 _05774_ _05852_ _05861_ _05851_ VGND VGND VPWR VPWR _05862_ sky130_fd_sc_hd__o311a_1
X_25578_ clknet_leaf_98_clk _00451_ net8383 VGND VGND VPWR VPWR cordic0.sin\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire8220 net8221 VGND VGND VPWR VPWR net8220 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15331_ _07403_ _07404_ VGND VGND VPWR VPWR _07405_ sky130_fd_sc_hd__and2_1
Xwire8231 net8232 VGND VGND VPWR VPWR net8231 sky130_fd_sc_hd__clkbuf_1
X_24529_ net328 _04385_ VGND VGND VPWR VPWR _04386_ sky130_fd_sc_hd__and2_1
Xwire8242 net28 VGND VGND VPWR VPWR net8242 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8253 net8254 VGND VGND VPWR VPWR net8253 sky130_fd_sc_hd__clkbuf_1
Xwire8264 net8265 VGND VGND VPWR VPWR net8264 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18050_ _09893_ _09900_ VGND VGND VPWR VPWR _09901_ sky130_fd_sc_hd__xnor2_4
Xwire8275 net8276 VGND VGND VPWR VPWR net8275 sky130_fd_sc_hd__clkbuf_1
Xfanout7479 net7487 VGND VGND VPWR VPWR net7479 sky130_fd_sc_hd__buf_1
XFILLER_0_136_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8286 net8287 VGND VGND VPWR VPWR net8286 sky130_fd_sc_hd__clkbuf_1
X_15262_ _07267_ _07299_ net829 _07335_ VGND VGND VPWR VPWR _07336_ sky130_fd_sc_hd__a2bb2o_1
Xwire7541 net7542 VGND VGND VPWR VPWR net7541 sky130_fd_sc_hd__clkbuf_1
Xwire7552 matmul0.op_in\[0\] VGND VGND VPWR VPWR net7552 sky130_fd_sc_hd__clkbuf_1
Xwire8297 net8298 VGND VGND VPWR VPWR net8297 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17001_ _08959_ _08962_ VGND VGND VPWR VPWR _08963_ sky130_fd_sc_hd__xnor2_1
X_14213_ net1121 net1304 net7629 VGND VGND VPWR VPWR _06472_ sky130_fd_sc_hd__o21a_1
Xmax_length3261 net3262 VGND VGND VPWR VPWR net3261 sky130_fd_sc_hd__buf_1
Xwire7574 matmul0.b_in\[1\] VGND VGND VPWR VPWR net7574 sky130_fd_sc_hd__clkbuf_1
Xwire6840 net6841 VGND VGND VPWR VPWR net6840 sky130_fd_sc_hd__buf_1
Xwire7585 net7586 VGND VGND VPWR VPWR net7585 sky130_fd_sc_hd__clkbuf_1
X_15193_ _07255_ _07266_ VGND VGND VPWR VPWR _07267_ sky130_fd_sc_hd__xnor2_1
Xwire6851 net6852 VGND VGND VPWR VPWR net6851 sky130_fd_sc_hd__buf_1
Xwire7596 net7597 VGND VGND VPWR VPWR net7596 sky130_fd_sc_hd__clkbuf_1
Xwire6862 net6863 VGND VGND VPWR VPWR net6862 sky130_fd_sc_hd__buf_1
XFILLER_0_104_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6873 net6874 VGND VGND VPWR VPWR net6873 sky130_fd_sc_hd__buf_1
X_14144_ net1314 VGND VGND VPWR VPWR _06405_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2593 net2594 VGND VGND VPWR VPWR net2593 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_158_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14075_ net1125 _06222_ net7604 VGND VGND VPWR VPWR _06338_ sky130_fd_sc_hd__a21o_1
X_18952_ net3917 _10788_ VGND VGND VPWR VPWR _10789_ sky130_fd_sc_hd__nor2_1
X_13026_ _05292_ _05295_ _05298_ VGND VGND VPWR VPWR _05299_ sky130_fd_sc_hd__a21oi_1
X_17903_ net7133 net2557 VGND VGND VPWR VPWR _09754_ sky130_fd_sc_hd__xnor2_4
X_18883_ net6781 _10682_ _10724_ _10666_ VGND VGND VPWR VPWR _10725_ sky130_fd_sc_hd__a2bb2o_1
X_17834_ net6974 net6995 VGND VGND VPWR VPWR _09685_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14977_ net3544 net3541 VGND VGND VPWR VPWR _07051_ sky130_fd_sc_hd__nor2_1
X_17765_ net7135 _09613_ net3265 net3346 VGND VGND VPWR VPWR _09616_ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1180 _01482_ VGND VGND VPWR VPWR net1180 sky130_fd_sc_hd__buf_1
X_19504_ _11327_ net1419 VGND VGND VPWR VPWR _11341_ sky130_fd_sc_hd__xnor2_1
Xwire1191 _11475_ VGND VGND VPWR VPWR net1191 sky130_fd_sc_hd__dlymetal6s2s_1
X_13928_ net7704 net2953 net3672 VGND VGND VPWR VPWR _06194_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16716_ matmul0.matmul_stage_inst.mult2\[14\] matmul0.matmul_stage_inst.mult1\[14\]
+ VGND VGND VPWR VPWR _08743_ sky130_fd_sc_hd__xor2_1
X_17696_ net3389 net1796 net6655 VGND VGND VPWR VPWR _09573_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_92_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19435_ net6145 net6163 VGND VGND VPWR VPWR _11272_ sky130_fd_sc_hd__or2_1
X_16647_ _08682_ _08683_ VGND VGND VPWR VPWR _08684_ sky130_fd_sc_hd__xnor2_1
X_13859_ net841 _06048_ VGND VGND VPWR VPWR _06126_ sky130_fd_sc_hd__nand2_1
XFILLER_0_186_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19366_ _11185_ _11200_ _11201_ _11202_ VGND VGND VPWR VPWR _11203_ sky130_fd_sc_hd__a2bb2o_1
X_16578_ net3471 VGND VGND VPWR VPWR _08636_ sky130_fd_sc_hd__buf_1
XFILLER_0_8_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18317_ _10166_ _10167_ VGND VGND VPWR VPWR _10168_ sky130_fd_sc_hd__xnor2_1
X_15529_ net6542 matmul0.matmul_stage_inst.c\[14\] matmul0.matmul_stage_inst.b\[14\]
+ net6614 VGND VGND VPWR VPWR _07602_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19297_ net3167 _11133_ VGND VGND VPWR VPWR _11134_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8692 net8698 VGND VGND VPWR VPWR net8692 sky130_fd_sc_hd__buf_1
XFILLER_0_115_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18248_ net4044 _09648_ net3267 net6964 VGND VGND VPWR VPWR _10099_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_154_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18179_ net3340 net7142 VGND VGND VPWR VPWR _10030_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20210_ net1770 _12032_ _12033_ VGND VGND VPWR VPWR _00466_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21190_ _01163_ _01204_ _01205_ VGND VGND VPWR VPWR _01206_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20141_ _11889_ _11891_ VGND VGND VPWR VPWR _11968_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2809 _07100_ VGND VGND VPWR VPWR net2809 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20072_ net1404 _11899_ VGND VGND VPWR VPWR _11901_ sky130_fd_sc_hd__nor2_1
X_23900_ pid_q.prev_error\[5\] pid_q.curr_error\[5\] VGND VGND VPWR VPWR _03765_ sky130_fd_sc_hd__xnor2_1
X_24880_ pid_q.ki\[8\] net2397 net3009 pid_q.kp\[8\] VGND VGND VPWR VPWR _04678_ sky130_fd_sc_hd__a22o_1
X_23831_ net5036 net4499 VGND VGND VPWR VPWR _03696_ sky130_fd_sc_hd__nand2_1
XFILLER_0_164_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23762_ _03622_ _03627_ VGND VGND VPWR VPWR _03628_ sky130_fd_sc_hd__xnor2_1
X_20974_ _00987_ _00988_ VGND VGND VPWR VPWR _00990_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25501_ clknet_leaf_41_clk _00381_ net8768 VGND VGND VPWR VPWR svm0.delta\[6\] sky130_fd_sc_hd__dfrtp_1
X_22713_ _02650_ VGND VGND VPWR VPWR _00597_ sky130_fd_sc_hd__clkbuf_1
Xmax_length6826 net6827 VGND VGND VPWR VPWR net6826 sky130_fd_sc_hd__buf_1
XFILLER_0_94_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23693_ _03451_ _03461_ _03449_ VGND VGND VPWR VPWR _03560_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25432_ clknet_leaf_96_clk _00315_ net8399 VGND VGND VPWR VPWR matmul0.sin\[5\] sky130_fd_sc_hd__dfrtp_1
X_22644_ net3090 _02564_ _02565_ net3080 VGND VGND VPWR VPWR _02607_ sky130_fd_sc_hd__a31o_1
XFILLER_0_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25363_ clknet_leaf_72_clk _00246_ net8478 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult2\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22575_ net3091 _02554_ _02555_ VGND VGND VPWR VPWR _02556_ sky130_fd_sc_hd__and3_1
XFILLER_0_180_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24314_ _04171_ _04040_ _04173_ VGND VGND VPWR VPWR _04174_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21526_ net4357 _01537_ _01538_ VGND VGND VPWR VPWR _01539_ sky130_fd_sc_hd__and3_1
Xwire6103 net6100 VGND VGND VPWR VPWR net6103 sky130_fd_sc_hd__buf_1
X_25294_ clknet_leaf_88_clk _00177_ net8431 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.d\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6125 net6126 VGND VGND VPWR VPWR net6125 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6136 net6137 VGND VGND VPWR VPWR net6136 sky130_fd_sc_hd__buf_1
XFILLER_0_32_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5402 net5403 VGND VGND VPWR VPWR net5402 sky130_fd_sc_hd__clkbuf_1
X_24245_ _04048_ net589 VGND VGND VPWR VPWR _04106_ sky130_fd_sc_hd__and2_1
Xwire6147 net6148 VGND VGND VPWR VPWR net6147 sky130_fd_sc_hd__clkbuf_2
X_21457_ _01466_ _01469_ VGND VGND VPWR VPWR _01470_ sky130_fd_sc_hd__xnor2_1
Xwire6158 net6156 VGND VGND VPWR VPWR net6158 sky130_fd_sc_hd__buf_1
Xwire5424 net5425 VGND VGND VPWR VPWR net5424 sky130_fd_sc_hd__clkbuf_1
Xfanout4639 net4643 VGND VGND VPWR VPWR net4639 sky130_fd_sc_hd__buf_1
Xwire5435 net5430 VGND VGND VPWR VPWR net5435 sky130_fd_sc_hd__buf_1
Xwire5446 net5447 VGND VGND VPWR VPWR net5446 sky130_fd_sc_hd__clkbuf_1
X_20408_ _12145_ net2089 VGND VGND VPWR VPWR _12205_ sky130_fd_sc_hd__xnor2_2
Xwire4712 net4713 VGND VGND VPWR VPWR net4712 sky130_fd_sc_hd__clkbuf_1
X_24176_ pid_q.prev_int\[8\] VGND VGND VPWR VPWR _04037_ sky130_fd_sc_hd__inv_2
Xwire5457 net5458 VGND VGND VPWR VPWR net5457 sky130_fd_sc_hd__buf_1
X_21388_ _01265_ _01266_ _01401_ VGND VGND VPWR VPWR _01402_ sky130_fd_sc_hd__a21oi_2
Xwire4723 net4721 VGND VGND VPWR VPWR net4723 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire5468 net5469 VGND VGND VPWR VPWR net5468 sky130_fd_sc_hd__clkbuf_1
Xwire5479 net5480 VGND VGND VPWR VPWR net5479 sky130_fd_sc_hd__buf_1
Xwire4745 net4746 VGND VGND VPWR VPWR net4745 sky130_fd_sc_hd__clkbuf_1
X_23127_ net5085 net4683 VGND VGND VPWR VPWR _02997_ sky130_fd_sc_hd__nand2_1
Xwire4756 net4757 VGND VGND VPWR VPWR net4756 sky130_fd_sc_hd__clkbuf_1
X_20339_ net1817 VGND VGND VPWR VPWR _12142_ sky130_fd_sc_hd__buf_1
Xwire4767 net4761 VGND VGND VPWR VPWR net4767 sky130_fd_sc_hd__buf_1
Xmax_length1199 net1200 VGND VGND VPWR VPWR net1199 sky130_fd_sc_hd__clkbuf_1
Xwire4778 net4773 VGND VGND VPWR VPWR net4778 sky130_fd_sc_hd__buf_1
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4789 net4791 VGND VGND VPWR VPWR net4789 sky130_fd_sc_hd__dlymetal6s2s_1
X_23058_ net4887 net4760 VGND VGND VPWR VPWR _02928_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput100 pid_d_data[12] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
Xinput111 pid_d_data[8] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_1
Xinput122 pid_q_addr[2] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_1
X_14900_ net6620 net6644 matmul0.matmul_stage_inst.f\[1\] VGND VGND VPWR VPWR _06974_
+ sky130_fd_sc_hd__o21a_1
X_22009_ pid_d.prev_int\[8\] VGND VGND VPWR VPWR _02016_ sky130_fd_sc_hd__inv_2
Xinput133 pid_q_data[12] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_1
X_15880_ _07940_ _07948_ VGND VGND VPWR VPWR _07949_ sky130_fd_sc_hd__xnor2_1
Xinput144 pid_q_data[8] VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_1
X_14831_ _06932_ VGND VGND VPWR VPWR _00187_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17550_ _09430_ _09431_ VGND VGND VPWR VPWR _09432_ sky130_fd_sc_hd__nor2_1
X_14762_ net9128 net2858 net2865 _06891_ VGND VGND VPWR VPWR _00159_ sky130_fd_sc_hd__a22o_1
X_16501_ net2750 net2744 VGND VGND VPWR VPWR _08561_ sky130_fd_sc_hd__nand2_1
X_13713_ _05906_ _05980_ _05981_ VGND VGND VPWR VPWR _05982_ sky130_fd_sc_hd__o21ai_1
X_17481_ _09295_ _09367_ _09371_ VGND VGND VPWR VPWR _09372_ sky130_fd_sc_hd__a21o_1
X_14693_ net7454 _06839_ VGND VGND VPWR VPWR _06840_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19220_ net3178 _11056_ net3890 VGND VGND VPWR VPWR _11057_ sky130_fd_sc_hd__a21o_1
X_16432_ _08480_ _08491_ _08492_ VGND VGND VPWR VPWR _08493_ sky130_fd_sc_hd__o21a_1
X_13644_ _05906_ _05913_ VGND VGND VPWR VPWR _05914_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_160_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19151_ _10984_ _10987_ VGND VGND VPWR VPWR _10988_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_184_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16363_ _08311_ net1083 _08425_ VGND VGND VPWR VPWR _08426_ sky130_fd_sc_hd__o21ai_1
X_13575_ net679 _05845_ VGND VGND VPWR VPWR _05846_ sky130_fd_sc_hd__xor2_1
XFILLER_0_87_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18102_ _09872_ _09873_ VGND VGND VPWR VPWR _09953_ sky130_fd_sc_hd__and2_1
Xwire8050 net8051 VGND VGND VPWR VPWR net8050 sky130_fd_sc_hd__buf_1
Xwire8061 net8058 VGND VGND VPWR VPWR net8061 sky130_fd_sc_hd__buf_1
X_15314_ net3545 net3558 VGND VGND VPWR VPWR _07388_ sky130_fd_sc_hd__nor2_1
X_19082_ _10917_ _10918_ VGND VGND VPWR VPWR _10919_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8072 net8073 VGND VGND VPWR VPWR net8072 sky130_fd_sc_hd__clkbuf_1
X_16294_ _08356_ _08357_ VGND VGND VPWR VPWR _08358_ sky130_fd_sc_hd__and2b_1
Xfanout6531 net6538 VGND VGND VPWR VPWR net6531 sky130_fd_sc_hd__buf_1
Xwire8083 net152 VGND VGND VPWR VPWR net8083 sky130_fd_sc_hd__clkbuf_1
Xwire8094 net8095 VGND VGND VPWR VPWR net8094 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout6553 net6564 VGND VGND VPWR VPWR net6553 sky130_fd_sc_hd__clkbuf_1
X_18033_ _09856_ _09883_ VGND VGND VPWR VPWR _09884_ sky130_fd_sc_hd__nor2_1
Xwire7360 matmul0.alpha_pass\[1\] VGND VGND VPWR VPWR net7360 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15245_ net3576 net3572 net4221 net4219 VGND VGND VPWR VPWR _07319_ sky130_fd_sc_hd__o22a_1
Xwire7371 net7372 VGND VGND VPWR VPWR net7371 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5830 net5847 VGND VGND VPWR VPWR net5830 sky130_fd_sc_hd__buf_1
Xfanout6586 net6591 VGND VGND VPWR VPWR net6586 sky130_fd_sc_hd__buf_1
Xwire7393 net7394 VGND VGND VPWR VPWR net7393 sky130_fd_sc_hd__clkbuf_1
Xfanout6597 net6608 VGND VGND VPWR VPWR net6597 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_112_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3091 _02553_ VGND VGND VPWR VPWR net3091 sky130_fd_sc_hd__buf_1
Xwire6670 net6663 VGND VGND VPWR VPWR net6670 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6681 svm0.state\[0\] VGND VGND VPWR VPWR net6681 sky130_fd_sc_hd__clkbuf_1
X_15176_ _07229_ net2242 VGND VGND VPWR VPWR _07250_ sky130_fd_sc_hd__xor2_2
Xwire6692 net6690 VGND VGND VPWR VPWR net6692 sky130_fd_sc_hd__buf_1
XFILLER_0_105_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14127_ net7625 _06387_ _06388_ VGND VGND VPWR VPWR _06389_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5980 pid_d.curr_int\[5\] VGND VGND VPWR VPWR net5980 sky130_fd_sc_hd__buf_1
X_19984_ net3862 net2095 VGND VGND VPWR VPWR _11815_ sky130_fd_sc_hd__nor2_1
XFILLER_0_185_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14058_ net9161 net1127 net219 net1927 VGND VGND VPWR VPWR _00025_ sky130_fd_sc_hd__a22o_1
X_18935_ net6816 net6779 _10773_ net6830 net6794 VGND VGND VPWR VPWR _10774_ sky130_fd_sc_hd__o221a_1
XFILLER_0_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13009_ net1336 _05100_ _05093_ VGND VGND VPWR VPWR _05282_ sky130_fd_sc_hd__a21o_1
XFILLER_0_193_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18866_ _10706_ _10707_ net6834 VGND VGND VPWR VPWR _10708_ sky130_fd_sc_hd__mux2_1
X_17817_ net3259 net2563 VGND VGND VPWR VPWR _09668_ sky130_fd_sc_hd__and2_1
X_18797_ net6867 net6878 VGND VGND VPWR VPWR _10641_ sky130_fd_sc_hd__nand2_1
XFILLER_0_179_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17748_ net7019 net6995 VGND VGND VPWR VPWR _09599_ sky130_fd_sc_hd__and2b_1
XFILLER_0_178_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17679_ svm0.tA\[7\] _09539_ VGND VGND VPWR VPWR _09559_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19418_ net6265 net3886 VGND VGND VPWR VPWR _11255_ sky130_fd_sc_hd__nand2_1
X_20690_ _08993_ _12464_ VGND VGND VPWR VPWR _12465_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19349_ net2108 _11151_ VGND VGND VPWR VPWR _11186_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22360_ net2471 _02362_ VGND VGND VPWR VPWR _02363_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21311_ _00877_ _00933_ _00931_ VGND VGND VPWR VPWR _01326_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_170_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22291_ _02291_ _02294_ VGND VGND VPWR VPWR _02295_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24030_ net4591 net4881 VGND VGND VPWR VPWR _03893_ sky130_fd_sc_hd__nand2_2
XFILLER_0_14_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21242_ net5861 net5475 VGND VGND VPWR VPWR _01257_ sky130_fd_sc_hd__nand2_2
Xwire4008 _09358_ VGND VGND VPWR VPWR net4008 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4019 _09243_ VGND VGND VPWR VPWR net4019 sky130_fd_sc_hd__buf_1
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21173_ _01181_ _01183_ net3807 VGND VGND VPWR VPWR _01189_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3307 net3309 VGND VGND VPWR VPWR net3307 sky130_fd_sc_hd__buf_1
XFILLER_0_111_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3318 net3319 VGND VGND VPWR VPWR net3318 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3329 net3330 VGND VGND VPWR VPWR net3329 sky130_fd_sc_hd__clkbuf_1
X_20124_ net2582 _11901_ VGND VGND VPWR VPWR _11952_ sky130_fd_sc_hd__or2_1
Xwire2606 _08933_ VGND VGND VPWR VPWR net2606 sky130_fd_sc_hd__buf_1
Xwire2617 _08636_ VGND VGND VPWR VPWR net2617 sky130_fd_sc_hd__buf_1
Xwire2628 net2629 VGND VGND VPWR VPWR net2628 sky130_fd_sc_hd__clkbuf_2
Xwire2639 _07843_ VGND VGND VPWR VPWR net2639 sky130_fd_sc_hd__buf_1
X_24932_ _04715_ VGND VGND VPWR VPWR _00751_ sky130_fd_sc_hd__clkbuf_1
X_20055_ net6077 _11490_ VGND VGND VPWR VPWR _11884_ sky130_fd_sc_hd__and2_1
Xwire1905 _06991_ VGND VGND VPWR VPWR net1905 sky130_fd_sc_hd__clkbuf_1
Xwire1916 net1917 VGND VGND VPWR VPWR net1916 sky130_fd_sc_hd__buf_1
Xwire1927 _05857_ VGND VGND VPWR VPWR net1927 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1938 net1939 VGND VGND VPWR VPWR net1938 sky130_fd_sc_hd__buf_1
Xwire1949 _05191_ VGND VGND VPWR VPWR net1949 sky130_fd_sc_hd__buf_1
X_24863_ _04666_ VGND VGND VPWR VPWR _00731_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23814_ _03652_ _03654_ _03653_ VGND VGND VPWR VPWR _03679_ sky130_fd_sc_hd__a21o_1
XFILLER_0_139_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length8047 net8048 VGND VGND VPWR VPWR net8047 sky130_fd_sc_hd__clkbuf_1
X_24794_ _04614_ _04613_ net5206 VGND VGND VPWR VPWR _04619_ sky130_fd_sc_hd__o21ai_1
X_23745_ net1662 _03610_ VGND VGND VPWR VPWR _03611_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20957_ _00970_ _00972_ _00883_ VGND VGND VPWR VPWR _00973_ sky130_fd_sc_hd__mux2_1
Xmax_length7379 matmul0.matmul_stage_inst.f\[15\] VGND VGND VPWR VPWR net7379 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23676_ _03423_ _03447_ _03446_ VGND VGND VPWR VPWR _03543_ sky130_fd_sc_hd__a21o_1
Xmax_length6678 net6677 VGND VGND VPWR VPWR net6678 sky130_fd_sc_hd__clkbuf_2
X_20888_ _00901_ _00902_ _00903_ VGND VGND VPWR VPWR _00904_ sky130_fd_sc_hd__o21ai_1
Xmax_length5944 net5945 VGND VGND VPWR VPWR net5944 sky130_fd_sc_hd__buf_1
X_25415_ clknet_leaf_89_clk _00298_ net8424 VGND VGND VPWR VPWR matmul0.cos\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_192_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22627_ net8905 _02596_ VGND VGND VPWR VPWR _02597_ sky130_fd_sc_hd__and2_1
XFILLER_0_165_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13360_ net843 _05632_ VGND VGND VPWR VPWR _05633_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_24_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25346_ clknet_leaf_72_clk _00229_ net8470 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_22558_ _04865_ net3775 VGND VGND VPWR VPWR _02542_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_165_Right_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21509_ net806 net757 VGND VGND VPWR VPWR _01522_ sky130_fd_sc_hd__or2_1
X_13291_ _05486_ _05563_ VGND VGND VPWR VPWR _05564_ sky130_fd_sc_hd__xor2_1
XFILLER_0_51_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25277_ clknet_leaf_71_clk _00160_ net8457 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.c\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22489_ net5390 _02486_ _02489_ net5647 VGND VGND VPWR VPWR _02490_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5210 net5211 VGND VGND VPWR VPWR net5210 sky130_fd_sc_hd__clkbuf_1
Xwire5221 net5222 VGND VGND VPWR VPWR net5221 sky130_fd_sc_hd__clkbuf_1
X_15030_ _07094_ net1895 VGND VGND VPWR VPWR _07104_ sky130_fd_sc_hd__xnor2_1
X_24228_ _03994_ _03998_ _03999_ VGND VGND VPWR VPWR _04089_ sky130_fd_sc_hd__o21ai_1
Xwire5232 net5233 VGND VGND VPWR VPWR net5232 sky130_fd_sc_hd__buf_1
XFILLER_0_47_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5254 net5255 VGND VGND VPWR VPWR net5254 sky130_fd_sc_hd__buf_1
Xwire5265 net5266 VGND VGND VPWR VPWR net5265 sky130_fd_sc_hd__buf_1
Xwire4531 net4532 VGND VGND VPWR VPWR net4531 sky130_fd_sc_hd__buf_1
Xwire5276 net5278 VGND VGND VPWR VPWR net5276 sky130_fd_sc_hd__clkbuf_1
Xwire4542 net4543 VGND VGND VPWR VPWR net4542 sky130_fd_sc_hd__buf_1
X_24159_ net739 net930 VGND VGND VPWR VPWR _04021_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5287 net5288 VGND VGND VPWR VPWR net5287 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4553 net4554 VGND VGND VPWR VPWR net4553 sky130_fd_sc_hd__buf_1
Xwire5298 matmul0.beta_pass\[2\] VGND VGND VPWR VPWR net5298 sky130_fd_sc_hd__clkbuf_1
Xwire4564 net4556 VGND VGND VPWR VPWR net4564 sky130_fd_sc_hd__clkbuf_1
Xwire4575 net4576 VGND VGND VPWR VPWR net4575 sky130_fd_sc_hd__buf_1
Xwire3830 net3831 VGND VGND VPWR VPWR net3830 sky130_fd_sc_hd__buf_1
Xwire3841 _00871_ VGND VGND VPWR VPWR net3841 sky130_fd_sc_hd__buf_1
Xwire4597 net4598 VGND VGND VPWR VPWR net4597 sky130_fd_sc_hd__buf_1
X_16981_ net6493 net6475 net6467 VGND VGND VPWR VPWR _08943_ sky130_fd_sc_hd__and3_1
Xwire3852 _12266_ VGND VGND VPWR VPWR net3852 sky130_fd_sc_hd__buf_1
Xwire3863 _11490_ VGND VGND VPWR VPWR net3863 sky130_fd_sc_hd__buf_1
XFILLER_0_101_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3874 net3875 VGND VGND VPWR VPWR net3874 sky130_fd_sc_hd__clkbuf_1
X_18720_ _10564_ _10565_ VGND VGND VPWR VPWR _10566_ sky130_fd_sc_hd__nand2_1
Xwire3885 _10930_ VGND VGND VPWR VPWR net3885 sky130_fd_sc_hd__clkbuf_1
X_15932_ _07894_ net1263 _08000_ VGND VGND VPWR VPWR _08001_ sky130_fd_sc_hd__a21oi_1
Xwire3896 _10878_ VGND VGND VPWR VPWR net3896 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_155_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18651_ _10495_ net1195 VGND VGND VPWR VPWR _10498_ sky130_fd_sc_hd__xnor2_1
X_15863_ net4075 net4068 VGND VGND VPWR VPWR _07932_ sky130_fd_sc_hd__nor2_2
X_17602_ net4015 svm0.tB\[10\] VGND VGND VPWR VPWR _09483_ sky130_fd_sc_hd__and2_1
X_14814_ net7446 net7168 net3627 VGND VGND VPWR VPWR _06924_ sky130_fd_sc_hd__a21o_1
XFILLER_0_192_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15794_ net3439 VGND VGND VPWR VPWR _07864_ sky130_fd_sc_hd__buf_1
X_18582_ net3945 _10429_ net6919 VGND VGND VPWR VPWR _10430_ sky130_fd_sc_hd__mux2_1
X_17533_ net6686 svm0.delta\[14\] _09414_ _09415_ VGND VGND VPWR VPWR _09416_ sky130_fd_sc_hd__a211o_1
X_14745_ net3616 matmul0.sin\[4\] _06832_ VGND VGND VPWR VPWR _06878_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17464_ svm0.counter\[4\] _09356_ _09357_ _09355_ VGND VGND VPWR VPWR _00395_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14676_ net7160 net7164 VGND VGND VPWR VPWR _06827_ sky130_fd_sc_hd__nor2_1
X_19203_ _11034_ _11039_ VGND VGND VPWR VPWR _11040_ sky130_fd_sc_hd__nand2_1
X_16415_ _08421_ _08413_ _08422_ VGND VGND VPWR VPWR _08477_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_95_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13627_ net7709 net3685 net2967 VGND VGND VPWR VPWR _05897_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17395_ net612 _09301_ _09299_ VGND VGND VPWR VPWR _09302_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_184_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_8__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_4_8__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_183_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19134_ net6119 net6086 VGND VGND VPWR VPWR _10971_ sky130_fd_sc_hd__xor2_2
XFILLER_0_55_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16346_ net2682 net3561 _08343_ VGND VGND VPWR VPWR _08409_ sky130_fd_sc_hd__a21oi_1
X_13558_ _05823_ _05828_ VGND VGND VPWR VPWR _05829_ sky130_fd_sc_hd__xnor2_1
Xfanout7062 net7067 VGND VGND VPWR VPWR net7062 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_132_Right_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout7073 cordic0.vec\[1\]\[4\] VGND VGND VPWR VPWR net7073 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19065_ _10900_ _10901_ VGND VGND VPWR VPWR _10902_ sky130_fd_sc_hd__nor2_1
X_16277_ net2707 _08258_ net2721 VGND VGND VPWR VPWR _08341_ sky130_fd_sc_hd__a21oi_1
X_13489_ net625 _05761_ VGND VGND VPWR VPWR _05762_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_164_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7190 net7191 VGND VGND VPWR VPWR net7190 sky130_fd_sc_hd__clkbuf_1
X_18016_ _09860_ net2550 VGND VGND VPWR VPWR _09867_ sky130_fd_sc_hd__nor2_1
X_15228_ net3451 net3487 VGND VGND VPWR VPWR _07302_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15159_ _07223_ net1884 _07232_ VGND VGND VPWR VPWR _07233_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_50_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19967_ net6166 net6093 VGND VGND VPWR VPWR _11798_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18918_ net6828 _10279_ _10710_ _10757_ net6814 VGND VGND VPWR VPWR _10758_ sky130_fd_sc_hd__a221o_1
X_19898_ net1768 _11728_ _11729_ _11730_ VGND VGND VPWR VPWR _00457_ sky130_fd_sc_hd__a31o_1
X_18849_ _10686_ _10691_ VGND VGND VPWR VPWR _10692_ sky130_fd_sc_hd__xor2_1
X_21860_ net5406 net3786 VGND VGND VPWR VPWR _01869_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20811_ net5830 net5510 VGND VGND VPWR VPWR _00827_ sky130_fd_sc_hd__nand2_1
X_21791_ _01794_ _01800_ VGND VGND VPWR VPWR _01801_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23530_ _03330_ _03331_ _03329_ VGND VGND VPWR VPWR _03398_ sky130_fd_sc_hd__o21ai_1
Xmax_length5218 matmul0.beta_pass\[11\] VGND VGND VPWR VPWR net5218 sky130_fd_sc_hd__clkbuf_1
X_20742_ _12509_ _12510_ _12512_ VGND VGND VPWR VPWR _12513_ sky130_fd_sc_hd__a21o_1
XFILLER_0_159_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length4506 net4503 VGND VGND VPWR VPWR net4506 sky130_fd_sc_hd__buf_1
Xwire8819 net8820 VGND VGND VPWR VPWR net8819 sky130_fd_sc_hd__clkbuf_1
X_23461_ net4550 net5099 VGND VGND VPWR VPWR _03330_ sky130_fd_sc_hd__nand2_1
XFILLER_0_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20673_ net1473 _12448_ net3357 VGND VGND VPWR VPWR _12450_ sky130_fd_sc_hd__a21oi_1
X_25200_ clknet_leaf_58_clk _00089_ net8710 VGND VGND VPWR VPWR matmul0.b_in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_22412_ _02382_ _02412_ VGND VGND VPWR VPWR _02414_ sky130_fd_sc_hd__nor2_1
Xwire509 _04497_ VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__buf_1
XFILLER_0_45_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23392_ _03254_ _03261_ VGND VGND VPWR VPWR _03262_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25131_ clknet_leaf_52_clk _00020_ net8805 VGND VGND VPWR VPWR svm0.tC\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22343_ _02291_ _02292_ _02293_ VGND VGND VPWR VPWR _02346_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25062_ net3732 _04806_ net4430 VGND VGND VPWR VPWR _04810_ sky130_fd_sc_hd__o21ba_1
X_22274_ _02242_ _02243_ _02199_ VGND VGND VPWR VPWR _02278_ sky130_fd_sc_hd__o21ba_1
X_24013_ net4488 _03875_ VGND VGND VPWR VPWR _03876_ sky130_fd_sc_hd__nand2_1
Xhold140 svm0.tA\[6\] VGND VGND VPWR VPWR net9093 sky130_fd_sc_hd__dlygate4sd3_1
X_21225_ _00938_ _00968_ _01232_ _01240_ VGND VGND VPWR VPWR _01241_ sky130_fd_sc_hd__o31a_1
Xhold151 matmul0.matmul_stage_inst.c\[2\] VGND VGND VPWR VPWR net9104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 svm0.vC\[12\] VGND VGND VPWR VPWR net9115 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3104 _02519_ VGND VGND VPWR VPWR net3104 sky130_fd_sc_hd__buf_1
Xhold173 svm0.tC\[12\] VGND VGND VPWR VPWR net9126 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3126 net3127 VGND VGND VPWR VPWR net3126 sky130_fd_sc_hd__clkbuf_2
Xhold184 svm0.tC\[4\] VGND VGND VPWR VPWR net9137 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3137 net3138 VGND VGND VPWR VPWR net3137 sky130_fd_sc_hd__buf_1
Xwire2403 _04527_ VGND VGND VPWR VPWR net2403 sky130_fd_sc_hd__buf_1
X_21156_ _01168_ _01171_ VGND VGND VPWR VPWR _01172_ sky130_fd_sc_hd__xnor2_1
Xhold195 matmul0.matmul_stage_inst.state\[0\] VGND VGND VPWR VPWR net9148 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3148 net3149 VGND VGND VPWR VPWR net3148 sky130_fd_sc_hd__clkbuf_1
Xwire2414 net2415 VGND VGND VPWR VPWR net2414 sky130_fd_sc_hd__clkbuf_1
Xwire3159 net3160 VGND VGND VPWR VPWR net3159 sky130_fd_sc_hd__clkbuf_1
Xwire2425 _03343_ VGND VGND VPWR VPWR net2425 sky130_fd_sc_hd__clkbuf_1
Xwire2436 net2437 VGND VGND VPWR VPWR net2436 sky130_fd_sc_hd__clkbuf_1
X_20107_ net6052 net6000 _11890_ VGND VGND VPWR VPWR _11935_ sky130_fd_sc_hd__mux2_1
Xwire1702 _02297_ VGND VGND VPWR VPWR net1702 sky130_fd_sc_hd__buf_1
X_21087_ _01062_ net1731 _01061_ VGND VGND VPWR VPWR _01103_ sky130_fd_sc_hd__and3b_1
Xwire1713 _01961_ VGND VGND VPWR VPWR net1713 sky130_fd_sc_hd__buf_1
Xwire2458 _02556_ VGND VGND VPWR VPWR net2458 sky130_fd_sc_hd__buf_1
Xwire2469 _02520_ VGND VGND VPWR VPWR net2469 sky130_fd_sc_hd__clkbuf_1
X_24915_ net8870 net137 VGND VGND VPWR VPWR _04704_ sky130_fd_sc_hd__and2b_1
X_20038_ net1404 _11867_ VGND VGND VPWR VPWR _11868_ sky130_fd_sc_hd__xnor2_2
Xwire1735 _00839_ VGND VGND VPWR VPWR net1735 sky130_fd_sc_hd__buf_1
Xwire1746 _12341_ VGND VGND VPWR VPWR net1746 sky130_fd_sc_hd__clkbuf_1
X_25895_ clknet_leaf_14_clk _00768_ net8621 VGND VGND VPWR VPWR pid_q.kp\[7\] sky130_fd_sc_hd__dfrtp_1
Xwire1757 _10921_ VGND VGND VPWR VPWR net1757 sky130_fd_sc_hd__buf_1
XFILLER_0_176_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1768 net1769 VGND VGND VPWR VPWR net1768 sky130_fd_sc_hd__buf_1
Xwire1779 _09725_ VGND VGND VPWR VPWR net1779 sky130_fd_sc_hd__buf_1
X_24846_ net7486 net372 _04327_ VGND VGND VPWR VPWR _04656_ sky130_fd_sc_hd__a21o_1
X_12860_ net4261 net1596 VGND VGND VPWR VPWR _05133_ sky130_fd_sc_hd__nor2_1
Xmax_length7121 net7118 VGND VGND VPWR VPWR net7121 sky130_fd_sc_hd__buf_1
X_24777_ net5228 net7980 VGND VGND VPWR VPWR _04604_ sky130_fd_sc_hd__and2b_1
X_12791_ _05063_ VGND VGND VPWR VPWR _05064_ sky130_fd_sc_hd__buf_1
XFILLER_0_179_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21989_ _01991_ _01996_ VGND VGND VPWR VPWR _01997_ sky130_fd_sc_hd__and2b_1
Xmax_length7154 matmul0.sin\[6\] VGND VGND VPWR VPWR net7154 sky130_fd_sc_hd__clkbuf_1
X_14530_ net726 _06703_ VGND VGND VPWR VPWR _06709_ sky130_fd_sc_hd__and2_1
X_23728_ _03512_ _03514_ _03513_ VGND VGND VPWR VPWR _03594_ sky130_fd_sc_hd__o21a_1
Xmax_length6453 net6454 VGND VGND VPWR VPWR net6453 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14461_ net9086 _06543_ _06649_ net6453 VGND VGND VPWR VPWR _00100_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23659_ net4615 net4934 VGND VGND VPWR VPWR _03526_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16200_ net1250 _08264_ VGND VGND VPWR VPWR _08265_ sky130_fd_sc_hd__xnor2_1
X_13412_ net731 _05633_ _05684_ VGND VGND VPWR VPWR _05685_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_138_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17180_ net6850 net1820 _09130_ VGND VGND VPWR VPWR _09132_ sky130_fd_sc_hd__or3_1
X_14392_ net8163 net3635 VGND VGND VPWR VPWR _06597_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16131_ net2645 net2659 _08194_ _08195_ VGND VGND VPWR VPWR _08197_ sky130_fd_sc_hd__o211ai_1
X_13343_ net7869 net4254 VGND VGND VPWR VPWR _05616_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25329_ clknet_leaf_80_clk _00212_ net8464 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.f\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16062_ _08025_ _08030_ _08128_ VGND VGND VPWR VPWR _08129_ sky130_fd_sc_hd__o21a_1
X_13274_ _05538_ _05545_ _05546_ VGND VGND VPWR VPWR _05547_ sky130_fd_sc_hd__or3_1
Xwire5040 net5042 VGND VGND VPWR VPWR net5040 sky130_fd_sc_hd__buf_1
XFILLER_0_20_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5051 net5052 VGND VGND VPWR VPWR net5051 sky130_fd_sc_hd__clkbuf_1
X_15013_ _07086_ VGND VGND VPWR VPWR _07087_ sky130_fd_sc_hd__buf_1
Xwire5062 net5063 VGND VGND VPWR VPWR net5062 sky130_fd_sc_hd__buf_1
XFILLER_0_103_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5084 net5090 VGND VGND VPWR VPWR net5084 sky130_fd_sc_hd__buf_1
Xwire4350 net4351 VGND VGND VPWR VPWR net4350 sky130_fd_sc_hd__clkbuf_1
X_19821_ net953 _11654_ VGND VGND VPWR VPWR _11655_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_102_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4372 net4373 VGND VGND VPWR VPWR net4372 sky130_fd_sc_hd__buf_1
XFILLER_0_166_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4394 net4395 VGND VGND VPWR VPWR net4394 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3660 net3661 VGND VGND VPWR VPWR net3660 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3671 net3672 VGND VGND VPWR VPWR net3671 sky130_fd_sc_hd__clkbuf_1
X_19752_ net6050 net6030 net3136 net6088 VGND VGND VPWR VPWR _11587_ sky130_fd_sc_hd__a211o_1
Xwire3682 net3683 VGND VGND VPWR VPWR net3682 sky130_fd_sc_hd__buf_1
X_16964_ _08842_ _08926_ net6522 VGND VGND VPWR VPWR _08927_ sky130_fd_sc_hd__mux2_1
Xwire3693 _04897_ VGND VGND VPWR VPWR net3693 sky130_fd_sc_hd__buf_1
X_18703_ _10545_ _10548_ VGND VGND VPWR VPWR _10549_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_142_Left_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2970 _05054_ VGND VGND VPWR VPWR net2970 sky130_fd_sc_hd__buf_1
X_15915_ net884 _07983_ VGND VGND VPWR VPWR _07984_ sky130_fd_sc_hd__or2_1
Xwire2981 net2983 VGND VGND VPWR VPWR net2981 sky130_fd_sc_hd__buf_1
X_19683_ _11164_ _11518_ net6176 VGND VGND VPWR VPWR _11519_ sky130_fd_sc_hd__mux2_1
Xwire2992 _04890_ VGND VGND VPWR VPWR net2992 sky130_fd_sc_hd__buf_1
X_16895_ net6369 _08858_ net6396 VGND VGND VPWR VPWR _08859_ sky130_fd_sc_hd__o21ba_1
X_18634_ net6827 net6862 _10480_ VGND VGND VPWR VPWR _10481_ sky130_fd_sc_hd__o21ai_1
X_15846_ _07819_ _07915_ VGND VGND VPWR VPWR _07916_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18565_ net663 net659 _10411_ _10412_ VGND VGND VPWR VPWR _10413_ sky130_fd_sc_hd__a31o_1
X_12989_ _05253_ _05261_ VGND VGND VPWR VPWR _05262_ sky130_fd_sc_hd__xnor2_2
X_15777_ net4138 net4131 net4198 net4197 VGND VGND VPWR VPWR _07847_ sky130_fd_sc_hd__o22a_1
X_17516_ net3275 _09401_ net6657 VGND VGND VPWR VPWR _09402_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14728_ net7437 net7162 net3697 VGND VGND VPWR VPWR _06865_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18496_ net1208 net1441 _10327_ VGND VGND VPWR VPWR _10345_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17447_ _09341_ _09342_ VGND VGND VPWR VPWR _09343_ sky130_fd_sc_hd__nand2_1
X_14659_ net3628 VGND VGND VPWR VPWR _06814_ sky130_fd_sc_hd__buf_1
XFILLER_0_144_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_151_Left_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17378_ svm0.delta\[3\] _09284_ VGND VGND VPWR VPWR _09288_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19117_ net6311 net3212 _10811_ VGND VGND VPWR VPWR _10954_ sky130_fd_sc_hd__o21a_1
X_16329_ _08319_ _08320_ _08321_ VGND VGND VPWR VPWR _08392_ sky130_fd_sc_hd__o21a_1
XFILLER_0_125_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19048_ net6356 _10813_ VGND VGND VPWR VPWR _10885_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5490 net5501 VGND VGND VPWR VPWR net5490 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21010_ net1185 _01024_ VGND VGND VPWR VPWR _01026_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_160_Left_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1009 _04569_ VGND VGND VPWR VPWR net1009 sky130_fd_sc_hd__buf_1
X_22961_ net5314 net3064 _02848_ net8910 VGND VGND VPWR VPWR _00647_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24700_ net5299 _04536_ VGND VGND VPWR VPWR _04537_ sky130_fd_sc_hd__xnor2_1
X_21912_ net5977 pid_d.prev_int\[8\] VGND VGND VPWR VPWR _01920_ sky130_fd_sc_hd__xor2_1
X_25680_ clknet_leaf_0_clk _00553_ net8409 VGND VGND VPWR VPWR pid_d.curr_error\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_22892_ _02017_ _02779_ net5357 VGND VGND VPWR VPWR _02786_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_78_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24631_ net4514 _04479_ _04480_ _04485_ VGND VGND VPWR VPWR _04486_ sky130_fd_sc_hd__o211a_1
X_21843_ _01756_ _01758_ _01851_ VGND VGND VPWR VPWR _01852_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_172_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24562_ net4545 _04417_ VGND VGND VPWR VPWR _04418_ sky130_fd_sc_hd__nand2_1
X_21774_ _01782_ _01783_ VGND VGND VPWR VPWR _01784_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23513_ _03379_ net745 VGND VGND VPWR VPWR _03382_ sky130_fd_sc_hd__xnor2_1
Xwire8616 net8615 VGND VGND VPWR VPWR net8616 sky130_fd_sc_hd__clkbuf_2
X_20725_ _12492_ _12496_ _12491_ VGND VGND VPWR VPWR _12497_ sky130_fd_sc_hd__mux2_1
X_24493_ net4894 net4871 VGND VGND VPWR VPWR _04350_ sky130_fd_sc_hd__or2_1
Xwire8638 net8639 VGND VGND VPWR VPWR net8638 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7904 svm0.periodTop\[2\] VGND VGND VPWR VPWR net7904 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23444_ net7466 net545 _03311_ net7526 net3056 VGND VGND VPWR VPWR _03314_ sky130_fd_sc_hd__a221o_1
Xwire7915 net7916 VGND VGND VPWR VPWR net7915 sky130_fd_sc_hd__clkbuf_1
Xwire306 net307 VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__clkbuf_1
Xwire7926 net7927 VGND VGND VPWR VPWR net7926 sky130_fd_sc_hd__clkbuf_1
X_20656_ _12422_ _12432_ _12433_ VGND VGND VPWR VPWR _12434_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length3613 net3614 VGND VGND VPWR VPWR net3613 sky130_fd_sc_hd__buf_1
XFILLER_0_162_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire317 _08236_ VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire328 _04384_ VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__buf_1
Xwire7937 net7938 VGND VGND VPWR VPWR net7937 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7948 net7942 VGND VGND VPWR VPWR net7948 sky130_fd_sc_hd__buf_1
Xwire339 net340 VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__buf_1
XFILLER_0_191_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7959 net7960 VGND VGND VPWR VPWR net7959 sky130_fd_sc_hd__clkbuf_1
X_23375_ _03241_ _03244_ VGND VGND VPWR VPWR _03245_ sky130_fd_sc_hd__xnor2_1
X_20587_ _12362_ _12369_ VGND VGND VPWR VPWR _12370_ sky130_fd_sc_hd__and2b_1
X_25114_ pid_d.prev_int\[2\] net2392 net1992 net9079 VGND VGND VPWR VPWR _00795_ sky130_fd_sc_hd__a22o_1
X_22326_ pid_d.curr_int\[12\] net3844 net2489 _02329_ VGND VGND VPWR VPWR _00531_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length2956 _05346_ VGND VGND VPWR VPWR net2956 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25045_ pid_q.out\[7\] net5178 VGND VGND VPWR VPWR _04796_ sky130_fd_sc_hd__xnor2_1
X_22257_ pid_d.curr_int\[11\] net3843 net2487 _02261_ VGND VGND VPWR VPWR _00530_
+ sky130_fd_sc_hd__a22o_1
X_21208_ _01223_ net1734 net1183 VGND VGND VPWR VPWR _01224_ sky130_fd_sc_hd__a21bo_1
X_22188_ net1710 _02057_ VGND VGND VPWR VPWR _02193_ sky130_fd_sc_hd__nand2_1
Xwire2200 net2201 VGND VGND VPWR VPWR net2200 sky130_fd_sc_hd__clkbuf_1
Xwire2211 net2212 VGND VGND VPWR VPWR net2211 sky130_fd_sc_hd__buf_1
Xwire2222 net2223 VGND VGND VPWR VPWR net2222 sky130_fd_sc_hd__buf_1
X_21139_ _01153_ _01154_ VGND VGND VPWR VPWR _01155_ sky130_fd_sc_hd__or2_1
Xwire2233 _07377_ VGND VGND VPWR VPWR net2233 sky130_fd_sc_hd__buf_1
Xwire2244 _07156_ VGND VGND VPWR VPWR net2244 sky130_fd_sc_hd__clkbuf_1
Xwire2255 _07006_ VGND VGND VPWR VPWR net2255 sky130_fd_sc_hd__clkbuf_1
Xwire2266 net2267 VGND VGND VPWR VPWR net2266 sky130_fd_sc_hd__buf_1
Xwire1521 _07992_ VGND VGND VPWR VPWR net1521 sky130_fd_sc_hd__buf_1
X_13961_ net7648 net1331 _06187_ _06218_ net7681 VGND VGND VPWR VPWR _06226_ sky130_fd_sc_hd__a32o_1
Xwire1532 net1533 VGND VGND VPWR VPWR net1532 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1543 _07349_ VGND VGND VPWR VPWR net1543 sky130_fd_sc_hd__buf_1
Xwire2288 net2289 VGND VGND VPWR VPWR net2288 sky130_fd_sc_hd__buf_1
Xwire2299 _05420_ VGND VGND VPWR VPWR net2299 sky130_fd_sc_hd__clkbuf_1
Xwire1554 net1555 VGND VGND VPWR VPWR net1554 sky130_fd_sc_hd__buf_1
Xwire1565 net1566 VGND VGND VPWR VPWR net1565 sky130_fd_sc_hd__clkbuf_1
X_12912_ net850 _05168_ _05169_ VGND VGND VPWR VPWR _05185_ sky130_fd_sc_hd__nand3_1
X_15700_ _07698_ _07699_ _07770_ VGND VGND VPWR VPWR _07771_ sky130_fd_sc_hd__o21a_1
Xwire1576 _05555_ VGND VGND VPWR VPWR net1576 sky130_fd_sc_hd__clkbuf_1
X_16680_ _08710_ _08706_ _08711_ VGND VGND VPWR VPWR _08712_ sky130_fd_sc_hd__a21o_1
X_25878_ clknet_leaf_14_clk _00751_ net8621 VGND VGND VPWR VPWR pid_q.ki\[6\] sky130_fd_sc_hd__dfrtp_1
X_13892_ net283 _06156_ _06157_ VGND VGND VPWR VPWR _06158_ sky130_fd_sc_hd__o21ai_1
Xwire1587 net1588 VGND VGND VPWR VPWR net1587 sky130_fd_sc_hd__buf_1
Xwire1598 net1599 VGND VGND VPWR VPWR net1598 sky130_fd_sc_hd__clkbuf_2
X_24829_ net5072 _04642_ net2000 net1363 VGND VGND VPWR VPWR _00716_ sky130_fd_sc_hd__a22o_1
XFILLER_0_158_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12843_ _05107_ _05114_ _05115_ VGND VGND VPWR VPWR _05116_ sky130_fd_sc_hd__and3_1
X_15631_ _07691_ _07702_ VGND VGND VPWR VPWR _07703_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15562_ _07627_ _07634_ VGND VGND VPWR VPWR _07635_ sky130_fd_sc_hd__xnor2_1
X_18350_ _10147_ _10199_ _10200_ net815 VGND VGND VPWR VPWR _10201_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12774_ _05038_ _05046_ VGND VGND VPWR VPWR _05047_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_51_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17301_ net6685 VGND VGND VPWR VPWR _09215_ sky130_fd_sc_hd__inv_2
X_14513_ net7313 net5267 _06685_ VGND VGND VPWR VPWR _06694_ sky130_fd_sc_hd__or3_1
XFILLER_0_51_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15493_ _07543_ _07546_ _07402_ VGND VGND VPWR VPWR _07566_ sky130_fd_sc_hd__a21o_1
X_18281_ net2546 _10062_ net2545 VGND VGND VPWR VPWR _10132_ sky130_fd_sc_hd__a21oi_1
Xmax_length6294 net6291 VGND VGND VPWR VPWR net6294 sky130_fd_sc_hd__buf_1
X_14444_ net8180 net3634 VGND VGND VPWR VPWR _06637_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17232_ _09178_ _09179_ _09162_ VGND VGND VPWR VPWR _09180_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_182_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17163_ _09113_ _09115_ VGND VGND VPWR VPWR _09116_ sky130_fd_sc_hd__xnor2_1
Xwire840 _06062_ VGND VGND VPWR VPWR net840 sky130_fd_sc_hd__buf_1
XFILLER_0_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14375_ _06584_ VGND VGND VPWR VPWR _00079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire851 _05019_ VGND VGND VPWR VPWR net851 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_10_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16114_ _08178_ _08179_ _07932_ VGND VGND VPWR VPWR _08180_ sky130_fd_sc_hd__a21oi_1
Xwire862 _01015_ VGND VGND VPWR VPWR net862 sky130_fd_sc_hd__buf_1
XFILLER_0_101_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13326_ net7710 net1605 net1339 net7687 VGND VGND VPWR VPWR _05599_ sky130_fd_sc_hd__a22o_1
Xwire873 _10725_ VGND VGND VPWR VPWR net873 sky130_fd_sc_hd__buf_1
Xwire884 net885 VGND VGND VPWR VPWR net884 sky130_fd_sc_hd__buf_1
XFILLER_0_52_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17094_ _09050_ VGND VGND VPWR VPWR _09051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire895 net896 VGND VGND VPWR VPWR net895 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_51_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16045_ net1518 _08047_ net1520 VGND VGND VPWR VPWR _08112_ sky130_fd_sc_hd__a21bo_1
X_13257_ net6677 net5193 net6672 VGND VGND VPWR VPWR _05530_ sky130_fd_sc_hd__and3b_1
XFILLER_0_86_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13188_ _05457_ _05460_ VGND VGND VPWR VPWR _05461_ sky130_fd_sc_hd__xnor2_2
Xwire4180 _06995_ VGND VGND VPWR VPWR net4180 sky130_fd_sc_hd__buf_1
X_19804_ net3174 _11634_ _11635_ _11637_ VGND VGND VPWR VPWR _11638_ sky130_fd_sc_hd__o211a_1
Xwire4191 net4192 VGND VGND VPWR VPWR net4191 sky130_fd_sc_hd__buf_1
X_17996_ net7004 _09846_ net2555 VGND VGND VPWR VPWR _09847_ sky130_fd_sc_hd__or3b_1
XFILLER_0_159_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3490 net3491 VGND VGND VPWR VPWR net3490 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19735_ _11560_ _11561_ _11564_ _11508_ _11569_ VGND VGND VPWR VPWR _11570_ sky130_fd_sc_hd__o221a_1
X_16947_ net2284 VGND VGND VPWR VPWR _08911_ sky130_fd_sc_hd__buf_1
XFILLER_0_159_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19666_ net3201 _11501_ _11409_ VGND VGND VPWR VPWR _11502_ sky130_fd_sc_hd__a21o_1
X_16878_ net6061 net6019 net6501 VGND VGND VPWR VPWR _08842_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18617_ net2128 _10462_ _10463_ VGND VGND VPWR VPWR _10464_ sky130_fd_sc_hd__o21ai_2
X_15829_ net3565 _07898_ net2221 net2821 VGND VGND VPWR VPWR _07899_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_149_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19597_ _11387_ _11430_ _11432_ _11433_ net6071 VGND VGND VPWR VPWR _11434_ sky130_fd_sc_hd__a311o_1
XFILLER_0_126_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18548_ _10395_ _10396_ VGND VGND VPWR VPWR _10397_ sky130_fd_sc_hd__nor2_1
XFILLER_0_191_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18479_ net1208 net1441 _10327_ VGND VGND VPWR VPWR _10329_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20510_ net7010 net6983 net6962 net6938 net6514 net6490 VGND VGND VPWR VPWR _12297_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21490_ net1049 _01502_ VGND VGND VPWR VPWR _01503_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20441_ net950 _12234_ VGND VGND VPWR VPWR _12235_ sky130_fd_sc_hd__xnor2_1
Xmax_length2208 net2209 VGND VGND VPWR VPWR net2208 sky130_fd_sc_hd__buf_1
X_23160_ net5064 net4735 VGND VGND VPWR VPWR _03030_ sky130_fd_sc_hd__nand2_1
X_20372_ net6508 _12109_ VGND VGND VPWR VPWR _12171_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22111_ net802 _02079_ _02070_ VGND VGND VPWR VPWR _02117_ sky130_fd_sc_hd__a21o_1
XFILLER_0_140_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23091_ _02953_ _02960_ VGND VGND VPWR VPWR _02961_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_2_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22042_ _02043_ _02048_ VGND VGND VPWR VPWR _02049_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25801_ clknet_leaf_30_clk _00674_ net8677 VGND VGND VPWR VPWR pid_q.curr_int\[9\]
+ sky130_fd_sc_hd__dfrtp_2
X_23993_ _03854_ _03855_ VGND VGND VPWR VPWR _03857_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25732_ clknet_leaf_9_clk _00605_ net8560 VGND VGND VPWR VPWR pid_d.ki\[6\] sky130_fd_sc_hd__dfrtp_1
X_22944_ pid_d.out\[14\] net2468 _02832_ net4331 VGND VGND VPWR VPWR _02833_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25663_ clknet_leaf_121_clk _00536_ net8396 VGND VGND VPWR VPWR pid_d.prev_error\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_22875_ net5360 net5978 VGND VGND VPWR VPWR _02771_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24614_ net1649 _04436_ VGND VGND VPWR VPWR _04469_ sky130_fd_sc_hd__nor2_1
X_21826_ _01833_ _01834_ VGND VGND VPWR VPWR _01835_ sky130_fd_sc_hd__xnor2_1
X_25594_ clknet_leaf_106_clk _00467_ net8356 VGND VGND VPWR VPWR cordic0.slte0.opB\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24545_ _04393_ _04396_ _04397_ _04400_ VGND VGND VPWR VPWR _04401_ sky130_fd_sc_hd__a211o_1
X_21757_ _01763_ _01766_ VGND VGND VPWR VPWR _01767_ sky130_fd_sc_hd__xnor2_2
Xwire8402 net8403 VGND VGND VPWR VPWR net8402 sky130_fd_sc_hd__buf_1
Xwire8413 net8410 VGND VGND VPWR VPWR net8413 sky130_fd_sc_hd__buf_1
Xwire8424 net8425 VGND VGND VPWR VPWR net8424 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout7628 net7633 VGND VGND VPWR VPWR net7628 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20708_ _12479_ _12480_ VGND VGND VPWR VPWR _12481_ sky130_fd_sc_hd__xnor2_2
X_24476_ _04331_ _04332_ VGND VGND VPWR VPWR _04333_ sky130_fd_sc_hd__nand2_1
Xfanout6905 cordic0.vec\[1\]\[11\] VGND VGND VPWR VPWR net6905 sky130_fd_sc_hd__buf_1
Xwire8446 net8449 VGND VGND VPWR VPWR net8446 sky130_fd_sc_hd__clkbuf_1
X_21688_ _01577_ _01579_ _01575_ VGND VGND VPWR VPWR _01699_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_164_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23427_ _03264_ net1167 VGND VGND VPWR VPWR _03297_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7756 net7757 VGND VGND VPWR VPWR net7756 sky130_fd_sc_hd__clkbuf_1
X_20639_ net6755 _12417_ net3305 VGND VGND VPWR VPWR _12418_ sky130_fd_sc_hd__mux2_1
Xwire158 net159 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__buf_1
Xwire7767 net7763 VGND VGND VPWR VPWR net7767 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7778 net7779 VGND VGND VPWR VPWR net7778 sky130_fd_sc_hd__buf_1
Xwire169 net170 VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_1
Xwire7789 net7790 VGND VGND VPWR VPWR net7789 sky130_fd_sc_hd__buf_1
X_14160_ _06401_ _06420_ VGND VGND VPWR VPWR _06421_ sky130_fd_sc_hd__xnor2_2
Xmax_length2731 net2733 VGND VGND VPWR VPWR net2731 sky130_fd_sc_hd__clkbuf_1
X_23358_ _03216_ _03227_ VGND VGND VPWR VPWR _03228_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13111_ net7822 _05053_ _05054_ VGND VGND VPWR VPWR _05384_ sky130_fd_sc_hd__and3_1
X_22309_ _02304_ _02312_ VGND VGND VPWR VPWR _02313_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_131_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14091_ _06284_ _06287_ _06353_ VGND VGND VPWR VPWR _06354_ sky130_fd_sc_hd__o21ai_1
X_23289_ _03147_ _03157_ VGND VGND VPWR VPWR _03159_ sky130_fd_sc_hd__nor2_1
X_25028_ _03671_ _04774_ net4457 VGND VGND VPWR VPWR _04781_ sky130_fd_sc_hd__o21ba_1
X_13042_ _05313_ _05314_ _05203_ VGND VGND VPWR VPWR _05315_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17850_ net7043 net3347 VGND VGND VPWR VPWR _09701_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2030 net2031 VGND VGND VPWR VPWR net2030 sky130_fd_sc_hd__clkbuf_1
Xwire2041 _02559_ VGND VGND VPWR VPWR net2041 sky130_fd_sc_hd__clkbuf_1
X_16801_ _08790_ VGND VGND VPWR VPWR _00299_ sky130_fd_sc_hd__clkbuf_1
Xwire2052 net2053 VGND VGND VPWR VPWR net2052 sky130_fd_sc_hd__clkbuf_2
Xwire2063 _01798_ VGND VGND VPWR VPWR net2063 sky130_fd_sc_hd__dlymetal6s2s_1
X_17781_ net7090 net7104 VGND VGND VPWR VPWR _09632_ sky130_fd_sc_hd__and2b_1
Xwire2074 _01046_ VGND VGND VPWR VPWR net2074 sky130_fd_sc_hd__clkbuf_2
X_14993_ net3603 net3521 _07064_ VGND VGND VPWR VPWR _07067_ sky130_fd_sc_hd__or3b_1
Xwire1340 net1341 VGND VGND VPWR VPWR net1340 sky130_fd_sc_hd__buf_1
Xwire2085 _12294_ VGND VGND VPWR VPWR net2085 sky130_fd_sc_hd__clkbuf_1
Xwire1351 _04921_ VGND VGND VPWR VPWR net1351 sky130_fd_sc_hd__buf_1
Xwire2096 _11694_ VGND VGND VPWR VPWR net2096 sky130_fd_sc_hd__buf_1
X_19520_ _11284_ _11285_ _11298_ VGND VGND VPWR VPWR _11357_ sky130_fd_sc_hd__or3_1
Xwire1362 _04702_ VGND VGND VPWR VPWR net1362 sky130_fd_sc_hd__buf_1
X_16732_ _08754_ VGND VGND VPWR VPWR _00266_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13944_ _06165_ _06209_ VGND VGND VPWR VPWR _06210_ sky130_fd_sc_hd__xor2_1
XFILLER_0_163_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1373 _04510_ VGND VGND VPWR VPWR net1373 sky130_fd_sc_hd__buf_1
Xwire1384 _03408_ VGND VGND VPWR VPWR net1384 sky130_fd_sc_hd__buf_1
Xwire1395 _12396_ VGND VGND VPWR VPWR net1395 sky130_fd_sc_hd__buf_1
X_19451_ _10982_ net2520 _11287_ VGND VGND VPWR VPWR _11288_ sky130_fd_sc_hd__o21a_1
X_13875_ net530 _06141_ VGND VGND VPWR VPWR _06142_ sky130_fd_sc_hd__xnor2_2
X_16663_ _08697_ VGND VGND VPWR VPWR _00254_ sky130_fd_sc_hd__clkbuf_1
X_18402_ net1073 _10157_ net1211 VGND VGND VPWR VPWR _10253_ sky130_fd_sc_hd__o21ba_1
X_12826_ net7784 _04919_ _05040_ _05041_ VGND VGND VPWR VPWR _05099_ sky130_fd_sc_hd__a22o_1
X_15614_ net4076 net4069 VGND VGND VPWR VPWR _07686_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19382_ net6152 _11047_ VGND VGND VPWR VPWR _11219_ sky130_fd_sc_hd__xnor2_1
X_16594_ net5185 net4253 VGND VGND VPWR VPWR _08645_ sky130_fd_sc_hd__and2_1
XFILLER_0_96_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18333_ _10106_ _10107_ _10182_ _10183_ VGND VGND VPWR VPWR _10184_ sky130_fd_sc_hd__a31oi_1
X_12757_ _04979_ _05029_ VGND VGND VPWR VPWR _05030_ sky130_fd_sc_hd__xor2_2
X_15545_ net2713 net3494 net3423 net2689 VGND VGND VPWR VPWR _07618_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15476_ net1875 _07544_ _07546_ VGND VGND VPWR VPWR _07550_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18264_ _10093_ _10113_ _10114_ VGND VGND VPWR VPWR _10115_ sky130_fd_sc_hd__nand3_1
X_12688_ net7948 _04960_ VGND VGND VPWR VPWR _04961_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17215_ _08835_ _09006_ VGND VGND VPWR VPWR _09164_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14427_ _06624_ VGND VGND VPWR VPWR _00091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18195_ _09793_ net3936 net6973 VGND VGND VPWR VPWR _10046_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14358_ net7271 net1303 net2895 net5351 _06570_ VGND VGND VPWR VPWR _06571_ sky130_fd_sc_hd__a221o_1
X_17146_ _09083_ _09084_ VGND VGND VPWR VPWR _09100_ sky130_fd_sc_hd__nor2_1
Xwire670 _09116_ VGND VGND VPWR VPWR net670 sky130_fd_sc_hd__buf_1
Xwire681 _05808_ VGND VGND VPWR VPWR net681 sky130_fd_sc_hd__buf_1
XFILLER_0_141_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire692 net693 VGND VGND VPWR VPWR net692 sky130_fd_sc_hd__buf_1
XFILLER_0_13_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13309_ _05495_ _05496_ _05497_ VGND VGND VPWR VPWR _05582_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17077_ net2609 _09034_ VGND VGND VPWR VPWR _09035_ sky130_fd_sc_hd__nand2_1
X_14289_ net78 net2901 net2264 net7771 VGND VGND VPWR VPWR _00058_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16028_ net2649 net2624 VGND VGND VPWR VPWR _08095_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17979_ net1214 _09826_ _09827_ _09829_ VGND VGND VPWR VPWR _09830_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_58_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19718_ _11488_ _11542_ VGND VGND VPWR VPWR _11553_ sky130_fd_sc_hd__or2_1
X_20990_ _00880_ _01005_ VGND VGND VPWR VPWR _01006_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19649_ _10344_ net568 VGND VGND VPWR VPWR _11486_ sky130_fd_sc_hd__nor2_1
XFILLER_0_177_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22660_ pid_d.mult0.b\[13\] net3775 VGND VGND VPWR VPWR _02615_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21611_ _01506_ _01622_ _01621_ net1179 VGND VGND VPWR VPWR _01623_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_118_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22591_ net5968 net2044 net3093 net1698 VGND VGND VPWR VPWR _00557_ sky130_fd_sc_hd__a22o_1
XFILLER_0_192_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24330_ _04187_ _04174_ _04188_ VGND VGND VPWR VPWR _04189_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_7_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21542_ _01501_ net1049 _01553_ VGND VGND VPWR VPWR _01554_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_29_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire7019 net7021 VGND VGND VPWR VPWR net7019 sky130_fd_sc_hd__buf_1
XFILLER_0_62_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24261_ net793 _04095_ _04120_ VGND VGND VPWR VPWR _04121_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21473_ _01484_ _01485_ VGND VGND VPWR VPWR _01486_ sky130_fd_sc_hd__xor2_1
Xwire6307 net6308 VGND VGND VPWR VPWR net6307 sky130_fd_sc_hd__clkbuf_1
Xwire6329 net6330 VGND VGND VPWR VPWR net6329 sky130_fd_sc_hd__clkbuf_1
X_23212_ _03075_ _03078_ _03081_ VGND VGND VPWR VPWR _03082_ sky130_fd_sc_hd__o21a_1
Xmax_length2038 net2039 VGND VGND VPWR VPWR net2038 sky130_fd_sc_hd__buf_1
XFILLER_0_15_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20424_ _12205_ _12210_ _12219_ VGND VGND VPWR VPWR _12220_ sky130_fd_sc_hd__a21oi_1
X_24192_ _04051_ _04001_ _04052_ VGND VGND VPWR VPWR _04053_ sky130_fd_sc_hd__a21o_1
Xwire4905 net4906 VGND VGND VPWR VPWR net4905 sky130_fd_sc_hd__buf_1
Xmax_length1337 net1338 VGND VGND VPWR VPWR net1337 sky130_fd_sc_hd__clkbuf_1
X_23143_ _03011_ _03012_ VGND VGND VPWR VPWR _03013_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20355_ _12151_ _12155_ VGND VGND VPWR VPWR _12156_ sky130_fd_sc_hd__nand2_1
Xwire4927 net4929 VGND VGND VPWR VPWR net4927 sky130_fd_sc_hd__buf_1
XFILLER_0_140_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4938 net4933 VGND VGND VPWR VPWR net4938 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4949 net4950 VGND VGND VPWR VPWR net4949 sky130_fd_sc_hd__buf_1
XFILLER_0_105_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23074_ _02940_ _02943_ VGND VGND VPWR VPWR _02944_ sky130_fd_sc_hd__xnor2_2
X_20286_ _09032_ net1485 VGND VGND VPWR VPWR _12092_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22025_ net5721 net5464 VGND VGND VPWR VPWR _02032_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold11 svm0.vC\[9\] VGND VGND VPWR VPWR net8964 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 cordic0.cos\[6\] VGND VGND VPWR VPWR net8975 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 pid_q.target\[1\] VGND VGND VPWR VPWR net8986 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 cordic0.cos\[5\] VGND VGND VPWR VPWR net8997 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 matmul0.matmul_stage_inst.d\[7\] VGND VGND VPWR VPWR net9008 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_length8900 net8901 VGND VGND VPWR VPWR net8900 sky130_fd_sc_hd__clkbuf_1
Xhold66 matmul0.matmul_stage_inst.d\[4\] VGND VGND VPWR VPWR net9019 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 svm0.vC\[8\] VGND VGND VPWR VPWR net9030 sky130_fd_sc_hd__dlygate4sd3_1
X_23976_ _03737_ _03743_ _03744_ VGND VGND VPWR VPWR _03840_ sky130_fd_sc_hd__o21a_1
Xhold88 svm0.counter\[15\] VGND VGND VPWR VPWR net9041 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 matmul0.matmul_stage_inst.d\[1\] VGND VGND VPWR VPWR net9052 sky130_fd_sc_hd__dlygate4sd3_1
X_25715_ clknet_leaf_9_clk _00588_ net8559 VGND VGND VPWR VPWR pid_d.mult0.a\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_22927_ net5339 net2467 _02816_ net4333 _02817_ VGND VGND VPWR VPWR _02818_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13660_ _05927_ _05929_ VGND VGND VPWR VPWR _05930_ sky130_fd_sc_hd__nand2_1
XFILLER_0_196_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25646_ clknet_leaf_1_clk _00519_ net8403 VGND VGND VPWR VPWR pid_d.curr_int\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_22858_ net4337 _02754_ _02755_ net523 net4359 VGND VGND VPWR VPWR _02756_ sky130_fd_sc_hd__a32o_1
X_12611_ _04885_ VGND VGND VPWR VPWR _04886_ sky130_fd_sc_hd__clkbuf_2
X_21809_ pid_d.prev_int\[6\] VGND VGND VPWR VPWR _01818_ sky130_fd_sc_hd__inv_2
X_13591_ _05858_ net534 _05859_ _05860_ VGND VGND VPWR VPWR _05861_ sky130_fd_sc_hd__o31a_1
Xclkbuf_leaf_117_clk clknet_4_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_117_clk
+ sky130_fd_sc_hd__clkbuf_16
X_25577_ clknet_leaf_98_clk _00450_ net8383 VGND VGND VPWR VPWR cordic0.sin\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_22789_ _02702_ VGND VGND VPWR VPWR _00621_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15330_ _07402_ _07366_ _07367_ VGND VGND VPWR VPWR _07404_ sky130_fd_sc_hd__or3_1
Xwire8210 net8211 VGND VGND VPWR VPWR net8210 sky130_fd_sc_hd__clkbuf_1
X_24528_ pid_q.prev_error\[13\] net5166 VGND VGND VPWR VPWR _04385_ sky130_fd_sc_hd__xnor2_1
Xwire8221 net8222 VGND VGND VPWR VPWR net8221 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout7436 net7443 VGND VGND VPWR VPWR net7436 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8232 net29 VGND VGND VPWR VPWR net8232 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8243 net8244 VGND VGND VPWR VPWR net8243 sky130_fd_sc_hd__clkbuf_1
Xwire8254 net8255 VGND VGND VPWR VPWR net8254 sky130_fd_sc_hd__clkbuf_1
Xwire7520 pid_q.state\[2\] VGND VGND VPWR VPWR net7520 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout7458 matmul0.op\[0\] VGND VGND VPWR VPWR net7458 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15261_ _07267_ _07299_ _07334_ VGND VGND VPWR VPWR _07335_ sky130_fd_sc_hd__a21oi_1
Xwire8265 net8266 VGND VGND VPWR VPWR net8265 sky130_fd_sc_hd__clkbuf_1
X_24459_ net792 _04316_ VGND VGND VPWR VPWR _04317_ sky130_fd_sc_hd__xnor2_1
Xwire7531 net7532 VGND VGND VPWR VPWR net7531 sky130_fd_sc_hd__clkbuf_2
Xwire8276 net8277 VGND VGND VPWR VPWR net8276 sky130_fd_sc_hd__clkbuf_1
Xwire8287 net8288 VGND VGND VPWR VPWR net8287 sky130_fd_sc_hd__clkbuf_1
Xwire7542 net7543 VGND VGND VPWR VPWR net7542 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8298 net8299 VGND VGND VPWR VPWR net8298 sky130_fd_sc_hd__clkbuf_1
Xmax_length3240 net3241 VGND VGND VPWR VPWR net3240 sky130_fd_sc_hd__buf_1
Xwire7553 net7554 VGND VGND VPWR VPWR net7553 sky130_fd_sc_hd__clkbuf_1
X_14212_ net7602 net1119 VGND VGND VPWR VPWR _06471_ sky130_fd_sc_hd__nand2_1
X_17000_ _08960_ _08961_ VGND VGND VPWR VPWR _08962_ sky130_fd_sc_hd__nand2_1
Xwire7564 net7565 VGND VGND VPWR VPWR net7564 sky130_fd_sc_hd__clkbuf_1
Xmax_length3262 net3263 VGND VGND VPWR VPWR net3262 sky130_fd_sc_hd__buf_1
Xwire7575 net7576 VGND VGND VPWR VPWR net7575 sky130_fd_sc_hd__clkbuf_1
X_15192_ _07259_ _07257_ VGND VGND VPWR VPWR _07266_ sky130_fd_sc_hd__xnor2_1
Xwire6841 net6839 VGND VGND VPWR VPWR net6841 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_85_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7586 net7587 VGND VGND VPWR VPWR net7586 sky130_fd_sc_hd__clkbuf_1
Xwire7597 matmul0.a_in\[10\] VGND VGND VPWR VPWR net7597 sky130_fd_sc_hd__clkbuf_1
Xwire6852 net6850 VGND VGND VPWR VPWR net6852 sky130_fd_sc_hd__clkbuf_2
Xmax_length3284 net3285 VGND VGND VPWR VPWR net3284 sky130_fd_sc_hd__clkbuf_2
Xmax_length3295 _09097_ VGND VGND VPWR VPWR net3295 sky130_fd_sc_hd__buf_1
Xwire6863 net6864 VGND VGND VPWR VPWR net6863 sky130_fd_sc_hd__buf_1
X_14143_ net7626 net1121 VGND VGND VPWR VPWR _06404_ sky130_fd_sc_hd__nand2_1
Xwire6874 net6872 VGND VGND VPWR VPWR net6874 sky130_fd_sc_hd__buf_1
XFILLER_0_21_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6885 net6886 VGND VGND VPWR VPWR net6885 sky130_fd_sc_hd__buf_1
XFILLER_0_132_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6896 net6897 VGND VGND VPWR VPWR net6896 sky130_fd_sc_hd__buf_1
XFILLER_0_158_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14074_ net1332 _06221_ net7604 VGND VGND VPWR VPWR _06337_ sky130_fd_sc_hd__o21a_1
X_18951_ net6166 net6093 VGND VGND VPWR VPWR _10788_ sky130_fd_sc_hd__nand2_1
X_13025_ _05290_ _05297_ VGND VGND VPWR VPWR _05298_ sky130_fd_sc_hd__nor2_1
X_17902_ net2553 _09752_ VGND VGND VPWR VPWR _09753_ sky130_fd_sc_hd__xnor2_1
X_18882_ _10682_ _10683_ net6781 VGND VGND VPWR VPWR _10724_ sky130_fd_sc_hd__o21ai_1
X_17833_ _09600_ _09602_ VGND VGND VPWR VPWR _09684_ sky130_fd_sc_hd__and2b_1
XFILLER_0_174_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17764_ _09614_ VGND VGND VPWR VPWR _09615_ sky130_fd_sc_hd__buf_1
X_14976_ net3544 net3541 net3539 VGND VGND VPWR VPWR _07050_ sky130_fd_sc_hd__a21oi_1
Xwire1170 _01971_ VGND VGND VPWR VPWR net1170 sky130_fd_sc_hd__clkbuf_2
X_19503_ _11332_ _11339_ VGND VGND VPWR VPWR _11340_ sky130_fd_sc_hd__xnor2_1
Xwire1181 _01394_ VGND VGND VPWR VPWR net1181 sky130_fd_sc_hd__buf_1
X_16715_ _08740_ _08736_ _08741_ VGND VGND VPWR VPWR _08742_ sky130_fd_sc_hd__a21o_1
X_13927_ net7743 net1571 VGND VGND VPWR VPWR _06193_ sky130_fd_sc_hd__nand2_1
Xwire1192 _11218_ VGND VGND VPWR VPWR net1192 sky130_fd_sc_hd__buf_1
X_17695_ net2571 _09202_ net1925 VGND VGND VPWR VPWR _00412_ sky130_fd_sc_hd__a21o_1
XFILLER_0_156_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19434_ net6148 VGND VGND VPWR VPWR _11271_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_179_Right_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16646_ matmul0.matmul_stage_inst.mult2\[4\] matmul0.matmul_stage_inst.mult1\[4\]
+ VGND VGND VPWR VPWR _08683_ sky130_fd_sc_hd__xor2_1
X_13858_ _06112_ _06124_ VGND VGND VPWR VPWR _06125_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_88_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12809_ _04979_ _04994_ _04997_ net1611 VGND VGND VPWR VPWR _05082_ sky130_fd_sc_hd__o31a_1
X_19365_ _11196_ _11199_ _11185_ VGND VGND VPWR VPWR _11202_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_108_clk clknet_4_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_108_clk
+ sky130_fd_sc_hd__clkbuf_16
X_16577_ _08635_ VGND VGND VPWR VPWR _00230_ sky130_fd_sc_hd__clkbuf_1
X_13789_ net7653 net1962 _05975_ _05974_ VGND VGND VPWR VPWR _06057_ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18316_ net3241 _09909_ VGND VGND VPWR VPWR _10167_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15528_ net6642 net6593 net7401 VGND VGND VPWR VPWR _07601_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19296_ net6290 net6334 VGND VGND VPWR VPWR _11133_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18247_ net3973 _10097_ VGND VGND VPWR VPWR _10098_ sky130_fd_sc_hd__and2_1
XFILLER_0_167_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15459_ _07381_ _07382_ _07532_ VGND VGND VPWR VPWR _07533_ sky130_fd_sc_hd__o21a_1
XFILLER_0_26_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18178_ _09817_ _10024_ _10028_ VGND VGND VPWR VPWR _10029_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17129_ net1476 _09073_ _09072_ VGND VGND VPWR VPWR _09084_ sky130_fd_sc_hd__or3_1
X_20140_ net274 _11963_ VGND VGND VPWR VPWR _11967_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20071_ net1404 _11898_ _11899_ VGND VGND VPWR VPWR _11900_ sky130_fd_sc_hd__o21a_1
XFILLER_0_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23830_ net4526 net5020 VGND VGND VPWR VPWR _03695_ sky130_fd_sc_hd__nand2_1
X_23761_ _03623_ _03626_ VGND VGND VPWR VPWR _03627_ sky130_fd_sc_hd__xnor2_2
X_20973_ _00987_ _00988_ VGND VGND VPWR VPWR _00989_ sky130_fd_sc_hd__nand2_1
X_25500_ clknet_leaf_41_clk _00380_ net8768 VGND VGND VPWR VPWR svm0.delta\[5\] sky130_fd_sc_hd__dfrtp_1
X_22712_ _02649_ net5391 net3094 VGND VGND VPWR VPWR _02650_ sky130_fd_sc_hd__mux2_1
Xmax_length6816 net6817 VGND VGND VPWR VPWR net6816 sky130_fd_sc_hd__buf_1
X_23692_ _03542_ _03558_ VGND VGND VPWR VPWR _03559_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_146_Right_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25431_ clknet_leaf_94_clk _00314_ net8445 VGND VGND VPWR VPWR matmul0.sin\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_94_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22643_ _01642_ net3076 net2040 _02606_ net8891 VGND VGND VPWR VPWR _00571_ sky130_fd_sc_hd__o311a_1
XFILLER_0_94_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25362_ clknet_leaf_72_clk _00245_ net8472 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult2\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22574_ net7329 _02551_ VGND VGND VPWR VPWR _02555_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24313_ _04171_ _04040_ _04172_ VGND VGND VPWR VPWR _04173_ sky130_fd_sc_hd__o21a_1
XFILLER_0_119_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21525_ _01535_ _01536_ VGND VGND VPWR VPWR _01538_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25293_ clknet_leaf_88_clk _00176_ net8435 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.d\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire6115 net6116 VGND VGND VPWR VPWR net6115 sky130_fd_sc_hd__buf_1
XFILLER_0_17_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24244_ _04048_ net589 VGND VGND VPWR VPWR _04105_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6126 net6122 VGND VGND VPWR VPWR net6126 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21456_ _01467_ _01468_ VGND VGND VPWR VPWR _01469_ sky130_fd_sc_hd__xnor2_1
Xwire6137 net6132 VGND VGND VPWR VPWR net6137 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire5403 net5405 VGND VGND VPWR VPWR net5403 sky130_fd_sc_hd__clkbuf_1
Xwire6148 net6149 VGND VGND VPWR VPWR net6148 sky130_fd_sc_hd__buf_1
Xwire5414 net5415 VGND VGND VPWR VPWR net5414 sky130_fd_sc_hd__clkbuf_1
Xwire5425 net5426 VGND VGND VPWR VPWR net5425 sky130_fd_sc_hd__buf_1
X_20407_ _09082_ _12203_ VGND VGND VPWR VPWR _12204_ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24175_ pid_q.curr_int\[8\] net3757 _02870_ _04036_ VGND VGND VPWR VPWR _00673_ sky130_fd_sc_hd__a22o_1
Xwire4702 net4703 VGND VGND VPWR VPWR net4702 sky130_fd_sc_hd__buf_1
Xwire5447 net5448 VGND VGND VPWR VPWR net5447 sky130_fd_sc_hd__clkbuf_1
X_21387_ _01265_ _01266_ _01264_ VGND VGND VPWR VPWR _01401_ sky130_fd_sc_hd__o21ba_1
Xwire5458 net5453 VGND VGND VPWR VPWR net5458 sky130_fd_sc_hd__buf_1
Xwire5469 net5470 VGND VGND VPWR VPWR net5469 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23126_ net5130 net4657 VGND VGND VPWR VPWR _02996_ sky130_fd_sc_hd__nand2_1
Xwire4735 net4736 VGND VGND VPWR VPWR net4735 sky130_fd_sc_hd__clkbuf_1
Xwire4746 net4747 VGND VGND VPWR VPWR net4746 sky130_fd_sc_hd__clkbuf_1
X_20338_ _12139_ _12140_ VGND VGND VPWR VPWR _12141_ sky130_fd_sc_hd__and2b_1
Xwire4757 net4758 VGND VGND VPWR VPWR net4757 sky130_fd_sc_hd__buf_1
Xwire4768 net4769 VGND VGND VPWR VPWR net4768 sky130_fd_sc_hd__buf_1
X_23057_ _02925_ net4865 net4772 _02926_ VGND VGND VPWR VPWR _02927_ sky130_fd_sc_hd__a31o_1
X_20269_ net3 net4 _12072_ net8121 VGND VGND VPWR VPWR _12079_ sky130_fd_sc_hd__a31o_1
Xinput101 pid_d_data[13] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_1
Xinput112 pid_d_data[9] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22008_ net9035 net3123 net2078 _02015_ VGND VGND VPWR VPWR _00527_ sky130_fd_sc_hd__a22o_1
Xinput123 pid_q_addr[3] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_1
Xinput134 pid_q_data[13] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_1
Xinput145 pid_q_data[9] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_1
X_14830_ net9231 matmul0.matmul_stage_inst.e\[4\] net3610 VGND VGND VPWR VPWR _06932_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length8752 net8753 VGND VGND VPWR VPWR net8752 sky130_fd_sc_hd__buf_1
XFILLER_0_53_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14761_ net7152 _06890_ VGND VGND VPWR VPWR _06891_ sky130_fd_sc_hd__xor2_1
X_23959_ _03817_ _03822_ VGND VGND VPWR VPWR _03823_ sky130_fd_sc_hd__xor2_1
X_16500_ net2772 net2783 VGND VGND VPWR VPWR _08560_ sky130_fd_sc_hd__nand2_1
X_13712_ _05911_ _05912_ VGND VGND VPWR VPWR _05981_ sky130_fd_sc_hd__or2_1
X_17480_ _09295_ _09367_ net6718 VGND VGND VPWR VPWR _09371_ sky130_fd_sc_hd__o21ba_1
X_14692_ matmul0.sin\[4\] net7155 _06832_ VGND VGND VPWR VPWR _06839_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_113_Right_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16431_ _08480_ _08481_ net303 VGND VGND VPWR VPWR _08492_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_195_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13643_ _05911_ _05912_ VGND VGND VPWR VPWR _05913_ sky130_fd_sc_hd__xnor2_1
X_25629_ clknet_leaf_108_clk _00502_ net8350 VGND VGND VPWR VPWR cordic0.vec\[0\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_27_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19150_ net6355 _10986_ VGND VGND VPWR VPWR _10987_ sky130_fd_sc_hd__xnor2_1
X_13574_ _05842_ net783 VGND VGND VPWR VPWR _05845_ sky130_fd_sc_hd__xnor2_2
X_16362_ _08311_ net1083 net1509 VGND VGND VPWR VPWR _08425_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18101_ _09872_ _09873_ VGND VGND VPWR VPWR _09952_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8051 net8052 VGND VGND VPWR VPWR net8051 sky130_fd_sc_hd__clkbuf_1
X_15313_ net1872 _07386_ VGND VGND VPWR VPWR _07387_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_147_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19081_ net6247 net6321 VGND VGND VPWR VPWR _10918_ sky130_fd_sc_hd__nand2_1
Xfanout6521 net6526 VGND VGND VPWR VPWR net6521 sky130_fd_sc_hd__clkbuf_2
Xwire8062 net8063 VGND VGND VPWR VPWR net8062 sky130_fd_sc_hd__buf_1
X_16293_ _08353_ net724 VGND VGND VPWR VPWR _08357_ sky130_fd_sc_hd__nand2_1
Xwire8084 net8085 VGND VGND VPWR VPWR net8084 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8095 net98 VGND VGND VPWR VPWR net8095 sky130_fd_sc_hd__clkbuf_1
X_18032_ _09868_ _09882_ VGND VGND VPWR VPWR _09883_ sky130_fd_sc_hd__xnor2_2
Xwire7350 net7351 VGND VGND VPWR VPWR net7350 sky130_fd_sc_hd__clkbuf_1
X_15244_ _07316_ _07317_ VGND VGND VPWR VPWR _07318_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_83_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7372 net7373 VGND VGND VPWR VPWR net7372 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7394 net7395 VGND VGND VPWR VPWR net7394 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15175_ net2849 net2730 net3446 _07246_ _07248_ VGND VGND VPWR VPWR _07249_ sky130_fd_sc_hd__a32o_1
XFILLER_0_105_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6682 net149 VGND VGND VPWR VPWR net6682 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14126_ net1332 _06221_ _06235_ VGND VGND VPWR VPWR _06388_ sky130_fd_sc_hd__and3_1
Xwire5970 pid_d.curr_error\[3\] VGND VGND VPWR VPWR net5970 sky130_fd_sc_hd__buf_1
XFILLER_0_162_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19983_ _11768_ net1408 _11813_ VGND VGND VPWR VPWR _11814_ sky130_fd_sc_hd__a21o_1
Xwire5981 pid_d.curr_int\[4\] VGND VGND VPWR VPWR net5981 sky130_fd_sc_hd__clkbuf_2
X_14057_ _06277_ _06320_ VGND VGND VPWR VPWR _06321_ sky130_fd_sc_hd__xnor2_1
X_18934_ net3982 _10751_ net3224 VGND VGND VPWR VPWR _10773_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13008_ net1336 _05100_ VGND VGND VPWR VPWR _05281_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18865_ net6770 _10677_ net2589 VGND VGND VPWR VPWR _10707_ sky130_fd_sc_hd__o21a_1
XFILLER_0_158_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17816_ net3259 net2563 VGND VGND VPWR VPWR _09667_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_19_Left_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18796_ _10637_ _10639_ VGND VGND VPWR VPWR _10640_ sky130_fd_sc_hd__xnor2_1
X_17747_ net1786 VGND VGND VPWR VPWR _09598_ sky130_fd_sc_hd__buf_1
XFILLER_0_178_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14959_ _07017_ _07032_ VGND VGND VPWR VPWR _07033_ sky130_fd_sc_hd__xnor2_1
X_17678_ svm0.tA\[7\] _09539_ svm0.counter\[7\] VGND VGND VPWR VPWR _09558_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_187_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19417_ _11009_ _10994_ _11253_ VGND VGND VPWR VPWR _11254_ sky130_fd_sc_hd__a21o_1
X_16629_ matmul0.matmul_stage_inst.mult2\[2\] matmul0.matmul_stage_inst.mult1\[2\]
+ VGND VGND VPWR VPWR _08668_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19348_ _11168_ _11184_ VGND VGND VPWR VPWR _11185_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19279_ _11109_ _11110_ net872 VGND VGND VPWR VPWR _11116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_28_Left_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21310_ _01315_ _01324_ VGND VGND VPWR VPWR _01325_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_170_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22290_ _02292_ _02293_ VGND VGND VPWR VPWR _02294_ sky130_fd_sc_hd__xor2_1
XFILLER_0_14_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21241_ _00838_ net1393 _01255_ VGND VGND VPWR VPWR _01256_ sky130_fd_sc_hd__a21o_1
Xwire4009 net4010 VGND VGND VPWR VPWR net4009 sky130_fd_sc_hd__buf_1
XFILLER_0_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21172_ net2073 _01156_ VGND VGND VPWR VPWR _01188_ sky130_fd_sc_hd__xor2_2
XFILLER_0_159_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3319 _09023_ VGND VGND VPWR VPWR net3319 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20123_ _11949_ _11950_ VGND VGND VPWR VPWR _11951_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2607 net2610 VGND VGND VPWR VPWR net2607 sky130_fd_sc_hd__buf_1
XFILLER_0_102_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2618 _08636_ VGND VGND VPWR VPWR net2618 sky130_fd_sc_hd__buf_1
Xwire2629 _07933_ VGND VGND VPWR VPWR net2629 sky130_fd_sc_hd__buf_1
X_24931_ pid_q.ki\[6\] _04714_ net1361 VGND VGND VPWR VPWR _04715_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_37_Left_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20054_ net3855 _11861_ _11879_ net6077 _11882_ VGND VGND VPWR VPWR _11883_ sky130_fd_sc_hd__a221o_1
Xwire1906 net1907 VGND VGND VPWR VPWR net1906 sky130_fd_sc_hd__clkbuf_1
Xwire1917 net1918 VGND VGND VPWR VPWR net1917 sky130_fd_sc_hd__buf_1
Xwire1928 net1929 VGND VGND VPWR VPWR net1928 sky130_fd_sc_hd__buf_1
Xwire1939 net1941 VGND VGND VPWR VPWR net1939 sky130_fd_sc_hd__buf_1
X_24862_ net1999 net4744 net2002 VGND VGND VPWR VPWR _04666_ sky130_fd_sc_hd__mux2_1
X_23813_ _03656_ _03676_ _03677_ VGND VGND VPWR VPWR _03678_ sky130_fd_sc_hd__a21o_1
X_24793_ net5198 VGND VGND VPWR VPWR _04618_ sky130_fd_sc_hd__inv_2
X_23744_ net2412 _03609_ VGND VGND VPWR VPWR _03610_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20956_ net5759 net5792 _00971_ VGND VGND VPWR VPWR _00972_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_184_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6624 net6625 VGND VGND VPWR VPWR net6624 sky130_fd_sc_hd__clkbuf_1
Xmax_length6635 net6636 VGND VGND VPWR VPWR net6635 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_177_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23675_ _03509_ _03541_ VGND VGND VPWR VPWR _03542_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_166_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20887_ net5601 net5821 VGND VGND VPWR VPWR _00903_ sky130_fd_sc_hd__nand2_1
X_22626_ pid_d.curr_error\[14\] net800 _02561_ VGND VGND VPWR VPWR _02596_ sky130_fd_sc_hd__mux2_1
X_25414_ clknet_leaf_86_clk _00297_ net8531 VGND VGND VPWR VPWR matmul0.cos\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_181_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_46_Left_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25345_ clknet_leaf_72_clk _00228_ net8472 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_22557_ net4390 net4380 net4315 net4327 VGND VGND VPWR VPWR _02541_ sky130_fd_sc_hd__nor4_1
XFILLER_0_9_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21508_ _01442_ _01520_ VGND VGND VPWR VPWR _01521_ sky130_fd_sc_hd__xnor2_1
X_13290_ _05553_ _05562_ VGND VGND VPWR VPWR _05563_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25276_ clknet_leaf_77_clk _00159_ net8457 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.c\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout5127 pid_q.mult0.b\[1\] VGND VGND VPWR VPWR net5127 sky130_fd_sc_hd__clkbuf_1
X_22488_ net5407 _02487_ _02488_ VGND VGND VPWR VPWR _02489_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5200 net5201 VGND VGND VPWR VPWR net5200 sky130_fd_sc_hd__buf_1
X_24227_ _04074_ _04087_ VGND VGND VPWR VPWR _04088_ sky130_fd_sc_hd__xnor2_1
Xwire5211 net5212 VGND VGND VPWR VPWR net5211 sky130_fd_sc_hd__clkbuf_1
X_21439_ _01448_ _01451_ VGND VGND VPWR VPWR _01452_ sky130_fd_sc_hd__xnor2_1
Xwire5233 net5234 VGND VGND VPWR VPWR net5233 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5244 net5245 VGND VGND VPWR VPWR net5244 sky130_fd_sc_hd__clkbuf_1
Xwire4510 net4511 VGND VGND VPWR VPWR net4510 sky130_fd_sc_hd__clkbuf_1
Xwire5255 net5256 VGND VGND VPWR VPWR net5255 sky130_fd_sc_hd__buf_1
X_24158_ net1160 _03927_ _04019_ VGND VGND VPWR VPWR _04020_ sky130_fd_sc_hd__a21oi_1
Xwire4521 net4522 VGND VGND VPWR VPWR net4521 sky130_fd_sc_hd__buf_1
Xwire5266 net5267 VGND VGND VPWR VPWR net5266 sky130_fd_sc_hd__clkbuf_1
Xwire4532 net4525 VGND VGND VPWR VPWR net4532 sky130_fd_sc_hd__buf_1
XFILLER_0_48_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4543 net4548 VGND VGND VPWR VPWR net4543 sky130_fd_sc_hd__buf_1
Xwire5288 net5289 VGND VGND VPWR VPWR net5288 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4554 net4555 VGND VGND VPWR VPWR net4554 sky130_fd_sc_hd__buf_1
Xwire5299 net5300 VGND VGND VPWR VPWR net5299 sky130_fd_sc_hd__buf_1
X_23109_ net5000 net4718 VGND VGND VPWR VPWR _02979_ sky130_fd_sc_hd__nand2_1
Xwire4565 net4566 VGND VGND VPWR VPWR net4565 sky130_fd_sc_hd__buf_1
Xwire3820 net3821 VGND VGND VPWR VPWR net3820 sky130_fd_sc_hd__clkbuf_1
Xwire3831 net3832 VGND VGND VPWR VPWR net3831 sky130_fd_sc_hd__clkbuf_1
Xwire4576 net4570 VGND VGND VPWR VPWR net4576 sky130_fd_sc_hd__buf_1
X_24089_ net7505 _03950_ _03951_ VGND VGND VPWR VPWR _03952_ sky130_fd_sc_hd__and3_1
X_16980_ net3349 net1232 net878 _08942_ VGND VGND VPWR VPWR _00326_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_55_Left_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4587 pid_q.mult0.a\[10\] VGND VGND VPWR VPWR net4587 sky130_fd_sc_hd__clkbuf_1
Xwire3842 _00851_ VGND VGND VPWR VPWR net3842 sky130_fd_sc_hd__buf_1
Xwire4598 net4599 VGND VGND VPWR VPWR net4598 sky130_fd_sc_hd__buf_1
Xwire3853 _12265_ VGND VGND VPWR VPWR net3853 sky130_fd_sc_hd__buf_1
Xwire3864 net3865 VGND VGND VPWR VPWR net3864 sky130_fd_sc_hd__buf_1
Xwire3875 _11054_ VGND VGND VPWR VPWR net3875 sky130_fd_sc_hd__clkbuf_1
X_15931_ _07894_ net1263 _07895_ VGND VGND VPWR VPWR _08000_ sky130_fd_sc_hd__o21a_1
Xwire3886 net3887 VGND VGND VPWR VPWR net3886 sky130_fd_sc_hd__buf_1
Xwire3897 _10839_ VGND VGND VPWR VPWR net3897 sky130_fd_sc_hd__buf_1
X_18650_ _10446_ _10496_ VGND VGND VPWR VPWR _10497_ sky130_fd_sc_hd__and2_1
X_15862_ net2727 _07928_ _07930_ net2234 VGND VGND VPWR VPWR _07931_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17601_ net4009 svm0.tB\[4\] svm0.tB\[3\] net4018 _09481_ VGND VGND VPWR VPWR _09482_
+ sky130_fd_sc_hd__o221a_1
X_14813_ net8978 net2871 _06923_ VGND VGND VPWR VPWR _00178_ sky130_fd_sc_hd__a21o_1
XFILLER_0_189_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18581_ net7016 net6952 VGND VGND VPWR VPWR _10429_ sky130_fd_sc_hd__or2_1
X_15793_ net2836 net2658 VGND VGND VPWR VPWR _07863_ sky130_fd_sc_hd__nor2_1
X_17532_ net6686 svm0.delta\[14\] net6742 net6694 VGND VGND VPWR VPWR _09415_ sky130_fd_sc_hd__o211a_1
Xmax_length8571 net8572 VGND VGND VPWR VPWR net8571 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14744_ net9063 net2860 net2259 _06877_ VGND VGND VPWR VPWR _00155_ sky130_fd_sc_hd__a22o_1
XFILLER_0_171_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17463_ svm0.counter\[4\] net2577 VGND VGND VPWR VPWR _09357_ sky130_fd_sc_hd__nor2_1
XFILLER_0_188_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_64_Left_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14675_ net7454 VGND VGND VPWR VPWR _06826_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19202_ net3180 _11038_ VGND VGND VPWR VPWR _11039_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16414_ _08440_ _08475_ VGND VGND VPWR VPWR _08476_ sky130_fd_sc_hd__xnor2_1
X_13626_ net7675 net2322 net2318 VGND VGND VPWR VPWR _05896_ sky130_fd_sc_hd__and3_1
X_17394_ net2572 _09300_ VGND VGND VPWR VPWR _09301_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout7030 net7037 VGND VGND VPWR VPWR net7030 sky130_fd_sc_hd__buf_1
X_19133_ _10862_ _10966_ _10969_ VGND VGND VPWR VPWR _10970_ sky130_fd_sc_hd__a21o_1
X_16345_ net882 _08407_ VGND VGND VPWR VPWR _08408_ sky130_fd_sc_hd__xnor2_2
X_13557_ _05824_ _05827_ VGND VGND VPWR VPWR _05828_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6351 net6354 VGND VGND VPWR VPWR net6351 sky130_fd_sc_hd__clkbuf_1
X_19064_ _10898_ net2525 VGND VGND VPWR VPWR _10901_ sky130_fd_sc_hd__and2_1
X_13488_ _05698_ net622 VGND VGND VPWR VPWR _05761_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout7096 net7100 VGND VGND VPWR VPWR net7096 sky130_fd_sc_hd__clkbuf_2
X_16276_ net1087 net981 VGND VGND VPWR VPWR _08340_ sky130_fd_sc_hd__and2b_1
XFILLER_0_81_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18015_ _09860_ net2550 VGND VGND VPWR VPWR _09866_ sky130_fd_sc_hd__nand2_1
Xfanout5650 pid_d.mult0.b\[15\] VGND VGND VPWR VPWR net5650 sky130_fd_sc_hd__clkbuf_1
X_15227_ net1276 _07300_ VGND VGND VPWR VPWR _07301_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6490 net6488 VGND VGND VPWR VPWR net6490 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15158_ net3568 net2742 _07229_ net2242 VGND VGND VPWR VPWR _07232_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_73_Left_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14109_ _06325_ _06329_ _06370_ VGND VGND VPWR VPWR _06371_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19966_ net4046 _11572_ VGND VGND VPWR VPWR _11797_ sky130_fd_sc_hd__xnor2_2
X_15089_ _07094_ net1895 _07162_ VGND VGND VPWR VPWR _07163_ sky130_fd_sc_hd__a21o_1
X_18917_ net6876 net6801 VGND VGND VPWR VPWR _10757_ sky130_fd_sc_hd__nand2_1
X_19897_ cordic0.cos\[4\] net2942 net1782 VGND VGND VPWR VPWR _11730_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18848_ net6781 _10687_ _10688_ _10690_ VGND VGND VPWR VPWR _10691_ sky130_fd_sc_hd__a31o_1
XFILLER_0_179_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18779_ _10407_ _10515_ _10622_ VGND VGND VPWR VPWR _10623_ sky130_fd_sc_hd__or3_1
XFILLER_0_179_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20810_ net5861 net5494 VGND VGND VPWR VPWR _00826_ sky130_fd_sc_hd__nand2_2
XFILLER_0_145_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21790_ _01795_ _01799_ VGND VGND VPWR VPWR _01800_ sky130_fd_sc_hd__xor2_1
XFILLER_0_166_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20741_ _12509_ _12510_ _12511_ VGND VGND VPWR VPWR _12512_ sky130_fd_sc_hd__o21a_1
XFILLER_0_175_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8809 net8810 VGND VGND VPWR VPWR net8809 sky130_fd_sc_hd__buf_1
X_23460_ net5162 net4513 VGND VGND VPWR VPWR _03329_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20672_ net6091 net1473 VGND VGND VPWR VPWR _12449_ sky130_fd_sc_hd__nand2_1
XFILLER_0_190_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22411_ _02382_ _02412_ VGND VGND VPWR VPWR _02413_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23391_ _03259_ _03260_ VGND VGND VPWR VPWR _03261_ sky130_fd_sc_hd__or2b_1
Xclkbuf_leaf_30_clk clknet_4_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_6_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25130_ clknet_leaf_52_clk _00019_ net8805 VGND VGND VPWR VPWR svm0.tC\[2\] sky130_fd_sc_hd__dfrtp_1
X_22342_ net944 _02344_ VGND VGND VPWR VPWR _02345_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_72_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25061_ net266 net1630 _04808_ net4430 _04809_ VGND VGND VPWR VPWR _00786_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22273_ _02248_ _02276_ _02249_ VGND VGND VPWR VPWR _02277_ sky130_fd_sc_hd__a21oi_1
X_24012_ net5067 _03873_ _03874_ VGND VGND VPWR VPWR _03875_ sky130_fd_sc_hd__a21o_1
XFILLER_0_130_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold130 pid_d.prev_error\[15\] VGND VGND VPWR VPWR net9083 sky130_fd_sc_hd__dlygate4sd3_1
X_21224_ _01221_ _01235_ _01238_ _01239_ VGND VGND VPWR VPWR _01240_ sky130_fd_sc_hd__a211o_1
Xhold141 matmul0.matmul_stage_inst.b\[7\] VGND VGND VPWR VPWR net9094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 pid_d.prev_error\[9\] VGND VGND VPWR VPWR net9105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 matmul0.matmul_stage_inst.c\[12\] VGND VGND VPWR VPWR net9116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 pid_q.prev_error\[10\] VGND VGND VPWR VPWR net9127 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3116 net3117 VGND VGND VPWR VPWR net3116 sky130_fd_sc_hd__buf_1
X_21155_ _01169_ _01170_ VGND VGND VPWR VPWR _01171_ sky130_fd_sc_hd__xor2_1
Xwire3127 _11620_ VGND VGND VPWR VPWR net3127 sky130_fd_sc_hd__buf_1
Xhold185 pid_d.prev_error\[4\] VGND VGND VPWR VPWR net9138 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3138 _11431_ VGND VGND VPWR VPWR net3138 sky130_fd_sc_hd__buf_1
Xhold196 svm0.tC\[2\] VGND VGND VPWR VPWR net9149 sky130_fd_sc_hd__dlygate4sd3_1
Xwire2404 _04224_ VGND VGND VPWR VPWR net2404 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2415 net2416 VGND VGND VPWR VPWR net2415 sky130_fd_sc_hd__clkbuf_1
X_20106_ _11906_ _11904_ _11933_ VGND VGND VPWR VPWR _11934_ sky130_fd_sc_hd__o21a_2
Xwire2426 _03333_ VGND VGND VPWR VPWR net2426 sky130_fd_sc_hd__buf_1
XFILLER_0_176_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2437 net2438 VGND VGND VPWR VPWR net2437 sky130_fd_sc_hd__clkbuf_1
X_21086_ _01101_ _01062_ net1731 VGND VGND VPWR VPWR _01102_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_186_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1703 _02231_ VGND VGND VPWR VPWR net1703 sky130_fd_sc_hd__buf_1
Xwire2448 net2449 VGND VGND VPWR VPWR net2448 sky130_fd_sc_hd__buf_2
XFILLER_0_95_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1714 _01939_ VGND VGND VPWR VPWR net1714 sky130_fd_sc_hd__buf_1
Xwire2459 _02543_ VGND VGND VPWR VPWR net2459 sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_97_clk clknet_4_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_97_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_77_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1725 _01497_ VGND VGND VPWR VPWR net1725 sky130_fd_sc_hd__buf_1
X_24914_ _04703_ VGND VGND VPWR VPWR _00745_ sky130_fd_sc_hd__clkbuf_1
X_20037_ _11863_ _11866_ VGND VGND VPWR VPWR _11867_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1736 _00836_ VGND VGND VPWR VPWR net1736 sky130_fd_sc_hd__buf_1
X_25894_ clknet_leaf_14_clk _00767_ net8621 VGND VGND VPWR VPWR pid_q.kp\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_176_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1747 net1748 VGND VGND VPWR VPWR net1747 sky130_fd_sc_hd__buf_1
Xwire1758 _10902_ VGND VGND VPWR VPWR net1758 sky130_fd_sc_hd__buf_1
Xwire1769 _10264_ VGND VGND VPWR VPWR net1769 sky130_fd_sc_hd__clkbuf_1
X_24845_ net4874 net2007 _04540_ net327 VGND VGND VPWR VPWR _00724_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length7111 net7112 VGND VGND VPWR VPWR net7111 sky130_fd_sc_hd__buf_1
X_12790_ net7875 _04962_ net2971 VGND VGND VPWR VPWR _05063_ sky130_fd_sc_hd__and3_1
X_24776_ net7479 _04535_ net457 net9193 _04529_ VGND VGND VPWR VPWR _00707_ sky130_fd_sc_hd__a32o_1
X_21988_ _01989_ _01995_ VGND VGND VPWR VPWR _01996_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23727_ _03589_ _03592_ VGND VGND VPWR VPWR _03593_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20939_ _00949_ _00951_ _00954_ VGND VGND VPWR VPWR _00955_ sky130_fd_sc_hd__a21o_1
XFILLER_0_166_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length6476 net6477 VGND VGND VPWR VPWR net6476 sky130_fd_sc_hd__clkbuf_1
X_14460_ net6443 _06541_ VGND VGND VPWR VPWR _06649_ sky130_fd_sc_hd__nor2_1
X_23658_ _03397_ _03406_ _03405_ VGND VGND VPWR VPWR _03525_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_165_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13411_ net731 _05633_ _05573_ VGND VGND VPWR VPWR _05684_ sky130_fd_sc_hd__a21o_1
Xmax_length5775 net5776 VGND VGND VPWR VPWR net5775 sky130_fd_sc_hd__buf_1
XFILLER_0_187_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22609_ net8888 _02582_ VGND VGND VPWR VPWR _02583_ sky130_fd_sc_hd__and2_1
X_14391_ _06596_ VGND VGND VPWR VPWR _00083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23589_ net4784 net3746 VGND VGND VPWR VPWR _03457_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13342_ _05343_ _05344_ _05052_ VGND VGND VPWR VPWR _05615_ sky130_fd_sc_hd__o21a_1
X_16130_ _08194_ _08195_ net2645 net2659 VGND VGND VPWR VPWR _08196_ sky130_fd_sc_hd__a211o_1
X_25328_ clknet_leaf_80_clk _00211_ net8497 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.f\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13273_ _05544_ _05541_ _05542_ VGND VGND VPWR VPWR _05546_ sky130_fd_sc_hd__and3_1
X_16061_ _08025_ _08030_ _08023_ VGND VGND VPWR VPWR _08128_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25259_ clknet_leaf_71_clk _00142_ net8457 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.b\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire5030 net5021 VGND VGND VPWR VPWR net5030 sky130_fd_sc_hd__buf_1
Xwire5041 net5042 VGND VGND VPWR VPWR net5041 sky130_fd_sc_hd__clkbuf_1
X_15012_ net4126 net4124 VGND VGND VPWR VPWR _07086_ sky130_fd_sc_hd__or2_1
Xwire5052 net5053 VGND VGND VPWR VPWR net5052 sky130_fd_sc_hd__buf_1
Xwire5063 net5064 VGND VGND VPWR VPWR net5063 sky130_fd_sc_hd__buf_1
Xwire5074 net5075 VGND VGND VPWR VPWR net5074 sky130_fd_sc_hd__buf_1
Xwire5085 net5088 VGND VGND VPWR VPWR net5085 sky130_fd_sc_hd__clkbuf_1
Xwire4340 pid_d.state\[4\] VGND VGND VPWR VPWR net4340 sky130_fd_sc_hd__clkbuf_1
X_19820_ _11631_ _11653_ VGND VGND VPWR VPWR _11654_ sky130_fd_sc_hd__xor2_2
Xwire5096 net5097 VGND VGND VPWR VPWR net5096 sky130_fd_sc_hd__buf_1
Xwire4351 pid_d.state\[3\] VGND VGND VPWR VPWR net4351 sky130_fd_sc_hd__buf_1
Xwire4362 net4363 VGND VGND VPWR VPWR net4362 sky130_fd_sc_hd__buf_1
Xwire4373 net4374 VGND VGND VPWR VPWR net4373 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4384 net4385 VGND VGND VPWR VPWR net4384 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3650 net3651 VGND VGND VPWR VPWR net3650 sky130_fd_sc_hd__clkbuf_1
Xwire4395 net4396 VGND VGND VPWR VPWR net4395 sky130_fd_sc_hd__clkbuf_1
X_19751_ net6097 _11329_ _11383_ _11585_ VGND VGND VPWR VPWR _11586_ sky130_fd_sc_hd__a211oi_2
Xwire3661 net3662 VGND VGND VPWR VPWR net3661 sky130_fd_sc_hd__clkbuf_1
X_16963_ net6055 net5996 net6501 VGND VGND VPWR VPWR _08926_ sky130_fd_sc_hd__mux2_1
Xwire3672 net3673 VGND VGND VPWR VPWR net3672 sky130_fd_sc_hd__clkbuf_1
Xwire3683 _05531_ VGND VGND VPWR VPWR net3683 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_88_clk clknet_4_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_88_clk sky130_fd_sc_hd__clkbuf_16
Xwire3694 _04897_ VGND VGND VPWR VPWR net3694 sky130_fd_sc_hd__buf_1
XFILLER_0_21_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18702_ net6779 net2126 _10547_ VGND VGND VPWR VPWR _10548_ sky130_fd_sc_hd__mux2_1
Xwire2960 net2961 VGND VGND VPWR VPWR net2960 sky130_fd_sc_hd__buf_1
X_15914_ _07977_ _07982_ VGND VGND VPWR VPWR _07983_ sky130_fd_sc_hd__xnor2_1
X_19682_ net6199 net6275 VGND VGND VPWR VPWR _11518_ sky130_fd_sc_hd__or2_1
XFILLER_0_194_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16894_ net6399 _08857_ VGND VGND VPWR VPWR _08858_ sky130_fd_sc_hd__nor2_1
Xwire2993 net2994 VGND VGND VPWR VPWR net2993 sky130_fd_sc_hd__buf_1
X_18633_ _10478_ net3938 net6878 _10479_ VGND VGND VPWR VPWR _10480_ sky130_fd_sc_hd__o2bb2a_1
X_15845_ _07821_ VGND VGND VPWR VPWR _07915_ sky130_fd_sc_hd__inv_2
XFILLER_0_182_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18564_ _10331_ net765 _10410_ _10396_ VGND VGND VPWR VPWR _10412_ sky130_fd_sc_hd__a31o_1
X_15776_ net3550 net3600 VGND VGND VPWR VPWR _07846_ sky130_fd_sc_hd__nor2_1
X_12988_ _05255_ _05260_ VGND VGND VPWR VPWR _05261_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17515_ svm0.delta\[12\] _09400_ VGND VGND VPWR VPWR _09401_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14727_ net8973 _06820_ net890 VGND VGND VPWR VPWR _00151_ sky130_fd_sc_hd__a21bo_1
X_18495_ net1784 VGND VGND VPWR VPWR _10344_ sky130_fd_sc_hd__buf_1
XFILLER_0_157_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17446_ net6738 net6744 VGND VGND VPWR VPWR _09342_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14658_ net8956 net2880 _06813_ VGND VGND VPWR VPWR _00133_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13609_ net7792 net1306 _05786_ _05787_ VGND VGND VPWR VPWR _05879_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_89_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17377_ svm0.delta\[4\] VGND VGND VPWR VPWR _09287_ sky130_fd_sc_hd__inv_2
XFILLER_0_184_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14589_ net2882 net281 _06763_ VGND VGND VPWR VPWR _06764_ sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_12_clk clknet_4_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_16
X_19116_ _10876_ _10899_ VGND VGND VPWR VPWR _10953_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_171_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16328_ _08387_ _08390_ VGND VGND VPWR VPWR _08391_ sky130_fd_sc_hd__xor2_1
XFILLER_0_131_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19047_ _10877_ _10883_ VGND VGND VPWR VPWR _10884_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16259_ _08319_ _08322_ VGND VGND VPWR VPWR _08323_ sky130_fd_sc_hd__xor2_2
XFILLER_0_3_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19949_ _11674_ _11710_ _11708_ VGND VGND VPWR VPWR _11781_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_96_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_79_clk clknet_4_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_79_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22960_ net4370 net201 _02847_ net4331 net2467 VGND VGND VPWR VPWR _02848_ sky130_fd_sc_hd__a221o_1
XFILLER_0_156_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21911_ _01916_ _01821_ _01918_ VGND VGND VPWR VPWR _01919_ sky130_fd_sc_hd__a21o_1
XFILLER_0_179_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22891_ net5354 net3103 VGND VGND VPWR VPWR _02785_ sky130_fd_sc_hd__nor2_1
X_24630_ _04481_ _04484_ _03705_ VGND VGND VPWR VPWR _04485_ sky130_fd_sc_hd__a21o_1
X_21842_ _01756_ _01758_ _01757_ VGND VGND VPWR VPWR _01851_ sky130_fd_sc_hd__o21a_1
XFILLER_0_136_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24561_ net4523 net4825 net4809 _04416_ VGND VGND VPWR VPWR _04417_ sky130_fd_sc_hd__a31o_1
XFILLER_0_136_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21773_ net5839 net5394 VGND VGND VPWR VPWR _01783_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23512_ net1166 net938 _03380_ VGND VGND VPWR VPWR _03381_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20724_ _12483_ _12492_ _12494_ VGND VGND VPWR VPWR _12496_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8606 net8607 VGND VGND VPWR VPWR net8606 sky130_fd_sc_hd__clkbuf_1
X_24492_ _04291_ net3037 VGND VGND VPWR VPWR _04349_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8628 net8627 VGND VGND VPWR VPWR net8628 sky130_fd_sc_hd__buf_1
Xwire8639 net8640 VGND VGND VPWR VPWR net8639 sky130_fd_sc_hd__buf_1
Xmax_length4326 net4327 VGND VGND VPWR VPWR net4326 sky130_fd_sc_hd__buf_1
XFILLER_0_162_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23443_ net3999 _03312_ VGND VGND VPWR VPWR _03313_ sky130_fd_sc_hd__nor2_1
X_20655_ net6132 _12421_ VGND VGND VPWR VPWR _12433_ sky130_fd_sc_hd__nor2_1
Xmax_length3603 _06964_ VGND VGND VPWR VPWR net3603 sky130_fd_sc_hd__buf_1
XFILLER_0_190_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire307 net308 VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__clkbuf_1
Xwire7927 net7928 VGND VGND VPWR VPWR net7927 sky130_fd_sc_hd__clkbuf_1
Xwire318 _06757_ VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7938 net7941 VGND VGND VPWR VPWR net7938 sky130_fd_sc_hd__clkbuf_1
Xwire329 net330 VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__buf_1
Xwire7949 net7950 VGND VGND VPWR VPWR net7949 sky130_fd_sc_hd__buf_1
XFILLER_0_61_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23374_ _03242_ _03243_ VGND VGND VPWR VPWR _03244_ sky130_fd_sc_hd__xnor2_1
X_20586_ _12366_ _12368_ VGND VGND VPWR VPWR _12369_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_33_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22325_ net4363 _02268_ _02274_ net4380 _02328_ VGND VGND VPWR VPWR _02329_ sky130_fd_sc_hd__a221o_1
Xmax_length2935 _06506_ VGND VGND VPWR VPWR net2935 sky130_fd_sc_hd__clkbuf_1
X_25113_ pid_d.prev_int\[1\] net2392 net1992 net5985 VGND VGND VPWR VPWR _00794_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25044_ net3738 _04790_ _04794_ VGND VGND VPWR VPWR _04795_ sky130_fd_sc_hd__a21o_1
X_22256_ net4381 _02187_ net299 net4317 net337 VGND VGND VPWR VPWR _02261_ sky130_fd_sc_hd__a221o_1
XFILLER_0_103_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21207_ net1732 VGND VGND VPWR VPWR _01223_ sky130_fd_sc_hd__inv_2
X_22187_ _02160_ _02189_ _02190_ _02191_ VGND VGND VPWR VPWR _02192_ sky130_fd_sc_hd__a22o_1
XFILLER_0_178_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21138_ net5634 net5872 VGND VGND VPWR VPWR _01154_ sky130_fd_sc_hd__nand2_1
Xwire2212 _07990_ VGND VGND VPWR VPWR net2212 sky130_fd_sc_hd__buf_1
Xwire2234 net2235 VGND VGND VPWR VPWR net2234 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1500 net1501 VGND VGND VPWR VPWR net1500 sky130_fd_sc_hd__buf_1
Xwire2245 net2246 VGND VGND VPWR VPWR net2245 sky130_fd_sc_hd__clkbuf_2
Xwire2256 net2257 VGND VGND VPWR VPWR net2256 sky130_fd_sc_hd__clkbuf_2
Xwire1511 _08220_ VGND VGND VPWR VPWR net1511 sky130_fd_sc_hd__buf_1
X_13960_ net7648 net1331 _06187_ VGND VGND VPWR VPWR _06225_ sky130_fd_sc_hd__a21o_1
Xwire2267 net2268 VGND VGND VPWR VPWR net2267 sky130_fd_sc_hd__clkbuf_1
X_21069_ _01037_ _01038_ VGND VGND VPWR VPWR _01085_ sky130_fd_sc_hd__xnor2_1
Xwire1522 _07975_ VGND VGND VPWR VPWR net1522 sky130_fd_sc_hd__buf_1
Xwire2278 _06515_ VGND VGND VPWR VPWR net2278 sky130_fd_sc_hd__buf_2
Xwire1533 net1534 VGND VGND VPWR VPWR net1533 sky130_fd_sc_hd__clkbuf_1
Xwire1544 _07277_ VGND VGND VPWR VPWR net1544 sky130_fd_sc_hd__buf_1
Xwire2289 net2290 VGND VGND VPWR VPWR net2289 sky130_fd_sc_hd__buf_1
Xwire1555 net1556 VGND VGND VPWR VPWR net1555 sky130_fd_sc_hd__clkbuf_1
X_12911_ _05168_ _05169_ net850 VGND VGND VPWR VPWR _05184_ sky130_fd_sc_hd__a21o_1
Xwire1566 net1567 VGND VGND VPWR VPWR net1566 sky130_fd_sc_hd__buf_1
X_25877_ clknet_leaf_14_clk _00750_ net8620 VGND VGND VPWR VPWR pid_q.ki\[5\] sky130_fd_sc_hd__dfrtp_1
X_13891_ _06142_ _06153_ _06155_ net449 VGND VGND VPWR VPWR _06157_ sky130_fd_sc_hd__o2bb2a_1
Xwire1577 net1578 VGND VGND VPWR VPWR net1577 sky130_fd_sc_hd__buf_1
Xwire1588 net1589 VGND VGND VPWR VPWR net1588 sky130_fd_sc_hd__buf_1
Xwire1599 net1600 VGND VGND VPWR VPWR net1599 sky130_fd_sc_hd__clkbuf_1
X_15630_ _07696_ _07701_ VGND VGND VPWR VPWR _07702_ sky130_fd_sc_hd__xnor2_1
X_24828_ net7480 net1640 _03575_ VGND VGND VPWR VPWR _04647_ sky130_fd_sc_hd__a21o_1
X_12842_ _05112_ _05113_ _05108_ _05109_ VGND VGND VPWR VPWR _05115_ sky130_fd_sc_hd__a211o_1
XFILLER_0_90_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15561_ _07631_ _07633_ VGND VGND VPWR VPWR _07634_ sky130_fd_sc_hd__xor2_1
XFILLER_0_61_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24759_ net5245 net2390 VGND VGND VPWR VPWR _04589_ sky130_fd_sc_hd__nand2_1
X_12773_ _05043_ net1147 VGND VGND VPWR VPWR _05046_ sky130_fd_sc_hd__xor2_1
XFILLER_0_96_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17300_ net7661 net7643 _09213_ VGND VGND VPWR VPWR _09214_ sky130_fd_sc_hd__or3_2
X_14512_ net7313 net5269 _06685_ VGND VGND VPWR VPWR _06693_ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18280_ _10129_ _10130_ VGND VGND VPWR VPWR _10131_ sky130_fd_sc_hd__nor2_1
X_15492_ _07543_ _07563_ _07564_ _07546_ VGND VGND VPWR VPWR _07565_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17231_ net3280 net1502 VGND VGND VPWR VPWR _09179_ sky130_fd_sc_hd__nand2_1
XFILLER_0_193_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14443_ _06636_ VGND VGND VPWR VPWR _00095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17162_ net1801 _09114_ net1076 VGND VGND VPWR VPWR _09115_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_107_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14374_ _06583_ matmul0.a_in\[12\] net900 VGND VGND VPWR VPWR _06584_ sky130_fd_sc_hd__mux2_1
Xwire830 _07166_ VGND VGND VPWR VPWR net830 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_49_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire841 _06045_ VGND VGND VPWR VPWR net841 sky130_fd_sc_hd__buf_1
Xwire852 net853 VGND VGND VPWR VPWR net852 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire863 net864 VGND VGND VPWR VPWR net863 sky130_fd_sc_hd__buf_1
X_16113_ net2712 net2239 VGND VGND VPWR VPWR _08179_ sky130_fd_sc_hd__nand2_1
X_13325_ _05596_ _05597_ VGND VGND VPWR VPWR _05598_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire874 net875 VGND VGND VPWR VPWR net874 sky130_fd_sc_hd__buf_1
X_17093_ net6974 VGND VGND VPWR VPWR _09050_ sky130_fd_sc_hd__inv_2
Xmax_length461 _04184_ VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire885 net886 VGND VGND VPWR VPWR net885 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire896 _06606_ VGND VGND VPWR VPWR net896 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_161_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16044_ _08105_ _08110_ VGND VGND VPWR VPWR _08111_ sky130_fd_sc_hd__xnor2_1
X_13256_ net6672 net6678 net7208 VGND VGND VPWR VPWR _05529_ sky130_fd_sc_hd__and3b_1
XFILLER_0_0_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13187_ _05458_ _05459_ VGND VGND VPWR VPWR _05460_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4170 net4172 VGND VGND VPWR VPWR net4170 sky130_fd_sc_hd__buf_1
X_19803_ net6151 _11582_ _11636_ VGND VGND VPWR VPWR _11637_ sky130_fd_sc_hd__nand3_1
Xwire4181 net4182 VGND VGND VPWR VPWR net4181 sky130_fd_sc_hd__buf_1
XFILLER_0_19_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4192 _06992_ VGND VGND VPWR VPWR net4192 sky130_fd_sc_hd__buf_1
X_17995_ net6940 _09843_ VGND VGND VPWR VPWR _09846_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19734_ _11565_ _11568_ net6084 VGND VGND VPWR VPWR _11569_ sky130_fd_sc_hd__o21ai_1
X_16946_ net2180 _08908_ net3351 VGND VGND VPWR VPWR _08910_ sky130_fd_sc_hd__a21o_1
Xwire3491 _07137_ VGND VGND VPWR VPWR net3491 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_1_clk clknet_4_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_16
Xwire2790 _07134_ VGND VGND VPWR VPWR net2790 sky130_fd_sc_hd__buf_1
XFILLER_0_189_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19665_ net3136 _11448_ VGND VGND VPWR VPWR _11501_ sky130_fd_sc_hd__or2_2
X_16877_ net2932 VGND VGND VPWR VPWR _08841_ sky130_fd_sc_hd__clkbuf_1
X_18616_ net2128 _10462_ net1762 VGND VGND VPWR VPWR _10463_ sky130_fd_sc_hd__a21o_1
X_15828_ _07864_ _07866_ VGND VGND VPWR VPWR _07898_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19596_ _11388_ VGND VGND VPWR VPWR _11433_ sky130_fd_sc_hd__inv_2
X_18547_ _10328_ _10394_ _10346_ VGND VGND VPWR VPWR _10396_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15759_ matmul0.matmul_stage_inst.mult1\[3\] net426 net2680 VGND VGND VPWR VPWR _07830_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18478_ net1208 net1441 _10327_ VGND VGND VPWR VPWR _10328_ sky130_fd_sc_hd__nand3_1
XFILLER_0_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17429_ _09328_ VGND VGND VPWR VPWR _00389_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20440_ net6369 _12233_ VGND VGND VPWR VPWR _12234_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20371_ net3355 cordic0.slte0.opA\[7\] net1228 _12170_ VGND VGND VPWR VPWR _00490_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22110_ _02081_ _02090_ _02091_ VGND VGND VPWR VPWR _02116_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23090_ _02956_ _02959_ VGND VGND VPWR VPWR _02960_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22041_ _02045_ _02047_ VGND VGND VPWR VPWR _02048_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_167_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25800_ clknet_leaf_30_clk _00673_ net8677 VGND VGND VPWR VPWR pid_q.curr_int\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_103_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23992_ _03854_ _03855_ VGND VGND VPWR VPWR _03856_ sky130_fd_sc_hd__nand2_1
X_25731_ clknet_leaf_9_clk _00604_ net8560 VGND VGND VPWR VPWR pid_d.ki\[5\] sky130_fd_sc_hd__dfrtp_1
X_22943_ pid_d.out\[14\] _02828_ _02831_ VGND VGND VPWR VPWR _02832_ sky130_fd_sc_hd__mux2_1
X_25662_ clknet_leaf_121_clk _00535_ net8406 VGND VGND VPWR VPWR pid_d.prev_error\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_74_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22874_ _01819_ _02762_ _02769_ VGND VGND VPWR VPWR _02770_ sky130_fd_sc_hd__a21o_1
X_24613_ net1651 net2018 net1649 VGND VGND VPWR VPWR _04468_ sky130_fd_sc_hd__mux2_1
X_21825_ net5548 net5679 VGND VGND VPWR VPWR _01834_ sky130_fd_sc_hd__nand2_1
X_25593_ clknet_leaf_91_clk _00466_ net8427 VGND VGND VPWR VPWR cordic0.cos\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_148_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21756_ _01764_ _01765_ VGND VGND VPWR VPWR _01766_ sky130_fd_sc_hd__xor2_1
X_24544_ _04315_ _04399_ VGND VGND VPWR VPWR _04400_ sky130_fd_sc_hd__and2_1
Xwire8403 net8404 VGND VGND VPWR VPWR net8403 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_164_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20707_ net6763 _12269_ net2583 VGND VGND VPWR VPWR _12480_ sky130_fd_sc_hd__mux2_1
Xwire8436 net8437 VGND VGND VPWR VPWR net8436 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire7702 net7703 VGND VGND VPWR VPWR net7702 sky130_fd_sc_hd__dlymetal6s2s_1
X_24475_ net5173 pid_q.prev_int\[13\] VGND VGND VPWR VPWR _04332_ sky130_fd_sc_hd__or2_1
X_21687_ _01593_ _01697_ VGND VGND VPWR VPWR _01698_ sky130_fd_sc_hd__xnor2_2
Xwire8447 net8448 VGND VGND VPWR VPWR net8447 sky130_fd_sc_hd__buf_1
Xwire7713 net7714 VGND VGND VPWR VPWR net7713 sky130_fd_sc_hd__buf_1
XFILLER_0_0_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8458 net8457 VGND VGND VPWR VPWR net8458 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_19_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8469 net8468 VGND VGND VPWR VPWR net8469 sky130_fd_sc_hd__clkbuf_2
X_23426_ _03264_ net1167 VGND VGND VPWR VPWR _03296_ sky130_fd_sc_hd__and2_1
Xwire7735 net7736 VGND VGND VPWR VPWR net7735 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20638_ _12295_ net3846 net2592 VGND VGND VPWR VPWR _12417_ sky130_fd_sc_hd__mux2_1
Xfanout6939 cordic0.vec\[1\]\[9\] VGND VGND VPWR VPWR net6939 sky130_fd_sc_hd__clkbuf_1
Xwire7746 net7747 VGND VGND VPWR VPWR net7746 sky130_fd_sc_hd__buf_1
XFILLER_0_163_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7757 net7758 VGND VGND VPWR VPWR net7757 sky130_fd_sc_hd__buf_1
XFILLER_0_110_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2710 _07309_ VGND VGND VPWR VPWR net2710 sky130_fd_sc_hd__clkbuf_1
Xwire159 net160 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23357_ _03221_ _03226_ VGND VGND VPWR VPWR _03227_ sky130_fd_sc_hd__xnor2_2
Xwire7779 net7783 VGND VGND VPWR VPWR net7779 sky130_fd_sc_hd__buf_1
Xmax_length2732 net2733 VGND VGND VPWR VPWR net2732 sky130_fd_sc_hd__buf_1
X_20569_ net6464 net3927 VGND VGND VPWR VPWR _12353_ sky130_fd_sc_hd__nand2_1
Xmax_length3488 net3489 VGND VGND VPWR VPWR net3488 sky130_fd_sc_hd__buf_1
XFILLER_0_33_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length2754 _07205_ VGND VGND VPWR VPWR net2754 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22308_ _02309_ _02311_ VGND VGND VPWR VPWR _02312_ sky130_fd_sc_hd__xor2_1
X_13110_ net7778 net2973 net2971 VGND VGND VPWR VPWR _05383_ sky130_fd_sc_hd__and3_1
X_14090_ _06284_ _06287_ _06288_ VGND VGND VPWR VPWR _06353_ sky130_fd_sc_hd__a21bo_1
Xmax_length2776 net2778 VGND VGND VPWR VPWR net2776 sky130_fd_sc_hd__buf_1
X_23288_ _03147_ _03157_ VGND VGND VPWR VPWR _03158_ sky130_fd_sc_hd__nand2_1
Xmax_length2798 _07129_ VGND VGND VPWR VPWR net2798 sky130_fd_sc_hd__clkbuf_1
X_13041_ _05184_ _05185_ net790 VGND VGND VPWR VPWR _05314_ sky130_fd_sc_hd__a21o_1
X_22239_ _02242_ _02243_ VGND VGND VPWR VPWR _02244_ sky130_fd_sc_hd__xnor2_1
X_25027_ _04779_ VGND VGND VPWR VPWR _04780_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2020 net2021 VGND VGND VPWR VPWR net2020 sky130_fd_sc_hd__buf_1
Xwire2031 net2032 VGND VGND VPWR VPWR net2031 sky130_fd_sc_hd__clkbuf_1
X_16800_ net8968 matmul0.cos\[3\] net3370 VGND VGND VPWR VPWR _08790_ sky130_fd_sc_hd__mux2_1
Xwire2042 _02548_ VGND VGND VPWR VPWR net2042 sky130_fd_sc_hd__buf_1
Xwire2053 net2054 VGND VGND VPWR VPWR net2053 sky130_fd_sc_hd__clkbuf_1
X_17780_ _09630_ _09607_ VGND VGND VPWR VPWR _09631_ sky130_fd_sc_hd__xnor2_1
Xwire2064 net2066 VGND VGND VPWR VPWR net2064 sky130_fd_sc_hd__buf_1
X_14992_ net4210 net4208 VGND VGND VPWR VPWR _07066_ sky130_fd_sc_hd__nor2_1
Xwire1330 _05526_ VGND VGND VPWR VPWR net1330 sky130_fd_sc_hd__buf_1
XFILLER_0_191_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2075 _01042_ VGND VGND VPWR VPWR net2075 sky130_fd_sc_hd__buf_1
Xwire2086 _12279_ VGND VGND VPWR VPWR net2086 sky130_fd_sc_hd__buf_1
X_16731_ matmul0.b_in\[2\] matmul0.b\[2\] net3703 VGND VGND VPWR VPWR _08754_ sky130_fd_sc_hd__mux2_1
X_13943_ _06205_ _06208_ VGND VGND VPWR VPWR _06209_ sky130_fd_sc_hd__xnor2_2
Xwire1352 net1353 VGND VGND VPWR VPWR net1352 sky130_fd_sc_hd__buf_1
X_25929_ clknet_leaf_2_clk _00802_ net8574 VGND VGND VPWR VPWR pid_d.prev_int\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire2097 net2098 VGND VGND VPWR VPWR net2097 sky130_fd_sc_hd__buf_1
Xwire1363 net1364 VGND VGND VPWR VPWR net1363 sky130_fd_sc_hd__clkbuf_1
Xwire1374 _04510_ VGND VGND VPWR VPWR net1374 sky130_fd_sc_hd__buf_1
Xwire1385 net1386 VGND VGND VPWR VPWR net1385 sky130_fd_sc_hd__buf_1
X_19450_ _10982_ net2520 _10988_ VGND VGND VPWR VPWR _11287_ sky130_fd_sc_hd__a21o_1
Xwire1396 net1397 VGND VGND VPWR VPWR net1396 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16662_ matmul0.alpha_pass\[6\] net972 net6563 VGND VGND VPWR VPWR _08697_ sky130_fd_sc_hd__mux2_1
X_13874_ _06137_ _06140_ VGND VGND VPWR VPWR _06141_ sky130_fd_sc_hd__xor2_1
X_18401_ net3926 _10250_ _10206_ _10251_ VGND VGND VPWR VPWR _10252_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15613_ net2851 net4076 net3397 net3444 VGND VGND VPWR VPWR _07685_ sky130_fd_sc_hd__a2bb2o_1
X_12825_ _05094_ _05097_ VGND VGND VPWR VPWR _05098_ sky130_fd_sc_hd__xnor2_1
X_19381_ net6218 _11208_ _11215_ _11217_ VGND VGND VPWR VPWR _11218_ sky130_fd_sc_hd__o22a_1
X_16593_ svm0.state\[1\] svm0.state\[0\] VGND VGND VPWR VPWR _08644_ sky130_fd_sc_hd__or2_1
XFILLER_0_189_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18332_ _10090_ net1777 net2138 VGND VGND VPWR VPWR _10183_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_167_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15544_ _07613_ _07616_ VGND VGND VPWR VPWR _07617_ sky130_fd_sc_hd__xnor2_2
X_12756_ _04994_ _05028_ VGND VGND VPWR VPWR _05029_ sky130_fd_sc_hd__xnor2_1
Xmax_length6070 net6071 VGND VGND VPWR VPWR net6070 sky130_fd_sc_hd__buf_1
XFILLER_0_16_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18263_ _10106_ _10107_ net2138 VGND VGND VPWR VPWR _10114_ sky130_fd_sc_hd__a21o_1
X_15475_ net1274 _07545_ VGND VGND VPWR VPWR _07549_ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12687_ net2330 net2325 VGND VGND VPWR VPWR _04960_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17214_ net966 _09145_ _09142_ VGND VGND VPWR VPWR _09163_ sky130_fd_sc_hd__a21oi_2
X_14426_ _06623_ matmul0.b_in\[8\] net897 VGND VGND VPWR VPWR _06624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18194_ net6920 net6949 VGND VGND VPWR VPWR _10045_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17145_ net6483 _09094_ _09096_ net3341 _09098_ VGND VGND VPWR VPWR _09099_ sky130_fd_sc_hd__a221o_1
X_14357_ net8204 _06527_ VGND VGND VPWR VPWR _06570_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire660 net661 VGND VGND VPWR VPWR net660 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire671 _08536_ VGND VGND VPWR VPWR net671 sky130_fd_sc_hd__clkbuf_1
Xwire682 _05470_ VGND VGND VPWR VPWR net682 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire693 _04050_ VGND VGND VPWR VPWR net693 sky130_fd_sc_hd__clkbuf_1
X_13308_ net1574 _05580_ VGND VGND VPWR VPWR _05581_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17076_ net6485 net2598 net6473 VGND VGND VPWR VPWR _09034_ sky130_fd_sc_hd__o21ai_1
X_14288_ net77 _06518_ _06519_ net7791 VGND VGND VPWR VPWR _00057_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16027_ net2708 net3400 VGND VGND VPWR VPWR _08094_ sky130_fd_sc_hd__nor2_1
X_13239_ _05441_ _05443_ _05442_ VGND VGND VPWR VPWR _05512_ sky130_fd_sc_hd__a21o_1
XFILLER_0_196_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_127_Right_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17978_ net1214 net1447 VGND VGND VPWR VPWR _09829_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16929_ net6418 _08891_ VGND VGND VPWR VPWR _08893_ sky130_fd_sc_hd__or2_1
X_19717_ net9029 net1199 _11552_ net1767 VGND VGND VPWR VPWR _00454_ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19648_ _11426_ _11484_ VGND VGND VPWR VPWR _11485_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19579_ _11413_ _11415_ VGND VGND VPWR VPWR _11416_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_172_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21610_ net5427 net5888 _01508_ VGND VGND VPWR VPWR _01622_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22590_ net3091 _02566_ _02567_ VGND VGND VPWR VPWR _02568_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21541_ _01501_ net1049 net1180 VGND VGND VPWR VPWR _01553_ sky130_fd_sc_hd__a21bo_1
Xwire7009 net7011 VGND VGND VPWR VPWR net7009 sky130_fd_sc_hd__clkbuf_1
X_24260_ net793 _04095_ _04088_ VGND VGND VPWR VPWR _04120_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21472_ net5843 net5458 VGND VGND VPWR VPWR _01485_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6308 net6306 VGND VGND VPWR VPWR net6308 sky130_fd_sc_hd__buf_1
XFILLER_0_15_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23211_ net5070 net4778 _03080_ VGND VGND VPWR VPWR _03081_ sky130_fd_sc_hd__a21o_1
XFILLER_0_145_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6319 net6316 VGND VGND VPWR VPWR net6319 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_7_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20423_ _12205_ _12210_ cordic0.slte0.opA\[10\] VGND VGND VPWR VPWR _12219_ sky130_fd_sc_hd__o21a_1
X_24191_ _04051_ _04001_ _03978_ VGND VGND VPWR VPWR _04052_ sky130_fd_sc_hd__o21a_1
Xwire5607 net5600 VGND VGND VPWR VPWR net5607 sky130_fd_sc_hd__buf_1
Xwire5618 net5619 VGND VGND VPWR VPWR net5618 sky130_fd_sc_hd__buf_1
Xwire5629 net5628 VGND VGND VPWR VPWR net5629 sky130_fd_sc_hd__buf_1
XFILLER_0_30_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23142_ net5112 net4681 VGND VGND VPWR VPWR _03012_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20354_ _12140_ _12148_ _12149_ cordic0.slte0.opA\[5\] VGND VGND VPWR VPWR _12155_
+ sky130_fd_sc_hd__a31o_1
Xwire4906 net4907 VGND VGND VPWR VPWR net4906 sky130_fd_sc_hd__buf_1
Xwire4917 net4918 VGND VGND VPWR VPWR net4917 sky130_fd_sc_hd__buf_1
XFILLER_0_105_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23073_ _02941_ _02942_ VGND VGND VPWR VPWR _02943_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_178_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20285_ net6499 _12090_ net1824 VGND VGND VPWR VPWR _12091_ sky130_fd_sc_hd__mux2_1
X_22024_ net5746 net5433 VGND VGND VPWR VPWR _02031_ sky130_fd_sc_hd__nand2_1
Xhold12 matmul0.matmul_stage_inst.a\[9\] VGND VGND VPWR VPWR net8965 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 matmul0.matmul_stage_inst.start VGND VGND VPWR VPWR net8976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 pid_d.curr_error\[0\] VGND VGND VPWR VPWR net8987 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 cordic0.out_valid VGND VGND VPWR VPWR net8998 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 pid_d.curr_int\[1\] VGND VGND VPWR VPWR net9009 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 matmul0.matmul_stage_inst.d\[5\] VGND VGND VPWR VPWR net9020 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 matmul0.matmul_stage_inst.b\[4\] VGND VGND VPWR VPWR net9031 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23975_ _03734_ _03746_ _03838_ VGND VGND VPWR VPWR _03839_ sky130_fd_sc_hd__o21ai_1
Xhold89 pid_q.target\[13\] VGND VGND VPWR VPWR net9042 sky130_fd_sc_hd__dlygate4sd3_1
X_25714_ clknet_leaf_9_clk _00587_ net8559 VGND VGND VPWR VPWR pid_d.mult0.a\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22926_ net295 _02793_ VGND VGND VPWR VPWR _02817_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25645_ clknet_leaf_100_clk _00518_ net8390 VGND VGND VPWR VPWR cordic0.vec\[0\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_22857_ _02752_ _02753_ VGND VGND VPWR VPWR _02755_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12610_ net8909 net4341 VGND VGND VPWR VPWR _04885_ sky130_fd_sc_hd__and2_1
XFILLER_0_183_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21808_ net9243 net3123 net2078 _01817_ VGND VGND VPWR VPWR _00525_ sky130_fd_sc_hd__a22o_1
X_13590_ _05849_ _05770_ net504 VGND VGND VPWR VPWR _05860_ sky130_fd_sc_hd__or3b_1
X_25576_ clknet_leaf_97_clk _00449_ net8385 VGND VGND VPWR VPWR cordic0.sin\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_22788_ pid_d.kp\[6\] _02674_ net1681 VGND VGND VPWR VPWR _02702_ sky130_fd_sc_hd__mux2_1
Xwire8200 net8201 VGND VGND VPWR VPWR net8200 sky130_fd_sc_hd__clkbuf_1
Xwire8211 net8212 VGND VGND VPWR VPWR net8211 sky130_fd_sc_hd__clkbuf_1
X_24527_ _04321_ _04325_ _04322_ VGND VGND VPWR VPWR _04384_ sky130_fd_sc_hd__a21bo_1
Xwire8222 net8223 VGND VGND VPWR VPWR net8222 sky130_fd_sc_hd__clkbuf_1
X_21739_ _01135_ net5645 VGND VGND VPWR VPWR _01749_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8233 net8234 VGND VGND VPWR VPWR net8233 sky130_fd_sc_hd__clkbuf_1
Xwire8244 net8245 VGND VGND VPWR VPWR net8244 sky130_fd_sc_hd__clkbuf_1
Xfanout7448 net7449 VGND VGND VPWR VPWR net7448 sky130_fd_sc_hd__buf_2
XFILLER_0_47_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8255 net8256 VGND VGND VPWR VPWR net8255 sky130_fd_sc_hd__clkbuf_1
X_15260_ _07280_ _07333_ VGND VGND VPWR VPWR _07334_ sky130_fd_sc_hd__xnor2_1
Xwire8266 net8267 VGND VGND VPWR VPWR net8266 sky130_fd_sc_hd__clkbuf_1
X_24458_ _04314_ _04315_ VGND VGND VPWR VPWR _04316_ sky130_fd_sc_hd__nand2_1
Xwire7532 net7533 VGND VGND VPWR VPWR net7532 sky130_fd_sc_hd__clkbuf_1
Xwire8277 net8278 VGND VGND VPWR VPWR net8277 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7543 net7544 VGND VGND VPWR VPWR net7543 sky130_fd_sc_hd__clkbuf_1
Xwire8288 net8289 VGND VGND VPWR VPWR net8288 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14211_ _06445_ _06467_ _06469_ _06447_ VGND VGND VPWR VPWR _06470_ sky130_fd_sc_hd__o2bb2a_2
Xwire8299 net20 VGND VGND VPWR VPWR net8299 sky130_fd_sc_hd__clkbuf_1
Xwire7554 net7555 VGND VGND VPWR VPWR net7554 sky130_fd_sc_hd__clkbuf_1
X_23409_ _03277_ _03278_ VGND VGND VPWR VPWR _03279_ sky130_fd_sc_hd__or2b_1
Xwire7565 matmul0.b_in\[10\] VGND VGND VPWR VPWR net7565 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout6769 net6772 VGND VGND VPWR VPWR net6769 sky130_fd_sc_hd__buf_1
X_15191_ _07235_ _07261_ _07262_ _07264_ VGND VGND VPWR VPWR _07265_ sky130_fd_sc_hd__o2bb2a_1
Xmax_length3263 _09620_ VGND VGND VPWR VPWR net3263 sky130_fd_sc_hd__clkbuf_2
X_24389_ _04162_ _04164_ _04247_ VGND VGND VPWR VPWR _04248_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire6842 net6839 VGND VGND VPWR VPWR net6842 sky130_fd_sc_hd__clkbuf_2
Xwire7587 net7588 VGND VGND VPWR VPWR net7587 sky130_fd_sc_hd__clkbuf_1
Xwire6853 net6850 VGND VGND VPWR VPWR net6853 sky130_fd_sc_hd__buf_1
Xmax_length3285 net3286 VGND VGND VPWR VPWR net3285 sky130_fd_sc_hd__buf_1
Xwire7598 net7599 VGND VGND VPWR VPWR net7598 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14142_ _06384_ _06391_ VGND VGND VPWR VPWR _06403_ sky130_fd_sc_hd__nor2_2
Xwire6864 net6865 VGND VGND VPWR VPWR net6864 sky130_fd_sc_hd__buf_1
XFILLER_0_85_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6875 net6872 VGND VGND VPWR VPWR net6875 sky130_fd_sc_hd__clkbuf_2
Xmax_length2573 net2574 VGND VGND VPWR VPWR net2573 sky130_fd_sc_hd__buf_1
Xwire6886 net6883 VGND VGND VPWR VPWR net6886 sky130_fd_sc_hd__buf_1
XFILLER_0_104_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6897 net6900 VGND VGND VPWR VPWR net6897 sky130_fd_sc_hd__clkbuf_2
X_14073_ net1332 _06174_ _06333_ _06221_ net7625 VGND VGND VPWR VPWR _06336_ sky130_fd_sc_hd__o32a_1
X_18950_ net6194 VGND VGND VPWR VPWR _10787_ sky130_fd_sc_hd__inv_2
X_13024_ net7933 _05296_ net1592 _05294_ VGND VGND VPWR VPWR _05297_ sky130_fd_sc_hd__o22a_1
X_17901_ _09695_ _09742_ VGND VGND VPWR VPWR _09752_ sky130_fd_sc_hd__xnor2_1
X_18881_ _10705_ _10722_ VGND VGND VPWR VPWR _10723_ sky130_fd_sc_hd__xnor2_2
X_17832_ net7032 _09679_ _09681_ _09648_ net3974 VGND VGND VPWR VPWR _09683_ sky130_fd_sc_hd__a221o_1
XFILLER_0_174_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17763_ net7121 net7133 VGND VGND VPWR VPWR _09614_ sky130_fd_sc_hd__nand2b_1
X_14975_ net4170 net4165 net4175 net4173 VGND VGND VPWR VPWR _07049_ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1160 _03923_ VGND VGND VPWR VPWR net1160 sky130_fd_sc_hd__buf_1
Xwire1171 _01858_ VGND VGND VPWR VPWR net1171 sky130_fd_sc_hd__buf_1
XFILLER_0_107_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19502_ _11335_ _11338_ VGND VGND VPWR VPWR _11339_ sky130_fd_sc_hd__xnor2_1
X_16714_ _08740_ _08736_ net7375 VGND VGND VPWR VPWR _08741_ sky130_fd_sc_hd__o21ba_1
X_13926_ net7721 net1581 VGND VGND VPWR VPWR _06192_ sky130_fd_sc_hd__and2_1
Xwire1182 _01372_ VGND VGND VPWR VPWR net1182 sky130_fd_sc_hd__clkbuf_2
X_17694_ svm0.state\[1\] net5185 _09187_ net3387 VGND VGND VPWR VPWR _00410_ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1193 _11081_ VGND VGND VPWR VPWR net1193 sky130_fd_sc_hd__buf_1
XFILLER_0_18_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19433_ _11267_ _11269_ VGND VGND VPWR VPWR _11270_ sky130_fd_sc_hd__xor2_1
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16645_ matmul0.matmul_stage_inst.mult1\[3\] _08675_ _08681_ VGND VGND VPWR VPWR
+ _08682_ sky130_fd_sc_hd__a21boi_2
X_13857_ net837 net907 VGND VGND VPWR VPWR _06124_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_190_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12808_ _04979_ _04997_ _05080_ VGND VGND VPWR VPWR _05081_ sky130_fd_sc_hd__o21a_1
X_19364_ _11186_ _11198_ VGND VGND VPWR VPWR _11201_ sky130_fd_sc_hd__xor2_1
XFILLER_0_128_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16576_ matmul0.matmul_stage_inst.mult1\[15\] net161 net3474 VGND VGND VPWR VPWR
+ _08635_ sky130_fd_sc_hd__mux2_1
X_13788_ _06052_ _06055_ VGND VGND VPWR VPWR _06056_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18315_ net3347 _09606_ net3226 VGND VGND VPWR VPWR _10166_ sky130_fd_sc_hd__a21oi_1
X_15527_ _07517_ _07518_ _07599_ VGND VGND VPWR VPWR _07600_ sky130_fd_sc_hd__o21a_1
XFILLER_0_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12739_ _05011_ VGND VGND VPWR VPWR _05012_ sky130_fd_sc_hd__buf_1
X_19295_ _10946_ VGND VGND VPWR VPWR _11132_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8661 net8664 VGND VGND VPWR VPWR net8661 sky130_fd_sc_hd__buf_1
XFILLER_0_155_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18246_ net7075 net7098 net7014 VGND VGND VPWR VPWR _10097_ sky130_fd_sc_hd__a21o_1
XFILLER_0_155_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15458_ net2814 _07063_ _07382_ _07383_ VGND VGND VPWR VPWR _07532_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14409_ net5282 net1295 net2891 net4452 _06610_ VGND VGND VPWR VPWR _06611_ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18177_ _09817_ _10024_ _10026_ _10027_ VGND VGND VPWR VPWR _10028_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15389_ _07313_ _07454_ net990 VGND VGND VPWR VPWR _07463_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17128_ net5990 net2169 _09082_ VGND VGND VPWR VPWR _09083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire490 _08378_ VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17059_ net3328 _09017_ net3336 VGND VGND VPWR VPWR _09018_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20070_ _11863_ net2494 VGND VGND VPWR VPWR _11899_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23760_ _03624_ _03625_ VGND VGND VPWR VPWR _03626_ sky130_fd_sc_hd__xnor2_1
X_20972_ net5602 net5868 VGND VGND VPWR VPWR _00988_ sky130_fd_sc_hd__nand2_1
XFILLER_0_196_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22711_ pid_d.ki\[14\] net3705 _04886_ pid_d.kp\[14\] VGND VGND VPWR VPWR _02649_
+ sky130_fd_sc_hd__a22o_1
Xmax_length6806 net6803 VGND VGND VPWR VPWR net6806 sky130_fd_sc_hd__buf_1
XFILLER_0_79_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23691_ _03556_ _03557_ VGND VGND VPWR VPWR _03558_ sky130_fd_sc_hd__or2b_1
Xmax_length6817 net6818 VGND VGND VPWR VPWR net6817 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_177_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25430_ clknet_leaf_97_clk _00313_ net8399 VGND VGND VPWR VPWR matmul0.sin\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22642_ net5860 net3083 VGND VGND VPWR VPWR _02606_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25361_ clknet_leaf_72_clk _00244_ net8477 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult2\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_22573_ net7329 _02551_ VGND VGND VPWR VPWR _02554_ sky130_fd_sc_hd__or2_1
XFILLER_0_192_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24312_ pid_q.curr_int\[9\] VGND VGND VPWR VPWR _04172_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21524_ _01535_ _01536_ VGND VGND VPWR VPWR _01537_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25292_ clknet_leaf_77_clk _00175_ net8438 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.d\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6105 net6106 VGND VGND VPWR VPWR net6105 sky130_fd_sc_hd__clkbuf_2
Xwire6116 net6113 VGND VGND VPWR VPWR net6116 sky130_fd_sc_hd__buf_1
X_24243_ net692 _04103_ VGND VGND VPWR VPWR _04104_ sky130_fd_sc_hd__xnor2_1
X_21455_ net5777 net5511 VGND VGND VPWR VPWR _01468_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6149 net6150 VGND VGND VPWR VPWR net6149 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20406_ net6485 net4050 _12109_ VGND VGND VPWR VPWR _12203_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5415 net5416 VGND VGND VPWR VPWR net5415 sky130_fd_sc_hd__buf_1
XFILLER_0_181_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24174_ net7525 _03959_ net241 net7467 net636 VGND VGND VPWR VPWR _04036_ sky130_fd_sc_hd__a221o_1
Xwire5426 net5427 VGND VGND VPWR VPWR net5426 sky130_fd_sc_hd__buf_1
XFILLER_0_160_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21386_ _01270_ _01274_ _01399_ VGND VGND VPWR VPWR _01400_ sky130_fd_sc_hd__o21ai_1
Xwire4703 net4704 VGND VGND VPWR VPWR net4703 sky130_fd_sc_hd__buf_1
Xwire5448 net5449 VGND VGND VPWR VPWR net5448 sky130_fd_sc_hd__buf_1
XFILLER_0_120_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4714 pid_q.mult0.a\[4\] VGND VGND VPWR VPWR net4714 sky130_fd_sc_hd__buf_1
X_23125_ _02911_ _02994_ VGND VGND VPWR VPWR _02995_ sky130_fd_sc_hd__xnor2_1
Xwire4725 net4726 VGND VGND VPWR VPWR net4725 sky130_fd_sc_hd__clkbuf_1
X_20337_ _12126_ _12138_ _12137_ VGND VGND VPWR VPWR _12140_ sky130_fd_sc_hd__a21o_1
Xwire4736 net4737 VGND VGND VPWR VPWR net4736 sky130_fd_sc_hd__buf_1
Xwire4747 net4744 VGND VGND VPWR VPWR net4747 sky130_fd_sc_hd__buf_1
Xwire4758 net4753 VGND VGND VPWR VPWR net4758 sky130_fd_sc_hd__buf_1
Xwire4769 net4770 VGND VGND VPWR VPWR net4769 sky130_fd_sc_hd__clkbuf_1
X_23056_ net4772 net4742 net4913 VGND VGND VPWR VPWR _02926_ sky130_fd_sc_hd__and3b_1
X_20268_ _12078_ VGND VGND VPWR VPWR _00479_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput102 pid_d_data[14] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_1
X_22007_ net4383 net698 net347 net4319 _02014_ VGND VGND VPWR VPWR _02015_ sky130_fd_sc_hd__a221o_1
Xinput113 pid_d_wen VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_1
Xinput124 pid_q_addr[4] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_1
X_20199_ net6042 net6000 _12023_ net6063 net6034 VGND VGND VPWR VPWR _12024_ sky130_fd_sc_hd__a221o_1
Xinput135 pid_q_data[14] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_1
Xinput146 pid_q_wen VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_1
Xmax_length8720 net8721 VGND VGND VPWR VPWR net8720 sky130_fd_sc_hd__buf_1
X_14760_ net3615 _06842_ VGND VGND VPWR VPWR _06890_ sky130_fd_sc_hd__and2_1
X_23958_ _03699_ _03821_ VGND VGND VPWR VPWR _03822_ sky130_fd_sc_hd__xor2_2
XFILLER_0_187_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length8775 net8776 VGND VGND VPWR VPWR net8775 sky130_fd_sc_hd__buf_1
X_13711_ _05911_ _05912_ VGND VGND VPWR VPWR _05980_ sky130_fd_sc_hd__and2_1
X_22909_ _02183_ _02797_ pid_d.out\[10\] VGND VGND VPWR VPWR _02801_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_6_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14691_ net3630 VGND VGND VPWR VPWR _06838_ sky130_fd_sc_hd__clkbuf_1
X_23889_ _03753_ VGND VGND VPWR VPWR _03754_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16430_ net490 net571 VGND VGND VPWR VPWR _08491_ sky130_fd_sc_hd__nor2_1
X_13642_ net1573 _05828_ net7617 net1347 VGND VGND VPWR VPWR _05912_ sky130_fd_sc_hd__o211a_1
X_25628_ clknet_leaf_104_clk _00501_ net8357 VGND VGND VPWR VPWR cordic0.vec\[0\]\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_78_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16361_ _08413_ _08423_ VGND VGND VPWR VPWR _08424_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_184_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13573_ net916 net913 _05843_ VGND VGND VPWR VPWR _05844_ sky130_fd_sc_hd__o21a_1
X_25559_ clknet_leaf_115_clk _00432_ net8335 VGND VGND VPWR VPWR cordic0.gm0.iter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8030 net8031 VGND VGND VPWR VPWR net8030 sky130_fd_sc_hd__clkbuf_1
X_18100_ _09754_ _09753_ VGND VGND VPWR VPWR _09951_ sky130_fd_sc_hd__xnor2_1
X_15312_ net1539 net1869 VGND VGND VPWR VPWR _07386_ sky130_fd_sc_hd__xnor2_2
X_19080_ net6247 net6328 VGND VGND VPWR VPWR _10917_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8052 net8053 VGND VGND VPWR VPWR net8052 sky130_fd_sc_hd__buf_1
X_16292_ _08353_ net724 VGND VGND VPWR VPWR _08356_ sky130_fd_sc_hd__nor2_1
Xwire8063 net8058 VGND VGND VPWR VPWR net8063 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8074 net8064 VGND VGND VPWR VPWR net8074 sky130_fd_sc_hd__buf_1
Xwire8085 _02657_ VGND VGND VPWR VPWR net8085 sky130_fd_sc_hd__clkbuf_1
Xwire7340 net7341 VGND VGND VPWR VPWR net7340 sky130_fd_sc_hd__buf_1
X_18031_ _09875_ _09881_ VGND VGND VPWR VPWR _09882_ sky130_fd_sc_hd__xnor2_1
Xfanout6544 net6566 VGND VGND VPWR VPWR net6544 sky130_fd_sc_hd__buf_1
Xwire8096 net8097 VGND VGND VPWR VPWR net8096 sky130_fd_sc_hd__clkbuf_1
X_15243_ _07195_ _07284_ VGND VGND VPWR VPWR _07317_ sky130_fd_sc_hd__xnor2_1
Xwire7351 matmul0.alpha_pass\[2\] VGND VGND VPWR VPWR net7351 sky130_fd_sc_hd__buf_1
Xwire7362 net7363 VGND VGND VPWR VPWR net7362 sky130_fd_sc_hd__buf_1
XFILLER_0_83_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7373 matmul0.alpha_pass\[0\] VGND VGND VPWR VPWR net7373 sky130_fd_sc_hd__buf_1
XFILLER_0_151_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire7384 matmul0.matmul_stage_inst.f\[6\] VGND VGND VPWR VPWR net7384 sky130_fd_sc_hd__clkbuf_1
Xwire6650 net6651 VGND VGND VPWR VPWR net6650 sky130_fd_sc_hd__buf_1
Xwire6661 net6662 VGND VGND VPWR VPWR net6661 sky130_fd_sc_hd__buf_1
X_15174_ net2849 net3453 _07247_ VGND VGND VPWR VPWR _07248_ sky130_fd_sc_hd__a21o_1
Xwire6683 net151 VGND VGND VPWR VPWR net6683 sky130_fd_sc_hd__clkbuf_1
Xmax_length2370 _04895_ VGND VGND VPWR VPWR net2370 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14125_ _06221_ _06386_ net7613 VGND VGND VPWR VPWR _06387_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5960 net5962 VGND VGND VPWR VPWR net5960 sky130_fd_sc_hd__buf_1
X_19982_ _11768_ net1408 _11744_ VGND VGND VPWR VPWR _11813_ sky130_fd_sc_hd__o21a_1
Xwire5971 pid_d.curr_error\[2\] VGND VGND VPWR VPWR net5971 sky130_fd_sc_hd__clkbuf_2
Xwire5982 pid_d.curr_int\[3\] VGND VGND VPWR VPWR net5982 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire5993 net5991 VGND VGND VPWR VPWR net5993 sky130_fd_sc_hd__buf_1
X_14056_ _06280_ net366 VGND VGND VPWR VPWR _06320_ sky130_fd_sc_hd__xnor2_1
X_18933_ net275 _10747_ net245 VGND VGND VPWR VPWR _10772_ sky130_fd_sc_hd__or3_1
X_13007_ _05153_ _05154_ VGND VGND VPWR VPWR _05280_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18864_ net6812 net6770 _10677_ VGND VGND VPWR VPWR _10706_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17815_ net3248 _09665_ VGND VGND VPWR VPWR _09666_ sky130_fd_sc_hd__xor2_2
X_18795_ net3920 _10638_ VGND VGND VPWR VPWR _10639_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17746_ net8062 net2195 VGND VGND VPWR VPWR _09597_ sky130_fd_sc_hd__nand2_1
XFILLER_0_168_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14958_ _07024_ _07031_ VGND VGND VPWR VPWR _07032_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13909_ _06173_ net1950 _06174_ VGND VGND VPWR VPWR _06175_ sky130_fd_sc_hd__or3_1
XFILLER_0_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17677_ _09552_ _09556_ _09547_ VGND VGND VPWR VPWR _09557_ sky130_fd_sc_hd__o21ai_1
X_14889_ net6539 net6590 matmul0.matmul_stage_inst.e\[0\] VGND VGND VPWR VPWR _06963_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19416_ _11009_ _10994_ net1426 VGND VGND VPWR VPWR _11253_ sky130_fd_sc_hd__o21a_1
X_16628_ _08665_ _08666_ VGND VGND VPWR VPWR _08667_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19347_ net1421 _11183_ VGND VGND VPWR VPWR _11184_ sky130_fd_sc_hd__xnor2_2
X_16559_ net881 _08617_ VGND VGND VPWR VPWR _08618_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19278_ _10862_ _11114_ VGND VGND VPWR VPWR _11115_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18229_ net7144 _09809_ VGND VGND VPWR VPWR _10080_ sky130_fd_sc_hd__or2b_1
XFILLER_0_182_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21240_ _00838_ net1393 net1735 VGND VGND VPWR VPWR _01255_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_4_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21171_ net5634 net5882 _01172_ _01180_ _01186_ VGND VGND VPWR VPWR _01187_ sky130_fd_sc_hd__a41o_1
XFILLER_0_68_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20122_ _11895_ _11894_ _11887_ VGND VGND VPWR VPWR _11950_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2608 net2610 VGND VGND VPWR VPWR net2608 sky130_fd_sc_hd__buf_1
Xwire2619 net2620 VGND VGND VPWR VPWR net2619 sky130_fd_sc_hd__buf_1
X_24930_ net8867 net142 VGND VGND VPWR VPWR _04714_ sky130_fd_sc_hd__and2b_1
XFILLER_0_102_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20053_ _11861_ _11881_ VGND VGND VPWR VPWR _11882_ sky130_fd_sc_hd__nor2_1
Xwire1907 _06885_ VGND VGND VPWR VPWR net1907 sky130_fd_sc_hd__clkbuf_1
Xwire1918 net1919 VGND VGND VPWR VPWR net1918 sky130_fd_sc_hd__buf_1
Xwire1929 net1930 VGND VGND VPWR VPWR net1929 sky130_fd_sc_hd__buf_1
XFILLER_0_175_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24861_ pid_q.ki\[2\] net2397 net3009 pid_q.kp\[2\] VGND VGND VPWR VPWR _04665_ sky130_fd_sc_hd__a22o_1
XFILLER_0_175_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length8016 pid_q.target\[4\] VGND VGND VPWR VPWR net8016 sky130_fd_sc_hd__clkbuf_1
Xmax_length8027 pid_q.target\[2\] VGND VGND VPWR VPWR net8027 sky130_fd_sc_hd__clkbuf_1
X_23812_ _03584_ _03585_ _03658_ VGND VGND VPWR VPWR _03677_ sky130_fd_sc_hd__and3_1
X_24792_ net5167 net1643 _04543_ net372 VGND VGND VPWR VPWR _00709_ sky130_fd_sc_hd__a22o_1
XFILLER_0_169_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23743_ net5096 _03607_ _03608_ VGND VGND VPWR VPWR _03609_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20955_ net5613 net5792 net5635 VGND VGND VPWR VPWR _00971_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23674_ net1019 net1018 VGND VGND VPWR VPWR _03541_ sky130_fd_sc_hd__xnor2_1
Xmax_length6647 net6648 VGND VGND VPWR VPWR net6647 sky130_fd_sc_hd__clkbuf_1
X_20886_ net5558 net5869 VGND VGND VPWR VPWR _00902_ sky130_fd_sc_hd__nand2_1
XFILLER_0_193_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25413_ clknet_leaf_90_clk _00296_ net8420 VGND VGND VPWR VPWR matmul0.cos\[0\] sky130_fd_sc_hd__dfrtp_1
X_22625_ net3770 _02593_ _02594_ VGND VGND VPWR VPWR _02595_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25344_ clknet_leaf_73_clk _00227_ net8471 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_22556_ net9083 _02521_ _02540_ VGND VGND VPWR VPWR _00550_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21507_ _01447_ _01519_ VGND VGND VPWR VPWR _01520_ sky130_fd_sc_hd__xor2_1
Xfanout5117 net5127 VGND VGND VPWR VPWR net5117 sky130_fd_sc_hd__buf_1
X_25275_ clknet_leaf_93_clk _00158_ net8447 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.c\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_22487_ net5434 net5390 net5671 VGND VGND VPWR VPWR _02488_ sky130_fd_sc_hd__or3b_1
XFILLER_0_134_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5139 net5157 VGND VGND VPWR VPWR net5139 sky130_fd_sc_hd__buf_1
XFILLER_0_1_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5201 net5203 VGND VGND VPWR VPWR net5201 sky130_fd_sc_hd__clkbuf_1
Xmax_length857 net858 VGND VGND VPWR VPWR net857 sky130_fd_sc_hd__clkbuf_1
X_24226_ net1159 _04086_ VGND VGND VPWR VPWR _04087_ sky130_fd_sc_hd__xnor2_1
Xwire5223 net5224 VGND VGND VPWR VPWR net5223 sky130_fd_sc_hd__clkbuf_2
X_21438_ _01449_ _01450_ VGND VGND VPWR VPWR _01451_ sky130_fd_sc_hd__xnor2_1
Xwire5234 matmul0.beta_pass\[10\] VGND VGND VPWR VPWR net5234 sky130_fd_sc_hd__clkbuf_1
Xwire4500 net4501 VGND VGND VPWR VPWR net4500 sky130_fd_sc_hd__buf_1
Xwire5245 net5246 VGND VGND VPWR VPWR net5245 sky130_fd_sc_hd__buf_1
Xwire4511 net4512 VGND VGND VPWR VPWR net4511 sky130_fd_sc_hd__buf_1
Xwire5256 net5257 VGND VGND VPWR VPWR net5256 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24157_ net1160 _03927_ _03928_ VGND VGND VPWR VPWR _04019_ sky130_fd_sc_hd__o21a_1
Xwire4522 net4524 VGND VGND VPWR VPWR net4522 sky130_fd_sc_hd__buf_1
Xwire5267 net5269 VGND VGND VPWR VPWR net5267 sky130_fd_sc_hd__buf_1
XFILLER_0_82_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21369_ _01381_ _01382_ VGND VGND VPWR VPWR _01383_ sky130_fd_sc_hd__xor2_1
Xwire5289 matmul0.beta_pass\[3\] VGND VGND VPWR VPWR net5289 sky130_fd_sc_hd__buf_1
X_23108_ net4981 net4739 _02976_ _02977_ VGND VGND VPWR VPWR _02978_ sky130_fd_sc_hd__a31o_1
Xwire4555 net4551 VGND VGND VPWR VPWR net4555 sky130_fd_sc_hd__clkbuf_2
Xwire3810 net3811 VGND VGND VPWR VPWR net3810 sky130_fd_sc_hd__clkbuf_1
Xwire4566 net4567 VGND VGND VPWR VPWR net4566 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_2_Left_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire3821 net3822 VGND VGND VPWR VPWR net3821 sky130_fd_sc_hd__buf_1
XFILLER_0_102_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24088_ _03948_ _03949_ VGND VGND VPWR VPWR _03951_ sky130_fd_sc_hd__or2_1
Xwire3832 net3833 VGND VGND VPWR VPWR net3832 sky130_fd_sc_hd__clkbuf_1
Xwire3843 net3844 VGND VGND VPWR VPWR net3843 sky130_fd_sc_hd__buf_1
Xwire3854 _12264_ VGND VGND VPWR VPWR net3854 sky130_fd_sc_hd__buf_1
Xwire4599 net4594 VGND VGND VPWR VPWR net4599 sky130_fd_sc_hd__buf_1
X_15930_ _07890_ _07907_ _07998_ VGND VGND VPWR VPWR _07999_ sky130_fd_sc_hd__o21ai_2
X_23039_ net5113 net4623 VGND VGND VPWR VPWR _02909_ sky130_fd_sc_hd__nand2_1
Xwire3876 _11035_ VGND VGND VPWR VPWR net3876 sky130_fd_sc_hd__clkbuf_1
Xwire3898 _10837_ VGND VGND VPWR VPWR net3898 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15861_ _07929_ net2671 _07837_ VGND VGND VPWR VPWR _07930_ sky130_fd_sc_hd__o21a_1
XFILLER_0_64_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17600_ net4006 svm0.tB\[7\] _09480_ VGND VGND VPWR VPWR _09481_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_157_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14812_ net3625 net7169 _06802_ net2855 VGND VGND VPWR VPWR _06923_ sky130_fd_sc_hd__o211a_1
X_18580_ net7044 _10423_ _10427_ VGND VGND VPWR VPWR _10428_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15792_ net1097 _07773_ _07861_ VGND VGND VPWR VPWR _07862_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17531_ net6694 net6742 svm0.delta\[14\] net6686 _09405_ VGND VGND VPWR VPWR _09414_
+ sky130_fd_sc_hd__o221a_1
X_14743_ net7453 _06876_ net2858 VGND VGND VPWR VPWR _06877_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17462_ net3273 _09355_ net6661 VGND VGND VPWR VPWR _09356_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14674_ net2865 VGND VGND VPWR VPWR _06825_ sky130_fd_sc_hd__buf_1
XFILLER_0_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19201_ net6207 net6141 net6244 VGND VGND VPWR VPWR _11038_ sky130_fd_sc_hd__and3_1
X_16413_ _08466_ _08474_ VGND VGND VPWR VPWR _08475_ sky130_fd_sc_hd__xor2_1
XFILLER_0_183_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13625_ _05888_ _05894_ VGND VGND VPWR VPWR _05895_ sky130_fd_sc_hd__xnor2_1
X_17393_ svm0.delta\[6\] _09296_ VGND VGND VPWR VPWR _09300_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19132_ _10862_ _10966_ _10908_ _10907_ VGND VGND VPWR VPWR _10969_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16344_ _08405_ _08406_ VGND VGND VPWR VPWR _08407_ sky130_fd_sc_hd__and2b_1
X_13556_ _05825_ _05826_ VGND VGND VPWR VPWR _05827_ sky130_fd_sc_hd__xor2_1
Xfanout7053 net7073 VGND VGND VPWR VPWR net7053 sky130_fd_sc_hd__buf_1
XFILLER_0_13_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19063_ _10898_ net2525 VGND VGND VPWR VPWR _10900_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout7086 net7102 VGND VGND VPWR VPWR net7086 sky130_fd_sc_hd__buf_1
Xfanout6341 net6345 VGND VGND VPWR VPWR net6341 sky130_fd_sc_hd__buf_1
X_16275_ _08333_ _08338_ VGND VGND VPWR VPWR _08339_ sky130_fd_sc_hd__xnor2_2
X_13487_ _05729_ _05759_ VGND VGND VPWR VPWR _05760_ sky130_fd_sc_hd__xor2_1
X_18014_ net7118 _09808_ _09862_ _09863_ _09864_ VGND VGND VPWR VPWR _09865_ sky130_fd_sc_hd__o221ai_1
Xwire7170 net7171 VGND VGND VPWR VPWR net7170 sky130_fd_sc_hd__buf_1
X_15226_ _07292_ _07296_ VGND VGND VPWR VPWR _07300_ sky130_fd_sc_hd__xor2_1
Xwire7181 matmul0.cos\[2\] VGND VGND VPWR VPWR net7181 sky130_fd_sc_hd__buf_1
XFILLER_0_125_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7192 net7193 VGND VGND VPWR VPWR net7192 sky130_fd_sc_hd__buf_1
XFILLER_0_124_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5673 net5681 VGND VGND VPWR VPWR net5673 sky130_fd_sc_hd__buf_1
Xwire6480 net6479 VGND VGND VPWR VPWR net6480 sky130_fd_sc_hd__buf_1
X_15157_ net3451 _07125_ VGND VGND VPWR VPWR _07231_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14108_ _06325_ _06329_ _06330_ VGND VGND VPWR VPWR _06370_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_129_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5790 net5791 VGND VGND VPWR VPWR net5790 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19965_ net6174 _11791_ _11795_ VGND VGND VPWR VPWR _11796_ sky130_fd_sc_hd__a21oi_1
X_15088_ _07094_ net1895 _07084_ VGND VGND VPWR VPWR _07162_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14039_ _06299_ _06302_ VGND VGND VPWR VPWR _06303_ sky130_fd_sc_hd__xnor2_2
X_18916_ net6814 _10755_ VGND VGND VPWR VPWR _10756_ sky130_fd_sc_hd__nand2_1
X_19896_ _11715_ _11727_ VGND VGND VPWR VPWR _11729_ sky130_fd_sc_hd__nand2_1
X_18847_ net6781 _10688_ _10689_ _10687_ VGND VGND VPWR VPWR _10690_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_98_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18778_ _10618_ _10619_ _10620_ _10621_ net421 _10561_ VGND VGND VPWR VPWR _10622_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17729_ net6502 _09587_ VGND VGND VPWR VPWR _00431_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20740_ net5557 net5823 VGND VGND VPWR VPWR _12511_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20671_ _12445_ _12447_ VGND VGND VPWR VPWR _12448_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22410_ _02380_ VGND VGND VPWR VPWR _02412_ sky130_fd_sc_hd__inv_2
X_23390_ _03256_ _03258_ VGND VGND VPWR VPWR _03260_ sky130_fd_sc_hd__nand2_1
XFILLER_0_161_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3829 _00960_ VGND VGND VPWR VPWR net3829 sky130_fd_sc_hd__buf_1
XFILLER_0_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22341_ net3778 _02343_ VGND VGND VPWR VPWR _02344_ sky130_fd_sc_hd__nor2_2
XFILLER_0_115_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22272_ _02095_ _02114_ _02170_ _02275_ VGND VGND VPWR VPWR _02276_ sky130_fd_sc_hd__a31o_1
X_25060_ net4430 net1995 _04807_ VGND VGND VPWR VPWR _04809_ sky130_fd_sc_hd__nor3_1
XFILLER_0_103_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24011_ net5048 net5027 net4500 VGND VGND VPWR VPWR _03874_ sky130_fd_sc_hd__and3_1
X_21223_ _01027_ _01234_ VGND VGND VPWR VPWR _01239_ sky130_fd_sc_hd__and2_1
Xhold120 cordic0.sin\[13\] VGND VGND VPWR VPWR net9073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 svm0.vC\[14\] VGND VGND VPWR VPWR net9084 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 svm0.vC\[2\] VGND VGND VPWR VPWR net9095 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 pid_d.prev_error\[3\] VGND VGND VPWR VPWR net9106 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3106 net3107 VGND VGND VPWR VPWR net3106 sky130_fd_sc_hd__clkbuf_1
X_21154_ net5628 net5912 VGND VGND VPWR VPWR _01170_ sky130_fd_sc_hd__nand2_1
Xwire3117 net3118 VGND VGND VPWR VPWR net3117 sky130_fd_sc_hd__clkbuf_1
Xhold164 pid_d.prev_error\[6\] VGND VGND VPWR VPWR net9117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 matmul0.matmul_stage_inst.c\[7\] VGND VGND VPWR VPWR net9128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 pid_q.prev_error\[4\] VGND VGND VPWR VPWR net9139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 matmul0.state\[0\] VGND VGND VPWR VPWR net9150 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3139 net3140 VGND VGND VPWR VPWR net3139 sky130_fd_sc_hd__clkbuf_1
Xwire2405 _04130_ VGND VGND VPWR VPWR net2405 sky130_fd_sc_hd__buf_1
X_20105_ _11906_ _11904_ _11907_ VGND VGND VPWR VPWR _11933_ sky130_fd_sc_hd__a21o_1
XFILLER_0_186_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2416 _03480_ VGND VGND VPWR VPWR net2416 sky130_fd_sc_hd__buf_1
XFILLER_0_10_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2427 _03271_ VGND VGND VPWR VPWR net2427 sky130_fd_sc_hd__buf_1
XFILLER_0_42_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21085_ net2075 net2074 net2480 VGND VGND VPWR VPWR _01101_ sky130_fd_sc_hd__a21oi_1
Xwire2438 _02660_ VGND VGND VPWR VPWR net2438 sky130_fd_sc_hd__clkbuf_1
Xwire1704 net1705 VGND VGND VPWR VPWR net1704 sky130_fd_sc_hd__buf_1
Xwire2449 net2450 VGND VGND VPWR VPWR net2449 sky130_fd_sc_hd__clkbuf_1
X_24913_ pid_q.ki\[0\] _04694_ _04702_ VGND VGND VPWR VPWR _04703_ sky130_fd_sc_hd__mux2_1
X_20036_ net3290 net2494 VGND VGND VPWR VPWR _11866_ sky130_fd_sc_hd__xnor2_1
Xwire1726 _01465_ VGND VGND VPWR VPWR net1726 sky130_fd_sc_hd__buf_1
X_25893_ clknet_leaf_14_clk _00766_ net8620 VGND VGND VPWR VPWR pid_q.kp\[5\] sky130_fd_sc_hd__dfrtp_1
Xwire1737 _00832_ VGND VGND VPWR VPWR net1737 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_137_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1748 _11644_ VGND VGND VPWR VPWR net1748 sky130_fd_sc_hd__clkbuf_1
Xwire1759 _10848_ VGND VGND VPWR VPWR net1759 sky130_fd_sc_hd__clkbuf_1
X_24844_ net7485 net455 _04257_ VGND VGND VPWR VPWR _04655_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24775_ _04602_ VGND VGND VPWR VPWR _04603_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21987_ net2477 net1046 _01994_ VGND VGND VPWR VPWR _01995_ sky130_fd_sc_hd__a21oi_1
X_23726_ _03590_ _03591_ VGND VGND VPWR VPWR _03592_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20938_ _00953_ _00941_ VGND VGND VPWR VPWR _00954_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23657_ _03516_ _03523_ VGND VGND VPWR VPWR _03524_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20869_ net5627 net5613 net5775 net5792 VGND VGND VPWR VPWR _00885_ sky130_fd_sc_hd__and4_1
XFILLER_0_187_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13410_ _05653_ _05682_ _05570_ _05652_ VGND VGND VPWR VPWR _05683_ sky130_fd_sc_hd__a2bb2o_1
X_22608_ pid_d.curr_error\[10\] net941 net3088 VGND VGND VPWR VPWR _02582_ sky130_fd_sc_hd__mux2_1
X_14390_ _06595_ matmul0.b_in\[0\] net900 VGND VGND VPWR VPWR _06596_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23588_ net4795 VGND VGND VPWR VPWR _03456_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13341_ _05520_ _05522_ VGND VGND VPWR VPWR _05614_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25327_ clknet_leaf_80_clk _00210_ net8491 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.f\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_22539_ pid_d.curr_error\[7\] net2381 net2048 VGND VGND VPWR VPWR _02532_ sky130_fd_sc_hd__and3_1
XFILLER_0_180_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16060_ _08118_ _08126_ VGND VGND VPWR VPWR _08127_ sky130_fd_sc_hd__xnor2_1
X_13272_ _05541_ _05542_ _05544_ VGND VGND VPWR VPWR _05545_ sky130_fd_sc_hd__a21oi_1
X_25258_ clknet_leaf_71_clk _00141_ net8458 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.b\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5031 net5032 VGND VGND VPWR VPWR net5031 sky130_fd_sc_hd__clkbuf_1
X_15011_ net3582 net3580 net4153 net4148 VGND VGND VPWR VPWR _07085_ sky130_fd_sc_hd__o22a_1
Xwire5042 net5036 VGND VGND VPWR VPWR net5042 sky130_fd_sc_hd__buf_1
X_24209_ _03983_ _03992_ _03991_ VGND VGND VPWR VPWR _04070_ sky130_fd_sc_hd__a21oi_1
Xwire5053 net5054 VGND VGND VPWR VPWR net5053 sky130_fd_sc_hd__buf_1
X_25189_ clknet_leaf_58_clk _00078_ net8720 VGND VGND VPWR VPWR matmul0.a_in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire5064 net5065 VGND VGND VPWR VPWR net5064 sky130_fd_sc_hd__buf_1
XFILLER_0_20_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5075 net5076 VGND VGND VPWR VPWR net5075 sky130_fd_sc_hd__buf_1
Xwire4330 net4324 VGND VGND VPWR VPWR net4330 sky130_fd_sc_hd__clkbuf_1
Xwire4341 net4342 VGND VGND VPWR VPWR net4341 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5097 net5098 VGND VGND VPWR VPWR net5097 sky130_fd_sc_hd__buf_1
XFILLER_0_20_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4374 net4375 VGND VGND VPWR VPWR net4374 sky130_fd_sc_hd__clkbuf_1
Xwire3640 net3641 VGND VGND VPWR VPWR net3640 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4385 net4383 VGND VGND VPWR VPWR net4385 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3651 net3652 VGND VGND VPWR VPWR net3651 sky130_fd_sc_hd__clkbuf_1
Xwire4396 pid_q.out\[15\] VGND VGND VPWR VPWR net4396 sky130_fd_sc_hd__clkbuf_1
X_19750_ net6171 net6198 net3150 net6097 VGND VGND VPWR VPWR _11585_ sky130_fd_sc_hd__o2bb2a_1
Xwire3662 net3663 VGND VGND VPWR VPWR net3662 sky130_fd_sc_hd__clkbuf_1
X_16962_ _08924_ VGND VGND VPWR VPWR _08925_ sky130_fd_sc_hd__buf_1
XFILLER_0_21_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3673 net3674 VGND VGND VPWR VPWR net3673 sky130_fd_sc_hd__buf_1
XFILLER_0_194_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3684 _05345_ VGND VGND VPWR VPWR net3684 sky130_fd_sc_hd__clkbuf_1
X_18701_ net3282 net2127 VGND VGND VPWR VPWR _10547_ sky130_fd_sc_hd__nor2_1
Xwire2950 net2951 VGND VGND VPWR VPWR net2950 sky130_fd_sc_hd__buf_1
Xwire3695 _04894_ VGND VGND VPWR VPWR net3695 sky130_fd_sc_hd__clkbuf_2
X_15913_ _07979_ net1094 VGND VGND VPWR VPWR _07982_ sky130_fd_sc_hd__xnor2_1
Xwire2961 net2962 VGND VGND VPWR VPWR net2961 sky130_fd_sc_hd__buf_1
X_19681_ net6200 _11512_ _11514_ _11515_ _11516_ VGND VGND VPWR VPWR _11517_ sky130_fd_sc_hd__o221a_1
X_16893_ net6370 VGND VGND VPWR VPWR _08857_ sky130_fd_sc_hd__inv_2
Xwire2972 _04963_ VGND VGND VPWR VPWR net2972 sky130_fd_sc_hd__buf_1
Xwire2983 net2984 VGND VGND VPWR VPWR net2983 sky130_fd_sc_hd__buf_1
Xwire2994 net2995 VGND VGND VPWR VPWR net2994 sky130_fd_sc_hd__clkbuf_2
X_15844_ _07909_ _07913_ VGND VGND VPWR VPWR _07914_ sky130_fd_sc_hd__xnor2_1
X_18632_ net6829 net6862 VGND VGND VPWR VPWR _10479_ sky130_fd_sc_hd__nand2_1
XFILLER_0_188_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15775_ _07837_ _07844_ VGND VGND VPWR VPWR _07845_ sky130_fd_sc_hd__xor2_1
X_18563_ _10331_ net765 _10410_ VGND VGND VPWR VPWR _10411_ sky130_fd_sc_hd__o21a_1
X_12987_ _05256_ _05259_ VGND VGND VPWR VPWR _05260_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_24_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17514_ _09315_ _09395_ _09399_ VGND VGND VPWR VPWR _09400_ sky130_fd_sc_hd__a21o_1
X_14726_ net9120 _06820_ net890 VGND VGND VPWR VPWR _00150_ sky130_fd_sc_hd__a21bo_1
X_18494_ net1771 net489 net1203 net9027 VGND VGND VPWR VPWR _00440_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17445_ net6741 net7376 net6744 net6738 VGND VGND VPWR VPWR _09341_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14657_ net7439 net7169 net2875 VGND VGND VPWR VPWR _06813_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13608_ _05874_ _05877_ VGND VGND VPWR VPWR _05878_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17376_ _09281_ _09282_ _09285_ net2567 VGND VGND VPWR VPWR _00378_ sky130_fd_sc_hd__a2bb2o_1
X_14588_ _06761_ _06762_ VGND VGND VPWR VPWR _06763_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19115_ _10949_ _10950_ _10940_ VGND VGND VPWR VPWR _10952_ sky130_fd_sc_hd__a21o_1
X_16327_ _08388_ _08389_ VGND VGND VPWR VPWR _08390_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13539_ net7686 net2321 net2317 VGND VGND VPWR VPWR _05810_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19046_ net6245 net3896 _10881_ _10882_ VGND VGND VPWR VPWR _10883_ sky130_fd_sc_hd__a211o_1
X_16258_ _08320_ _08321_ VGND VGND VPWR VPWR _08322_ sky130_fd_sc_hd__xnor2_1
Xfanout6182 net6185 VGND VGND VPWR VPWR net6182 sky130_fd_sc_hd__buf_1
XFILLER_0_3_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15209_ _07281_ _07282_ VGND VGND VPWR VPWR _07283_ sky130_fd_sc_hd__xnor2_1
X_16189_ net2691 net2731 net2645 _08253_ VGND VGND VPWR VPWR _08254_ sky130_fd_sc_hd__or4_1
XFILLER_0_49_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19948_ _11772_ _11779_ VGND VGND VPWR VPWR _11780_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19879_ _11674_ _11711_ VGND VGND VPWR VPWR _11712_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21910_ _01916_ _01821_ _01917_ VGND VGND VPWR VPWR _01918_ sky130_fd_sc_hd__o21a_1
XFILLER_0_65_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22890_ _02784_ VGND VGND VPWR VPWR _00640_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21841_ _01846_ _01849_ VGND VGND VPWR VPWR _01850_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_179_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24560_ _04415_ _04343_ _04345_ VGND VGND VPWR VPWR _04416_ sky130_fd_sc_hd__a21oi_1
X_21772_ net5812 net5406 VGND VGND VPWR VPWR _01782_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23511_ net1166 net938 _03299_ VGND VGND VPWR VPWR _03380_ sky130_fd_sc_hd__o21a_1
X_20723_ net1817 _12484_ _12491_ _12494_ VGND VGND VPWR VPWR _12495_ sky130_fd_sc_hd__nor4_1
X_24491_ _03197_ net4499 net3756 VGND VGND VPWR VPWR _04348_ sky130_fd_sc_hd__a21o_1
XFILLER_0_81_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23442_ pid_q.prev_error\[0\] pid_q.curr_error\[0\] VGND VGND VPWR VPWR _03312_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_163_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7906 net7907 VGND VGND VPWR VPWR net7906 sky130_fd_sc_hd__buf_1
X_20654_ net6133 _12421_ VGND VGND VPWR VPWR _12432_ sky130_fd_sc_hd__nand2_1
Xwire7917 net7914 VGND VGND VPWR VPWR net7917 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_74_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire308 net309 VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__clkbuf_1
Xwire319 _06276_ VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__buf_1
Xwire7928 net7929 VGND VGND VPWR VPWR net7928 sky130_fd_sc_hd__clkbuf_1
Xwire7939 net7940 VGND VGND VPWR VPWR net7939 sky130_fd_sc_hd__clkbuf_1
X_23373_ net4700 net4914 VGND VGND VPWR VPWR _03243_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20585_ _08991_ _12367_ VGND VGND VPWR VPWR _12368_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2914 _06516_ VGND VGND VPWR VPWR net2914 sky130_fd_sc_hd__dlymetal6s2s_1
X_25112_ net4392 net2392 net1992 net9206 VGND VGND VPWR VPWR _00793_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22324_ _04887_ net297 VGND VGND VPWR VPWR _02328_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25043_ net3738 _04790_ pid_q.out\[6\] VGND VGND VPWR VPWR _04794_ sky130_fd_sc_hd__o21ba_1
X_22255_ net4364 _02258_ _02259_ VGND VGND VPWR VPWR _02260_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21206_ net808 _01078_ _01221_ VGND VGND VPWR VPWR _01222_ sky130_fd_sc_hd__o21a_1
X_22186_ net859 _02159_ VGND VGND VPWR VPWR _02191_ sky130_fd_sc_hd__or2b_1
Xwire2202 net2203 VGND VGND VPWR VPWR net2202 sky130_fd_sc_hd__buf_1
XFILLER_0_100_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21137_ _01149_ _01152_ VGND VGND VPWR VPWR _01153_ sky130_fd_sc_hd__xnor2_1
Xwire2213 net2214 VGND VGND VPWR VPWR net2213 sky130_fd_sc_hd__clkbuf_1
Xwire2224 _07810_ VGND VGND VPWR VPWR net2224 sky130_fd_sc_hd__buf_1
Xwire1501 _08905_ VGND VGND VPWR VPWR net1501 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2246 net2247 VGND VGND VPWR VPWR net2246 sky130_fd_sc_hd__buf_1
X_21068_ net5835 net5871 _12556_ VGND VGND VPWR VPWR _01084_ sky130_fd_sc_hd__and3_1
Xwire2257 net2258 VGND VGND VPWR VPWR net2257 sky130_fd_sc_hd__clkbuf_1
Xwire1512 _08175_ VGND VGND VPWR VPWR net1512 sky130_fd_sc_hd__buf_1
Xwire1523 net1524 VGND VGND VPWR VPWR net1523 sky130_fd_sc_hd__buf_1
Xwire2268 net2269 VGND VGND VPWR VPWR net2268 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_92_Left_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2279 net2280 VGND VGND VPWR VPWR net2279 sky130_fd_sc_hd__clkbuf_1
Xwire1534 _07771_ VGND VGND VPWR VPWR net1534 sky130_fd_sc_hd__clkbuf_1
X_12910_ net1143 _05182_ VGND VGND VPWR VPWR _05183_ sky130_fd_sc_hd__xnor2_1
Xwire1545 net1546 VGND VGND VPWR VPWR net1545 sky130_fd_sc_hd__buf_1
X_20019_ net1406 net2093 _11808_ VGND VGND VPWR VPWR _11849_ sky130_fd_sc_hd__o21a_1
Xwire1556 net1557 VGND VGND VPWR VPWR net1556 sky130_fd_sc_hd__buf_1
X_25876_ clknet_leaf_15_clk _00749_ net8618 VGND VGND VPWR VPWR pid_q.ki\[4\] sky130_fd_sc_hd__dfrtp_1
X_13890_ _06142_ _06153_ _06155_ net449 VGND VGND VPWR VPWR _06156_ sky130_fd_sc_hd__a2bb2o_1
Xwire1567 _05764_ VGND VGND VPWR VPWR net1567 sky130_fd_sc_hd__buf_1
Xwire1578 net1579 VGND VGND VPWR VPWR net1578 sky130_fd_sc_hd__buf_1
Xwire1589 net1591 VGND VGND VPWR VPWR net1589 sky130_fd_sc_hd__buf_1
XFILLER_0_69_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24827_ net5091 _04642_ net2000 net926 VGND VGND VPWR VPWR _00715_ sky130_fd_sc_hd__a22o_1
X_12841_ _05108_ _05109_ _05112_ _05113_ VGND VGND VPWR VPWR _05114_ sky130_fd_sc_hd__o211ai_1
X_15560_ _07541_ _07502_ _07632_ VGND VGND VPWR VPWR _07633_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24758_ _04586_ _04587_ VGND VGND VPWR VPWR _04588_ sky130_fd_sc_hd__and2_1
X_12772_ _04927_ _04933_ _05044_ VGND VGND VPWR VPWR _05045_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14511_ net3032 _06691_ VGND VGND VPWR VPWR _06692_ sky130_fd_sc_hd__nand2_1
XFILLER_0_178_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23709_ net7527 _03485_ net467 net7468 net1663 VGND VGND VPWR VPWR _03576_ sky130_fd_sc_hd__a221o_1
XFILLER_0_83_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15491_ _07402_ _07544_ VGND VGND VPWR VPWR _07564_ sky130_fd_sc_hd__or2_1
Xmax_length6263 net6261 VGND VGND VPWR VPWR net6263 sky130_fd_sc_hd__clkbuf_1
X_24689_ net7475 net3269 net8875 VGND VGND VPWR VPWR _04527_ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length5540 net5532 VGND VGND VPWR VPWR net5540 sky130_fd_sc_hd__buf_1
X_17230_ net3280 _09165_ VGND VGND VPWR VPWR _09178_ sky130_fd_sc_hd__or2_1
X_14442_ _06635_ matmul0.b_in\[12\] net895 VGND VGND VPWR VPWR _06636_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17161_ net822 VGND VGND VPWR VPWR _09114_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire820 net821 VGND VGND VPWR VPWR net820 sky130_fd_sc_hd__clkbuf_1
X_14373_ net7225 net1297 net2894 net5333 _06582_ VGND VGND VPWR VPWR _06583_ sky130_fd_sc_hd__a221o_1
XFILLER_0_182_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire842 _05631_ VGND VGND VPWR VPWR net842 sky130_fd_sc_hd__buf_1
XFILLER_0_88_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16112_ net3449 net2719 net3499 VGND VGND VPWR VPWR _08178_ sky130_fd_sc_hd__a21o_1
Xwire853 _04100_ VGND VGND VPWR VPWR net853 sky130_fd_sc_hd__clkbuf_1
X_13324_ net7774 _04960_ _05507_ VGND VGND VPWR VPWR _05597_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire864 _12218_ VGND VGND VPWR VPWR net864 sky130_fd_sc_hd__clkbuf_1
X_17092_ net6981 _09048_ _09049_ _09047_ VGND VGND VPWR VPWR _00331_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire875 _10269_ VGND VGND VPWR VPWR net875 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire886 _07962_ VGND VGND VPWR VPWR net886 sky130_fd_sc_hd__clkbuf_1
Xwire897 net898 VGND VGND VPWR VPWR net897 sky130_fd_sc_hd__buf_1
X_16043_ net2640 _08109_ VGND VGND VPWR VPWR _08110_ sky130_fd_sc_hd__nand2_1
X_13255_ net7923 _05527_ VGND VGND VPWR VPWR _05528_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_108_Right_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13186_ net7689 net2350 net2346 VGND VGND VPWR VPWR _05459_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4160 net4161 VGND VGND VPWR VPWR net4160 sky130_fd_sc_hd__buf_1
X_19802_ net6170 net2104 VGND VGND VPWR VPWR _11636_ sky130_fd_sc_hd__xnor2_1
Xwire4182 net4183 VGND VGND VPWR VPWR net4182 sky130_fd_sc_hd__buf_1
X_17994_ _09843_ VGND VGND VPWR VPWR _09845_ sky130_fd_sc_hd__inv_2
Xwire3470 _07152_ VGND VGND VPWR VPWR net3470 sky130_fd_sc_hd__clkbuf_1
X_19733_ net6030 _11501_ _11566_ _11567_ VGND VGND VPWR VPWR _11568_ sky130_fd_sc_hd__o211a_1
Xwire3481 net3482 VGND VGND VPWR VPWR net3481 sky130_fd_sc_hd__dlymetal6s2s_1
X_16945_ net4241 VGND VGND VPWR VPWR _08909_ sky130_fd_sc_hd__buf_1
Xwire3492 net3493 VGND VGND VPWR VPWR net3492 sky130_fd_sc_hd__buf_1
X_19664_ net2502 _11499_ VGND VGND VPWR VPWR _11500_ sky130_fd_sc_hd__xnor2_2
Xwire2791 net2792 VGND VGND VPWR VPWR net2791 sky130_fd_sc_hd__clkbuf_2
X_16876_ net7134 _08839_ _08840_ net1828 VGND VGND VPWR VPWR _00324_ sky130_fd_sc_hd__a22o_1
X_18615_ _10439_ VGND VGND VPWR VPWR _10462_ sky130_fd_sc_hd__inv_2
X_15827_ net2799 net2216 net2225 VGND VGND VPWR VPWR _07897_ sky130_fd_sc_hd__or3_1
XFILLER_0_17_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19595_ _11431_ net2106 VGND VGND VPWR VPWR _11432_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15758_ _07737_ _07828_ VGND VGND VPWR VPWR _07829_ sky130_fd_sc_hd__xor2_1
X_18546_ _10328_ _10346_ _10394_ VGND VGND VPWR VPWR _10395_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_158_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14709_ matmul0.sin\[10\] _06851_ VGND VGND VPWR VPWR _06852_ sky130_fd_sc_hd__xnor2_1
X_15689_ net3550 _07759_ VGND VGND VPWR VPWR _07760_ sky130_fd_sc_hd__nor2_1
X_18477_ _10308_ _10326_ VGND VGND VPWR VPWR _10327_ sky130_fd_sc_hd__xnor2_1
X_17428_ _09326_ _09327_ svm0.delta\[14\] VGND VGND VPWR VPWR _09328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17359_ net3277 VGND VGND VPWR VPWR _09272_ sky130_fd_sc_hd__buf_1
XFILLER_0_67_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20370_ _12166_ _12169_ VGND VGND VPWR VPWR _12170_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_152_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19029_ _10817_ _10806_ _10807_ _10833_ _10865_ VGND VGND VPWR VPWR _10866_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_28_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22040_ _01942_ _01943_ _02046_ VGND VGND VPWR VPWR _02047_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23991_ pid_q.prev_error\[6\] pid_q.curr_error\[6\] VGND VGND VPWR VPWR _03855_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_177_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25730_ clknet_leaf_8_clk _00603_ net8554 VGND VGND VPWR VPWR pid_d.ki\[4\] sky130_fd_sc_hd__dfrtp_1
X_22942_ pid_d.curr_int\[14\] _02830_ VGND VGND VPWR VPWR _02831_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_183_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25661_ clknet_leaf_24_clk _00534_ net8584 VGND VGND VPWR VPWR pid_d.curr_int\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22873_ _01819_ _02762_ net5363 VGND VGND VPWR VPWR _02769_ sky130_fd_sc_hd__o21ba_1
X_24612_ _04423_ _04460_ _04462_ _04466_ VGND VGND VPWR VPWR _04467_ sky130_fd_sc_hd__o211a_1
X_21824_ net5686 net5539 VGND VGND VPWR VPWR _01833_ sky130_fd_sc_hd__nand2_1
XFILLER_0_195_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25592_ clknet_leaf_91_clk _00465_ net8428 VGND VGND VPWR VPWR cordic0.cos\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_24543_ _04373_ _04374_ _04398_ _04264_ VGND VGND VPWR VPWR _04399_ sky130_fd_sc_hd__a22o_1
X_21755_ net5785 net5461 VGND VGND VPWR VPWR _01765_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8404 net8401 VGND VGND VPWR VPWR net8404 sky130_fd_sc_hd__clkbuf_2
Xwire8415 net8416 VGND VGND VPWR VPWR net8415 sky130_fd_sc_hd__clkbuf_1
X_20706_ _12463_ _12464_ _12473_ _08993_ VGND VGND VPWR VPWR _12479_ sky130_fd_sc_hd__o31a_1
X_24474_ net5173 pid_q.prev_int\[13\] VGND VGND VPWR VPWR _04331_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21686_ _01695_ _01696_ VGND VGND VPWR VPWR _01697_ sky130_fd_sc_hd__or2b_1
XFILLER_0_53_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8437 net8435 VGND VGND VPWR VPWR net8437 sky130_fd_sc_hd__buf_1
XFILLER_0_81_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7703 net7704 VGND VGND VPWR VPWR net7703 sky130_fd_sc_hd__buf_1
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8448 net8449 VGND VGND VPWR VPWR net8448 sky130_fd_sc_hd__buf_1
XFILLER_0_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7714 net7716 VGND VGND VPWR VPWR net7714 sky130_fd_sc_hd__buf_1
X_23425_ net1385 _03294_ VGND VGND VPWR VPWR _03295_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_163_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7725 net7726 VGND VGND VPWR VPWR net7725 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7736 net7737 VGND VGND VPWR VPWR net7736 sky130_fd_sc_hd__buf_1
XFILLER_0_11_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20637_ _12416_ VGND VGND VPWR VPWR _00510_ sky130_fd_sc_hd__clkbuf_1
Xwire7747 net7745 VGND VGND VPWR VPWR net7747 sky130_fd_sc_hd__buf_1
XFILLER_0_184_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7758 net7759 VGND VGND VPWR VPWR net7758 sky130_fd_sc_hd__buf_1
XFILLER_0_117_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23356_ _03223_ net2428 VGND VGND VPWR VPWR _03226_ sky130_fd_sc_hd__xnor2_1
Xmax_length3467 net3468 VGND VGND VPWR VPWR net3467 sky130_fd_sc_hd__buf_1
XFILLER_0_6_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20568_ net3325 net3847 _12351_ VGND VGND VPWR VPWR _12352_ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22307_ net1704 net1703 _02310_ VGND VGND VPWR VPWR _02311_ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23287_ _03149_ _03156_ VGND VGND VPWR VPWR _03157_ sky130_fd_sc_hd__xnor2_1
Xmax_length2777 net2778 VGND VGND VPWR VPWR net2777 sky130_fd_sc_hd__clkbuf_1
X_20499_ _12284_ _12285_ _12286_ net6350 VGND VGND VPWR VPWR _00502_ sky130_fd_sc_hd__o22a_1
X_25026_ net7512 net2396 VGND VGND VPWR VPWR _04779_ sky130_fd_sc_hd__and2_1
X_13040_ net790 _05185_ _05184_ VGND VGND VPWR VPWR _05313_ sky130_fd_sc_hd__nand3b_1
X_22238_ _02160_ _02190_ net2062 VGND VGND VPWR VPWR _02243_ sky130_fd_sc_hd__o21a_1
X_22169_ _02174_ _02102_ pid_d.prev_error\[9\] VGND VGND VPWR VPWR _02175_ sky130_fd_sc_hd__o21ba_1
Xwire2010 _04583_ VGND VGND VPWR VPWR net2010 sky130_fd_sc_hd__clkbuf_1
Xwire2021 _04076_ VGND VGND VPWR VPWR net2021 sky130_fd_sc_hd__buf_1
XFILLER_0_79_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2032 _02715_ VGND VGND VPWR VPWR net2032 sky130_fd_sc_hd__clkbuf_1
X_14991_ net2850 net3525 _07064_ VGND VGND VPWR VPWR _07065_ sky130_fd_sc_hd__a21oi_1
Xwire2054 _02209_ VGND VGND VPWR VPWR net2054 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1320 _05611_ VGND VGND VPWR VPWR net1320 sky130_fd_sc_hd__buf_1
Xwire2065 net2066 VGND VGND VPWR VPWR net2065 sky130_fd_sc_hd__buf_1
Xwire1331 net1332 VGND VGND VPWR VPWR net1331 sky130_fd_sc_hd__buf_1
Xwire2076 _00974_ VGND VGND VPWR VPWR net2076 sky130_fd_sc_hd__buf_1
X_13942_ _06112_ _06206_ _06207_ VGND VGND VPWR VPWR _06208_ sky130_fd_sc_hd__o21ai_2
Xwire1342 _05012_ VGND VGND VPWR VPWR net1342 sky130_fd_sc_hd__buf_1
Xwire2087 net2088 VGND VGND VPWR VPWR net2087 sky130_fd_sc_hd__buf_1
X_16730_ _08753_ VGND VGND VPWR VPWR _00265_ sky130_fd_sc_hd__clkbuf_1
X_25928_ clknet_leaf_2_clk _00801_ net8574 VGND VGND VPWR VPWR pid_d.prev_int\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1353 net1354 VGND VGND VPWR VPWR net1353 sky130_fd_sc_hd__buf_1
Xwire2098 _11692_ VGND VGND VPWR VPWR net2098 sky130_fd_sc_hd__clkbuf_1
Xwire1364 _04647_ VGND VGND VPWR VPWR net1364 sky130_fd_sc_hd__clkbuf_1
Xwire1386 net1387 VGND VGND VPWR VPWR net1386 sky130_fd_sc_hd__clkbuf_1
X_16661_ _08694_ _08695_ VGND VGND VPWR VPWR _08696_ sky130_fd_sc_hd__xnor2_1
X_25859_ clknet_leaf_16_clk _00732_ net8619 VGND VGND VPWR VPWR pid_q.mult0.a\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13873_ net7807 net1568 net996 _06139_ VGND VGND VPWR VPWR _06140_ sky130_fd_sc_hd__a31o_1
Xwire1397 _12378_ VGND VGND VPWR VPWR net1397 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18400_ _10155_ net1775 VGND VGND VPWR VPWR _10251_ sky130_fd_sc_hd__or2_1
X_15612_ net4069 VGND VGND VPWR VPWR _07684_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12824_ _05095_ _05096_ VGND VGND VPWR VPWR _05097_ sky130_fd_sc_hd__xnor2_1
X_19380_ net2509 _11209_ _11216_ _11208_ net2518 VGND VGND VPWR VPWR _11217_ sky130_fd_sc_hd__o311a_1
X_16592_ _08643_ VGND VGND VPWR VPWR _00237_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15543_ _07614_ _07615_ VGND VGND VPWR VPWR _07616_ sky130_fd_sc_hd__xor2_1
X_18331_ _10093_ net2138 VGND VGND VPWR VPWR _10182_ sky130_fd_sc_hd__or2b_1
X_12755_ _04997_ _05027_ net1611 VGND VGND VPWR VPWR _05028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18262_ _10106_ _10107_ net2138 VGND VGND VPWR VPWR _10113_ sky130_fd_sc_hd__nand3_1
X_15474_ _07545_ _07547_ _07402_ VGND VGND VPWR VPWR _07548_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_155_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12686_ net2974 VGND VGND VPWR VPWR _04959_ sky130_fd_sc_hd__buf_1
XFILLER_0_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8887 net8890 VGND VGND VPWR VPWR net8887 sky130_fd_sc_hd__buf_1
X_17213_ _09160_ _09161_ VGND VGND VPWR VPWR _09162_ sky130_fd_sc_hd__and2_1
X_14425_ net5243 net1295 net2891 net4431 _06622_ VGND VGND VPWR VPWR _06623_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18193_ net3948 _09793_ _10043_ VGND VGND VPWR VPWR _10044_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_115_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17144_ _09097_ net3305 VGND VGND VPWR VPWR _09098_ sky130_fd_sc_hd__nor2_1
Xwire650 net651 VGND VGND VPWR VPWR net650 sky130_fd_sc_hd__clkbuf_1
X_14356_ net3647 VGND VGND VPWR VPWR _06569_ sky130_fd_sc_hd__buf_1
XFILLER_0_21_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire661 net662 VGND VGND VPWR VPWR net661 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_188_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire672 _08210_ VGND VGND VPWR VPWR net672 sky130_fd_sc_hd__dlymetal6s2s_1
X_13307_ net1572 net1945 VGND VGND VPWR VPWR _05580_ sky130_fd_sc_hd__xor2_1
Xwire683 _05337_ VGND VGND VPWR VPWR net683 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_97_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire694 net695 VGND VGND VPWR VPWR net694 sky130_fd_sc_hd__buf_1
X_17075_ net3313 net4040 VGND VGND VPWR VPWR _09033_ sky130_fd_sc_hd__nor2_1
X_14287_ net76 _06518_ _06519_ net7819 VGND VGND VPWR VPWR _00056_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16026_ _08014_ _08091_ _08092_ VGND VGND VPWR VPWR _08093_ sky130_fd_sc_hd__a21oi_1
X_13238_ _05451_ _05452_ _05510_ VGND VGND VPWR VPWR _05511_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_139_Left_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_196_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13169_ net7802 net3687 net2970 VGND VGND VPWR VPWR _05442_ sky130_fd_sc_hd__and3_1
XFILLER_0_137_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17977_ net2141 _09612_ net1780 VGND VGND VPWR VPWR _09828_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19716_ _11546_ _11551_ VGND VGND VPWR VPWR _11552_ sky130_fd_sc_hd__xnor2_1
X_16928_ net6418 _08891_ _08884_ VGND VGND VPWR VPWR _08892_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19647_ _11481_ _11483_ VGND VGND VPWR VPWR _11484_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16859_ net6525 VGND VGND VPWR VPWR _08824_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_148_Left_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19578_ _11327_ net1419 _11414_ VGND VGND VPWR VPWR _11415_ sky130_fd_sc_hd__o21a_1
XFILLER_0_153_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18529_ net1765 _10376_ VGND VGND VPWR VPWR _10378_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21540_ _01547_ net652 _01550_ _01551_ VGND VGND VPWR VPWR _01552_ sky130_fd_sc_hd__a31o_1
XFILLER_0_75_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21471_ net5864 net5429 VGND VGND VPWR VPWR _01484_ sky130_fd_sc_hd__nand2_1
Xwire6309 net6310 VGND VGND VPWR VPWR net6309 sky130_fd_sc_hd__buf_1
X_23210_ _03039_ _03079_ net5157 net5116 net3752 VGND VGND VPWR VPWR _03080_ sky130_fd_sc_hd__o2111a_1
X_20422_ _12215_ _12216_ _12217_ net6459 VGND VGND VPWR VPWR _12218_ sky130_fd_sc_hd__a31oi_1
X_24190_ _03976_ VGND VGND VPWR VPWR _04051_ sky130_fd_sc_hd__inv_2
Xwire5608 net5609 VGND VGND VPWR VPWR net5608 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23141_ net5084 net4697 VGND VGND VPWR VPWR _03011_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_157_Left_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20353_ net9168 _12153_ _12154_ VGND VGND VPWR VPWR _00488_ sky130_fd_sc_hd__a21bo_1
Xwire4907 net4908 VGND VGND VPWR VPWR net4907 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4918 net4919 VGND VGND VPWR VPWR net4918 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4929 net4930 VGND VGND VPWR VPWR net4929 sky130_fd_sc_hd__buf_1
X_23072_ net5041 net4634 VGND VGND VPWR VPWR _02942_ sky130_fd_sc_hd__nand2_1
X_20284_ net6499 net6468 VGND VGND VPWR VPWR _12090_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22023_ net5709 net5480 VGND VGND VPWR VPWR _02030_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold13 cordic0.sin\[3\] VGND VGND VPWR VPWR net8966 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 _00014_ VGND VGND VPWR VPWR net8977 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 pid_d.prev_error\[14\] VGND VGND VPWR VPWR net8988 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 pid_q.target\[9\] VGND VGND VPWR VPWR net8999 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold57 pid_q.target\[0\] VGND VGND VPWR VPWR net9010 sky130_fd_sc_hd__dlygate4sd3_1
X_23974_ _03734_ _03746_ _03736_ VGND VGND VPWR VPWR _03838_ sky130_fd_sc_hd__a21bo_1
Xhold68 matmul0.matmul_stage_inst.a\[11\] VGND VGND VPWR VPWR net9021 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 pid_q.prev_error\[12\] VGND VGND VPWR VPWR net9032 sky130_fd_sc_hd__dlygate4sd3_1
X_25713_ clknet_leaf_9_clk _00586_ net8552 VGND VGND VPWR VPWR pid_d.mult0.a\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_22925_ net5339 _02809_ _02815_ VGND VGND VPWR VPWR _02816_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_166_Left_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25644_ clknet_leaf_102_clk _00517_ net8367 VGND VGND VPWR VPWR cordic0.vec\[0\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_22856_ _02752_ _02753_ VGND VGND VPWR VPWR _02754_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21807_ net4385 _01740_ net473 net4319 net804 VGND VGND VPWR VPWR _01817_ sky130_fd_sc_hd__a221o_1
X_25575_ clknet_leaf_97_clk _00448_ net8398 VGND VGND VPWR VPWR cordic0.sin\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22787_ _02701_ VGND VGND VPWR VPWR _00620_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24526_ net7463 VGND VGND VPWR VPWR _04383_ sky130_fd_sc_hd__inv_2
Xwire8201 net8202 VGND VGND VPWR VPWR net8201 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21738_ _01660_ _01670_ _01747_ VGND VGND VPWR VPWR _01748_ sky130_fd_sc_hd__o21a_1
Xwire8212 net8213 VGND VGND VPWR VPWR net8212 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8223 net8224 VGND VGND VPWR VPWR net8223 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8234 net8235 VGND VGND VPWR VPWR net8234 sky130_fd_sc_hd__clkbuf_1
Xwire7500 net7496 VGND VGND VPWR VPWR net7500 sky130_fd_sc_hd__buf_1
Xwire8245 net8246 VGND VGND VPWR VPWR net8245 sky130_fd_sc_hd__clkbuf_1
Xwire7511 net7515 VGND VGND VPWR VPWR net7511 sky130_fd_sc_hd__buf_1
XFILLER_0_136_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24457_ _04313_ net928 VGND VGND VPWR VPWR _04315_ sky130_fd_sc_hd__or2b_2
Xwire8256 net8257 VGND VGND VPWR VPWR net8256 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7522 net7524 VGND VGND VPWR VPWR net7522 sky130_fd_sc_hd__buf_1
X_21669_ net5701 net5572 _01678_ _01679_ VGND VGND VPWR VPWR _01680_ sky130_fd_sc_hd__a31o_1
Xwire8267 net8268 VGND VGND VPWR VPWR net8267 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7533 net7534 VGND VGND VPWR VPWR net7533 sky130_fd_sc_hd__clkbuf_1
Xwire8278 net8279 VGND VGND VPWR VPWR net8278 sky130_fd_sc_hd__clkbuf_1
X_14210_ _06445_ _06468_ _06467_ VGND VGND VPWR VPWR _06469_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8289 net22 VGND VGND VPWR VPWR net8289 sky130_fd_sc_hd__clkbuf_1
Xwire7544 net7545 VGND VGND VPWR VPWR net7544 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_193_Right_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23408_ net2427 _03276_ VGND VGND VPWR VPWR _03278_ sky130_fd_sc_hd__nand2_1
Xwire7555 matmul0.b_in\[15\] VGND VGND VPWR VPWR net7555 sky130_fd_sc_hd__clkbuf_1
Xwire6810 net6811 VGND VGND VPWR VPWR net6810 sky130_fd_sc_hd__buf_1
X_15190_ net991 _07263_ VGND VGND VPWR VPWR _07264_ sky130_fd_sc_hd__xnor2_1
Xfanout6759 net6768 VGND VGND VPWR VPWR net6759 sky130_fd_sc_hd__buf_1
Xmax_length3253 net3254 VGND VGND VPWR VPWR net3253 sky130_fd_sc_hd__buf_1
Xwire6821 net6822 VGND VGND VPWR VPWR net6821 sky130_fd_sc_hd__buf_1
Xwire7566 matmul0.b_in\[9\] VGND VGND VPWR VPWR net7566 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_175_Left_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24388_ _04162_ _04164_ _04121_ VGND VGND VPWR VPWR _04247_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6832 net6833 VGND VGND VPWR VPWR net6832 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire7577 net7578 VGND VGND VPWR VPWR net7577 sky130_fd_sc_hd__clkbuf_1
Xwire7588 matmul0.a_in\[13\] VGND VGND VPWR VPWR net7588 sky130_fd_sc_hd__clkbuf_1
X_14141_ _06377_ _06392_ VGND VGND VPWR VPWR _06402_ sky130_fd_sc_hd__and2b_1
Xwire7599 matmul0.a_in\[9\] VGND VGND VPWR VPWR net7599 sky130_fd_sc_hd__clkbuf_1
Xmax_length3286 net3287 VGND VGND VPWR VPWR net3286 sky130_fd_sc_hd__buf_1
X_23339_ net5057 net4618 VGND VGND VPWR VPWR _03209_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6898 net6900 VGND VGND VPWR VPWR net6898 sky130_fd_sc_hd__clkbuf_1
X_14072_ _06117_ net1125 _06334_ net4249 VGND VGND VPWR VPWR _06335_ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13023_ net7878 net2966 net2305 VGND VGND VPWR VPWR _05296_ sky130_fd_sc_hd__and3_1
X_25009_ _04762_ _04763_ VGND VGND VPWR VPWR _04765_ sky130_fd_sc_hd__nand2_1
X_17900_ _09640_ _09750_ VGND VGND VPWR VPWR _09751_ sky130_fd_sc_hd__xnor2_2
X_18880_ _10680_ net1194 VGND VGND VPWR VPWR _10722_ sky130_fd_sc_hd__xnor2_1
X_17831_ net7060 net7027 VGND VGND VPWR VPWR _09682_ sky130_fd_sc_hd__nor2_1
X_17762_ net7103 net7121 VGND VGND VPWR VPWR _09613_ sky130_fd_sc_hd__or2b_1
XPHY_EDGE_ROW_184_Left_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14974_ net4178 _06998_ net4182 net4180 VGND VGND VPWR VPWR _07048_ sky130_fd_sc_hd__o22a_1
Xwire1150 net1151 VGND VGND VPWR VPWR net1150 sky130_fd_sc_hd__buf_1
Xwire1161 _03829_ VGND VGND VPWR VPWR net1161 sky130_fd_sc_hd__clkbuf_2
X_19501_ net6154 _11267_ _11336_ _11337_ VGND VGND VPWR VPWR _11338_ sky130_fd_sc_hd__o211a_1
Xwire1172 _01777_ VGND VGND VPWR VPWR net1172 sky130_fd_sc_hd__buf_1
XFILLER_0_92_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16713_ matmul0.matmul_stage_inst.mult1\[13\] VGND VGND VPWR VPWR _08740_ sky130_fd_sc_hd__inv_2
X_13925_ _06093_ _06094_ _06190_ VGND VGND VPWR VPWR _06191_ sky130_fd_sc_hd__a21oi_2
X_17693_ net9244 net2568 _09572_ net9048 net3384 VGND VGND VPWR VPWR _00409_ sky130_fd_sc_hd__a32o_1
Xwire1183 net1184 VGND VGND VPWR VPWR net1183 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_16_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1194 _10721_ VGND VGND VPWR VPWR net1194 sky130_fd_sc_hd__buf_1
X_19432_ _11035_ _11268_ VGND VGND VPWR VPWR _11269_ sky130_fd_sc_hd__xnor2_1
X_13856_ _06120_ _06122_ VGND VGND VPWR VPWR _06123_ sky130_fd_sc_hd__xnor2_1
X_16644_ _08679_ _08672_ _08674_ _08680_ VGND VGND VPWR VPWR _08681_ sky130_fd_sc_hd__a31o_1
XFILLER_0_190_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12807_ _04979_ _04997_ _04994_ VGND VGND VPWR VPWR _05080_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19363_ _11186_ _11196_ _11198_ _11199_ VGND VGND VPWR VPWR _11200_ sky130_fd_sc_hd__or4_1
X_13787_ _06053_ _06054_ VGND VGND VPWR VPWR _06055_ sky130_fd_sc_hd__xnor2_1
X_16575_ _08632_ _08633_ VGND VGND VPWR VPWR _08634_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18314_ _09026_ net7034 net7110 VGND VGND VPWR VPWR _10165_ sky130_fd_sc_hd__and3_1
X_12738_ net2358 net1980 VGND VGND VPWR VPWR _05011_ sky130_fd_sc_hd__and2_1
X_15526_ net2852 _07598_ _07518_ _07519_ VGND VGND VPWR VPWR _07599_ sky130_fd_sc_hd__a31o_1
X_19294_ net3173 _10986_ _10918_ VGND VGND VPWR VPWR _11131_ sky130_fd_sc_hd__or3_1
XFILLER_0_45_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8673 net8697 VGND VGND VPWR VPWR net8673 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_38_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout8684 net8701 VGND VGND VPWR VPWR net8684 sky130_fd_sc_hd__clkbuf_2
X_15457_ _07526_ _07530_ VGND VGND VPWR VPWR _07531_ sky130_fd_sc_hd__xnor2_1
X_18245_ _10039_ _10040_ net6911 VGND VGND VPWR VPWR _10096_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_193_Left_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12669_ net7836 net1974 net1971 VGND VGND VPWR VPWR _04942_ sky130_fd_sc_hd__and3_1
XFILLER_0_143_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14408_ net8146 net3633 VGND VGND VPWR VPWR _06610_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_160_Right_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15388_ _07327_ _07453_ VGND VGND VPWR VPWR _07462_ sky130_fd_sc_hd__nand2_1
X_18176_ _10025_ _09822_ VGND VGND VPWR VPWR _10027_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17127_ _09071_ VGND VGND VPWR VPWR _09082_ sky130_fd_sc_hd__buf_1
XFILLER_0_41_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire480 net481 VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__buf_1
X_14339_ _06556_ VGND VGND VPWR VPWR _00071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire491 _08243_ VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__buf_1
XFILLER_0_64_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17058_ net1807 net2171 VGND VGND VPWR VPWR _09017_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16009_ _08014_ _08076_ VGND VGND VPWR VPWR _08077_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20971_ net5621 net5831 VGND VGND VPWR VPWR _00987_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22710_ _02648_ VGND VGND VPWR VPWR _00596_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23690_ net933 _03555_ VGND VGND VPWR VPWR _03557_ sky130_fd_sc_hd__nand2_1
XFILLER_0_177_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_189_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6829 net6830 VGND VGND VPWR VPWR net6829 sky130_fd_sc_hd__buf_1
XFILLER_0_94_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22641_ net1724 net3076 net2457 _02605_ net8891 VGND VGND VPWR VPWR _00570_ sky130_fd_sc_hd__o311a_1
XFILLER_0_193_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25360_ clknet_leaf_57_clk _00243_ net8718 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult2\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_22572_ net3768 VGND VGND VPWR VPWR _02553_ sky130_fd_sc_hd__buf_1
XFILLER_0_111_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24311_ pid_q.prev_int\[9\] VGND VGND VPWR VPWR _04171_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21523_ pid_d.prev_error\[3\] net5970 VGND VGND VPWR VPWR _01536_ sky130_fd_sc_hd__xnor2_1
X_25291_ clknet_leaf_88_clk _00174_ net8420 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.d\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6106 net6107 VGND VGND VPWR VPWR net6106 sky130_fd_sc_hd__clkbuf_1
X_24242_ _04101_ _04102_ VGND VGND VPWR VPWR _04103_ sky130_fd_sc_hd__and2b_1
X_21454_ net5766 net5529 VGND VGND VPWR VPWR _01467_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6128 net6130 VGND VGND VPWR VPWR net6128 sky130_fd_sc_hd__buf_1
XFILLER_0_32_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6139 net6140 VGND VGND VPWR VPWR net6139 sky130_fd_sc_hd__buf_1
Xfanout4609 pid_q.mult0.a\[8\] VGND VGND VPWR VPWR net4609 sky130_fd_sc_hd__buf_1
Xwire5405 net5398 VGND VGND VPWR VPWR net5405 sky130_fd_sc_hd__buf_1
X_20405_ _12191_ _12201_ _12202_ VGND VGND VPWR VPWR _00492_ sky130_fd_sc_hd__o21ai_1
Xwire5416 net5417 VGND VGND VPWR VPWR net5416 sky130_fd_sc_hd__clkbuf_2
X_24173_ net7511 _04033_ _04034_ VGND VGND VPWR VPWR _04035_ sky130_fd_sc_hd__and3_1
X_21385_ _01270_ _01274_ net1730 VGND VGND VPWR VPWR _01399_ sky130_fd_sc_hd__a21o_1
Xwire5427 net5428 VGND VGND VPWR VPWR net5427 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire5438 net5439 VGND VGND VPWR VPWR net5438 sky130_fd_sc_hd__buf_1
XFILLER_0_142_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4704 net4705 VGND VGND VPWR VPWR net4704 sky130_fd_sc_hd__clkbuf_2
Xwire5449 net5450 VGND VGND VPWR VPWR net5449 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23124_ _02909_ _02910_ VGND VGND VPWR VPWR _02994_ sky130_fd_sc_hd__xnor2_1
Xwire4726 net4733 VGND VGND VPWR VPWR net4726 sky130_fd_sc_hd__clkbuf_1
X_20336_ _12126_ _12137_ _12138_ VGND VGND VPWR VPWR _12139_ sky130_fd_sc_hd__and3_1
Xwire4737 net4734 VGND VGND VPWR VPWR net4737 sky130_fd_sc_hd__clkbuf_1
Xwire4748 net4749 VGND VGND VPWR VPWR net4748 sky130_fd_sc_hd__buf_1
X_23055_ net4911 VGND VGND VPWR VPWR _02925_ sky130_fd_sc_hd__inv_2
X_20267_ _12077_ cordic0.slte0.opB\[14\] net2531 VGND VGND VPWR VPWR _12078_ sky130_fd_sc_hd__mux2_1
X_22006_ net4353 _02012_ _02013_ VGND VGND VPWR VPWR _02014_ sky130_fd_sc_hd__and3_1
Xinput103 pid_d_data[15] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_1
Xinput114 pid_q_addr[0] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_1
X_20198_ net6090 net6096 net6042 net6000 VGND VGND VPWR VPWR _12023_ sky130_fd_sc_hd__a31o_1
Xinput125 pid_q_addr[5] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_1
Xinput136 pid_q_data[15] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_1
Xinput147 rstb VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_1
Xmax_length8710 net8711 VGND VGND VPWR VPWR net8710 sky130_fd_sc_hd__clkbuf_2
X_23957_ _03818_ _03820_ VGND VGND VPWR VPWR _03821_ sky130_fd_sc_hd__xor2_2
X_13710_ net909 net781 VGND VGND VPWR VPWR _05979_ sky130_fd_sc_hd__xnor2_2
X_22908_ _02794_ _02800_ net8903 VGND VGND VPWR VPWR _00642_ sky130_fd_sc_hd__o21a_1
X_14690_ net8994 net2868 net2262 net2261 VGND VGND VPWR VPWR _00141_ sky130_fd_sc_hd__a22o_1
X_23888_ _03750_ _03752_ VGND VGND VPWR VPWR _03753_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13641_ _05907_ _05910_ VGND VGND VPWR VPWR _05911_ sky130_fd_sc_hd__xnor2_1
X_25627_ clknet_leaf_117_clk _00500_ net8331 VGND VGND VPWR VPWR cordic0.slte0.opA\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_22839_ _02737_ _02738_ VGND VGND VPWR VPWR _02739_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16360_ _08421_ _08422_ VGND VGND VPWR VPWR _08423_ sky130_fd_sc_hd__xor2_1
X_13572_ net916 net913 net915 VGND VGND VPWR VPWR _05843_ sky130_fd_sc_hd__a21o_1
X_25558_ clknet_leaf_111_clk _00431_ net8365 VGND VGND VPWR VPWR cordic0.gm0.iter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire8020 net8021 VGND VGND VPWR VPWR net8020 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15311_ _07381_ _07384_ VGND VGND VPWR VPWR _07385_ sky130_fd_sc_hd__xnor2_1
Xwire8031 net8032 VGND VGND VPWR VPWR net8031 sky130_fd_sc_hd__clkbuf_1
X_24509_ _04339_ _04365_ VGND VGND VPWR VPWR _04366_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_125_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8042 net8045 VGND VGND VPWR VPWR net8042 sky130_fd_sc_hd__clkbuf_1
Xfanout6501 net6503 VGND VGND VPWR VPWR net6501 sky130_fd_sc_hd__buf_2
X_16291_ _08249_ net1251 _08354_ VGND VGND VPWR VPWR _08355_ sky130_fd_sc_hd__o21a_1
X_25489_ clknet_leaf_48_clk _00369_ net8779 VGND VGND VPWR VPWR svm0.tA\[11\] sky130_fd_sc_hd__dfrtp_1
Xwire8053 net8046 VGND VGND VPWR VPWR net8053 sky130_fd_sc_hd__buf_1
Xfanout6512 net6528 VGND VGND VPWR VPWR net6512 sky130_fd_sc_hd__buf_1
XFILLER_0_13_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7330 net7331 VGND VGND VPWR VPWR net7330 sky130_fd_sc_hd__clkbuf_1
Xwire8075 net8076 VGND VGND VPWR VPWR net8075 sky130_fd_sc_hd__clkbuf_1
X_18030_ _09878_ net3235 VGND VGND VPWR VPWR _09881_ sky130_fd_sc_hd__xnor2_2
X_15242_ net3549 net3528 VGND VGND VPWR VPWR _07316_ sky130_fd_sc_hd__nor2_1
Xwire8086 net8087 VGND VGND VPWR VPWR net8086 sky130_fd_sc_hd__clkbuf_1
Xwire7341 net7342 VGND VGND VPWR VPWR net7341 sky130_fd_sc_hd__buf_1
XFILLER_0_48_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8097 net96 VGND VGND VPWR VPWR net8097 sky130_fd_sc_hd__clkbuf_1
Xfanout6567 net6576 VGND VGND VPWR VPWR net6567 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire7363 matmul0.alpha_pass\[1\] VGND VGND VPWR VPWR net7363 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6640 net6638 VGND VGND VPWR VPWR net6640 sky130_fd_sc_hd__buf_1
Xwire7385 matmul0.matmul_stage_inst.f\[5\] VGND VGND VPWR VPWR net7385 sky130_fd_sc_hd__clkbuf_1
Xwire6651 net6652 VGND VGND VPWR VPWR net6651 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15173_ net4221 net4219 net4181 net4179 VGND VGND VPWR VPWR _07247_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7396 net7397 VGND VGND VPWR VPWR net7396 sky130_fd_sc_hd__clkbuf_1
Xwire6662 net6660 VGND VGND VPWR VPWR net6662 sky130_fd_sc_hd__buf_1
Xwire6673 net6672 VGND VGND VPWR VPWR net6673 sky130_fd_sc_hd__clkbuf_2
Xwire6684 net6685 VGND VGND VPWR VPWR net6684 sky130_fd_sc_hd__buf_1
X_14124_ net1597 _06221_ VGND VGND VPWR VPWR _06386_ sky130_fd_sc_hd__nor2_1
Xfanout5888 net5895 VGND VGND VPWR VPWR net5888 sky130_fd_sc_hd__clkbuf_1
Xwire6695 net6696 VGND VGND VPWR VPWR net6695 sky130_fd_sc_hd__clkbuf_1
Xwire5950 net5951 VGND VGND VPWR VPWR net5950 sky130_fd_sc_hd__buf_1
XFILLER_0_104_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19981_ _11788_ _11811_ VGND VGND VPWR VPWR _11812_ sky130_fd_sc_hd__xnor2_2
Xwire5961 net5963 VGND VGND VPWR VPWR net5961 sky130_fd_sc_hd__buf_1
Xwire5972 pid_d.curr_error\[1\] VGND VGND VPWR VPWR net5972 sky130_fd_sc_hd__buf_1
Xwire5983 pid_d.curr_int\[2\] VGND VGND VPWR VPWR net5983 sky130_fd_sc_hd__clkbuf_2
X_14055_ _06282_ _06318_ VGND VGND VPWR VPWR _06319_ sky130_fd_sc_hd__xnor2_1
X_18932_ net2537 VGND VGND VPWR VPWR _10771_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13006_ _05262_ _05278_ VGND VGND VPWR VPWR _05279_ sky130_fd_sc_hd__xnor2_1
X_18863_ _10703_ _10680_ _10704_ VGND VGND VPWR VPWR _10705_ sky130_fd_sc_hd__a21o_1
XFILLER_0_193_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17814_ net3977 _09664_ VGND VGND VPWR VPWR _09665_ sky130_fd_sc_hd__xnor2_2
X_18794_ net6897 net6808 VGND VGND VPWR VPWR _10638_ sky130_fd_sc_hd__xnor2_2
X_17745_ net8998 _08819_ net8060 VGND VGND VPWR VPWR _00438_ sky130_fd_sc_hd__o21a_1
X_14957_ net3575 net3571 net4137 net4130 VGND VGND VPWR VPWR _07031_ sky130_fd_sc_hd__o22a_1
X_13908_ net7633 net7605 VGND VGND VPWR VPWR _06174_ sky130_fd_sc_hd__nand2_1
X_17676_ svm0.tA\[3\] _09554_ _09555_ VGND VGND VPWR VPWR _09556_ sky130_fd_sc_hd__a21oi_1
X_14888_ net6620 net6638 matmul0.matmul_stage_inst.f\[0\] VGND VGND VPWR VPWR _06962_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_134_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19415_ _11243_ _11251_ net763 VGND VGND VPWR VPWR _11252_ sky130_fd_sc_hd__or3b_1
XFILLER_0_76_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16627_ matmul0.matmul_stage_inst.mult2\[1\] matmul0.matmul_stage_inst.mult1\[1\]
+ matmul0.matmul_stage_inst.mult2\[0\] matmul0.matmul_stage_inst.mult1\[0\] VGND VGND
+ VPWR VPWR _08666_ sky130_fd_sc_hd__o211ai_2
X_13839_ net7615 net1148 net1563 VGND VGND VPWR VPWR _06106_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19346_ _11180_ _11182_ VGND VGND VPWR VPWR _11183_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16558_ _08604_ _08616_ VGND VGND VPWR VPWR _08617_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15509_ _07476_ _07581_ VGND VGND VPWR VPWR _07582_ sky130_fd_sc_hd__xnor2_2
X_19277_ _10907_ _10908_ VGND VGND VPWR VPWR _11114_ sky130_fd_sc_hd__nand2_1
X_16489_ _08521_ _08532_ _08504_ VGND VGND VPWR VPWR _08549_ sky130_fd_sc_hd__a21o_1
Xfanout8492 net8509 VGND VGND VPWR VPWR net8492 sky130_fd_sc_hd__clkbuf_1
X_18228_ _10053_ _10078_ VGND VGND VPWR VPWR _10079_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout7791 svm0.periodTop\[6\] VGND VGND VPWR VPWR net7791 sky130_fd_sc_hd__buf_1
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18159_ _09769_ _09770_ VGND VGND VPWR VPWR _10010_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21170_ net3807 _01184_ _01185_ VGND VGND VPWR VPWR _01186_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20121_ _11941_ _11948_ VGND VGND VPWR VPWR _11949_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2609 _08925_ VGND VGND VPWR VPWR net2609 sky130_fd_sc_hd__buf_1
X_20052_ net3132 net6077 _11880_ VGND VGND VPWR VPWR _11881_ sky130_fd_sc_hd__a21oi_1
Xwire1908 _06850_ VGND VGND VPWR VPWR net1908 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1919 net1920 VGND VGND VPWR VPWR net1919 sky130_fd_sc_hd__clkbuf_1
X_24860_ net3710 VGND VGND VPWR VPWR _04664_ sky130_fd_sc_hd__clkbuf_1
X_23811_ _03584_ _03585_ _03658_ VGND VGND VPWR VPWR _03676_ sky130_fd_sc_hd__a21o_1
XFILLER_0_84_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24791_ _04613_ _04616_ VGND VGND VPWR VPWR _04617_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length7305 matmul0.alpha_pass\[6\] VGND VGND VPWR VPWR net7305 sky130_fd_sc_hd__clkbuf_1
Xmax_length7316 matmul0.alpha_pass\[5\] VGND VGND VPWR VPWR net7316 sky130_fd_sc_hd__clkbuf_1
X_23742_ net5146 net5122 net5097 net4482 VGND VGND VPWR VPWR _03608_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_75_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20954_ net5635 net5759 net3836 _00969_ VGND VGND VPWR VPWR _00970_ sky130_fd_sc_hd__a31o_1
XFILLER_0_191_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23673_ _03524_ _03539_ VGND VGND VPWR VPWR _03540_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20885_ net5575 net5832 VGND VGND VPWR VPWR _00901_ sky130_fd_sc_hd__nand2_1
X_25412_ clknet_leaf_80_clk _00295_ net8494 VGND VGND VPWR VPWR matmul0.a\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_177_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22624_ net7203 _02590_ VGND VGND VPWR VPWR _02594_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25343_ clknet_leaf_56_clk _00226_ net8714 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22555_ net5964 net3017 net2461 VGND VGND VPWR VPWR _02540_ sky130_fd_sc_hd__and3_1
XFILLER_0_106_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21506_ net948 _01518_ VGND VGND VPWR VPWR _01519_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_173_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25274_ clknet_leaf_76_clk _00157_ net8458 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.c\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_22486_ net5671 _02483_ net5390 VGND VGND VPWR VPWR _02487_ sky130_fd_sc_hd__o21a_1
X_24225_ net2024 net1657 VGND VGND VPWR VPWR _04086_ sky130_fd_sc_hd__xnor2_2
X_21437_ net5618 net5673 VGND VGND VPWR VPWR _01450_ sky130_fd_sc_hd__nand2_1
Xwire5213 net5214 VGND VGND VPWR VPWR net5213 sky130_fd_sc_hd__buf_1
Xwire5224 net5225 VGND VGND VPWR VPWR net5224 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5235 net5237 VGND VGND VPWR VPWR net5235 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24156_ _03920_ _04017_ _03932_ VGND VGND VPWR VPWR _04018_ sky130_fd_sc_hd__o21ai_1
Xwire5246 net5247 VGND VGND VPWR VPWR net5246 sky130_fd_sc_hd__buf_1
Xwire4512 net4513 VGND VGND VPWR VPWR net4512 sky130_fd_sc_hd__buf_1
Xwire5257 net5258 VGND VGND VPWR VPWR net5257 sky130_fd_sc_hd__clkbuf_1
X_21368_ net5944 net5399 VGND VGND VPWR VPWR _01382_ sky130_fd_sc_hd__nand2_1
Xwire4523 net4524 VGND VGND VPWR VPWR net4523 sky130_fd_sc_hd__buf_1
Xwire5268 net5269 VGND VGND VPWR VPWR net5268 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4534 net4535 VGND VGND VPWR VPWR net4534 sky130_fd_sc_hd__buf_1
Xwire5279 net5280 VGND VGND VPWR VPWR net5279 sky130_fd_sc_hd__buf_1
XFILLER_0_102_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23107_ _02974_ _02975_ VGND VGND VPWR VPWR _02977_ sky130_fd_sc_hd__nor2_1
Xwire4545 net4546 VGND VGND VPWR VPWR net4545 sky130_fd_sc_hd__buf_1
Xwire3800 net3801 VGND VGND VPWR VPWR net3800 sky130_fd_sc_hd__clkbuf_1
X_20319_ cordic0.slte0.opA\[2\] _12112_ VGND VGND VPWR VPWR _12123_ sky130_fd_sc_hd__or2_1
Xwire3811 net3812 VGND VGND VPWR VPWR net3811 sky130_fd_sc_hd__buf_1
X_24087_ _03948_ _03949_ VGND VGND VPWR VPWR _03950_ sky130_fd_sc_hd__nand2_1
Xwire3822 _00978_ VGND VGND VPWR VPWR net3822 sky130_fd_sc_hd__clkbuf_1
Xwire4567 net4569 VGND VGND VPWR VPWR net4567 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21299_ net1050 _01313_ VGND VGND VPWR VPWR _01314_ sky130_fd_sc_hd__xor2_1
Xwire4578 net4579 VGND VGND VPWR VPWR net4578 sky130_fd_sc_hd__clkbuf_1
Xwire3833 net3834 VGND VGND VPWR VPWR net3833 sky130_fd_sc_hd__clkbuf_1
Xwire4589 net4590 VGND VGND VPWR VPWR net4589 sky130_fd_sc_hd__buf_1
X_23038_ _02894_ _02907_ VGND VGND VPWR VPWR _02908_ sky130_fd_sc_hd__xnor2_2
Xwire3855 _11559_ VGND VGND VPWR VPWR net3855 sky130_fd_sc_hd__clkbuf_1
Xwire3866 _11289_ VGND VGND VPWR VPWR net3866 sky130_fd_sc_hd__buf_1
Xwire3877 _11025_ VGND VGND VPWR VPWR net3877 sky130_fd_sc_hd__buf_1
Xwire3888 _10898_ VGND VGND VPWR VPWR net3888 sky130_fd_sc_hd__dlymetal6s2s_1
X_15860_ net2699 net2727 VGND VGND VPWR VPWR _07929_ sky130_fd_sc_hd__nand2_1
X_14811_ net9065 net2876 net2854 _06922_ VGND VGND VPWR VPWR _00177_ sky130_fd_sc_hd__o22a_1
XFILLER_0_192_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15791_ net1097 _07773_ net1099 VGND VGND VPWR VPWR _07861_ sky130_fd_sc_hd__o21a_1
X_24989_ _04749_ VGND VGND VPWR VPWR _00774_ sky130_fd_sc_hd__clkbuf_1
X_17530_ net6686 _09412_ _09413_ VGND VGND VPWR VPWR _00405_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_54_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14742_ net7448 net7156 VGND VGND VPWR VPWR _06876_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length8584 net8581 VGND VGND VPWR VPWR net8584 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_168_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17461_ svm0.delta\[4\] _09354_ VGND VGND VPWR VPWR _09355_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14673_ net9081 net2869 _06822_ net2865 VGND VGND VPWR VPWR _00137_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19200_ net3876 _11036_ VGND VGND VPWR VPWR _11037_ sky130_fd_sc_hd__xnor2_1
X_13624_ _05892_ _05893_ VGND VGND VPWR VPWR _05894_ sky130_fd_sc_hd__and2b_1
X_16412_ _08467_ _08473_ VGND VGND VPWR VPWR _08474_ sky130_fd_sc_hd__xnor2_2
X_17392_ svm0.delta\[7\] VGND VGND VPWR VPWR _09299_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19131_ net3216 _10808_ _10967_ VGND VGND VPWR VPWR _10968_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13555_ net7638 net1975 net2311 VGND VGND VPWR VPWR _05826_ sky130_fd_sc_hd__and3_1
XFILLER_0_109_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16343_ _08402_ _08404_ VGND VGND VPWR VPWR _08406_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_183_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout7043 net7047 VGND VGND VPWR VPWR net7043 sky130_fd_sc_hd__buf_1
Xfanout6320 net6330 VGND VGND VPWR VPWR net6320 sky130_fd_sc_hd__buf_1
X_19062_ _10827_ _10811_ VGND VGND VPWR VPWR _10899_ sky130_fd_sc_hd__xnor2_2
X_16274_ net978 _08337_ VGND VGND VPWR VPWR _08338_ sky130_fd_sc_hd__xnor2_1
X_13486_ _05741_ _05758_ VGND VGND VPWR VPWR _05759_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6353 net6361 VGND VGND VPWR VPWR net6353 sky130_fd_sc_hd__buf_1
X_18013_ net7082 net7108 VGND VGND VPWR VPWR _09864_ sky130_fd_sc_hd__or2_1
X_15225_ _07278_ _07280_ _07298_ VGND VGND VPWR VPWR _07299_ sky130_fd_sc_hd__o21a_1
Xwire7160 net7161 VGND VGND VPWR VPWR net7160 sky130_fd_sc_hd__clkbuf_2
Xfanout5630 pid_d.mult0.a\[1\] VGND VGND VPWR VPWR net5630 sky130_fd_sc_hd__buf_1
Xwire7171 matmul0.cos\[9\] VGND VGND VPWR VPWR net7171 sky130_fd_sc_hd__clkbuf_1
Xfanout6375 net6378 VGND VGND VPWR VPWR net6375 sky130_fd_sc_hd__buf_1
Xwire7182 matmul0.cos\[1\] VGND VGND VPWR VPWR net7182 sky130_fd_sc_hd__buf_1
Xwire7193 net7194 VGND VGND VPWR VPWR net7193 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6470 net6473 VGND VGND VPWR VPWR net6470 sky130_fd_sc_hd__buf_1
XFILLER_0_160_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15156_ _06992_ net4186 VGND VGND VPWR VPWR _07230_ sky130_fd_sc_hd__nor2_1
Xfanout4940 net4946 VGND VGND VPWR VPWR net4940 sky130_fd_sc_hd__clkbuf_1
Xfanout5685 net5697 VGND VGND VPWR VPWR net5685 sky130_fd_sc_hd__buf_1
XFILLER_0_196_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout4962 net4976 VGND VGND VPWR VPWR net4962 sky130_fd_sc_hd__buf_1
XFILLER_0_50_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14107_ _06332_ _06351_ VGND VGND VPWR VPWR _06369_ sky130_fd_sc_hd__nor2_2
Xwire5780 net5781 VGND VGND VPWR VPWR net5780 sky130_fd_sc_hd__buf_1
XFILLER_0_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19964_ net6107 _11758_ _11792_ _11793_ _11794_ VGND VGND VPWR VPWR _11795_ sky130_fd_sc_hd__a41o_1
X_15087_ net2800 _07148_ _07160_ VGND VGND VPWR VPWR _07161_ sky130_fd_sc_hd__a21bo_1
Xwire5791 pid_d.mult0.b\[8\] VGND VGND VPWR VPWR net5791 sky130_fd_sc_hd__clkbuf_1
X_14038_ _06300_ _06301_ VGND VGND VPWR VPWR _06302_ sky130_fd_sc_hd__xnor2_1
X_18915_ net6828 _10279_ _10754_ _10278_ VGND VGND VPWR VPWR _10755_ sky130_fd_sc_hd__a22o_1
X_19895_ _11715_ _11727_ VGND VGND VPWR VPWR _11728_ sky130_fd_sc_hd__or2_1
XFILLER_0_180_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18846_ _10629_ _10647_ VGND VGND VPWR VPWR _10689_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18777_ net764 _10603_ VGND VGND VPWR VPWR _10621_ sky130_fd_sc_hd__or2b_1
X_15989_ net2712 net3394 _08053_ VGND VGND VPWR VPWR _08057_ sky130_fd_sc_hd__nand3_1
XFILLER_0_179_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17728_ net8059 net6522 VGND VGND VPWR VPWR _09587_ sky130_fd_sc_hd__nand2_1
X_17659_ net6723 svm0.tA\[6\] VGND VGND VPWR VPWR _09539_ sky130_fd_sc_hd__and2b_1
XFILLER_0_159_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20670_ _12435_ _12446_ VGND VGND VPWR VPWR _12447_ sky130_fd_sc_hd__or2_1
XFILLER_0_174_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19329_ _11162_ _11165_ net6315 VGND VGND VPWR VPWR _11166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22340_ _02228_ net2472 _02342_ VGND VGND VPWR VPWR _02343_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22271_ _02169_ VGND VGND VPWR VPWR _02275_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24010_ net5027 net4500 net5048 VGND VGND VPWR VPWR _03873_ sky130_fd_sc_hd__a21o_1
X_21222_ net861 _01236_ _01237_ VGND VGND VPWR VPWR _01238_ sky130_fd_sc_hd__o21a_1
Xhold110 matmul0.matmul_stage_inst.c\[3\] VGND VGND VPWR VPWR net9063 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 cordic0.sin\[11\] VGND VGND VPWR VPWR net9074 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold132 cordic0.sin\[8\] VGND VGND VPWR VPWR net9085 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold143 svm0.tB\[14\] VGND VGND VPWR VPWR net9096 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 pid_q.prev_error\[15\] VGND VGND VPWR VPWR net9107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 svm0.tC\[6\] VGND VGND VPWR VPWR net9118 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3107 net3108 VGND VGND VPWR VPWR net3107 sky130_fd_sc_hd__buf_1
X_21153_ net5599 net5955 VGND VGND VPWR VPWR _01169_ sky130_fd_sc_hd__nand2_1
Xhold176 svm0.tB\[13\] VGND VGND VPWR VPWR net9129 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3118 net3119 VGND VGND VPWR VPWR net3118 sky130_fd_sc_hd__buf_1
Xwire3129 _11572_ VGND VGND VPWR VPWR net3129 sky130_fd_sc_hd__buf_1
Xhold187 svm0.tB\[4\] VGND VGND VPWR VPWR net9140 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2406 net2407 VGND VGND VPWR VPWR net2406 sky130_fd_sc_hd__clkbuf_1
Xhold198 pid_q.curr_error\[14\] VGND VGND VPWR VPWR net9151 sky130_fd_sc_hd__dlygate4sd3_1
X_20104_ _11878_ _11929_ _11931_ VGND VGND VPWR VPWR _11932_ sky130_fd_sc_hd__a21oi_1
Xwire2417 net2418 VGND VGND VPWR VPWR net2417 sky130_fd_sc_hd__clkbuf_1
X_21084_ _01088_ _01090_ VGND VGND VPWR VPWR _01100_ sky130_fd_sc_hd__xor2_2
Xwire2428 _03225_ VGND VGND VPWR VPWR net2428 sky130_fd_sc_hd__buf_1
Xwire2439 net2440 VGND VGND VPWR VPWR net2439 sky130_fd_sc_hd__buf_1
Xwire1705 _02223_ VGND VGND VPWR VPWR net1705 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24912_ net1636 VGND VGND VPWR VPWR _04702_ sky130_fd_sc_hd__buf_1
Xwire1716 _01887_ VGND VGND VPWR VPWR net1716 sky130_fd_sc_hd__buf_1
X_20035_ net6028 net3136 _11588_ _11451_ _11864_ VGND VGND VPWR VPWR _11865_ sky130_fd_sc_hd__a221o_1
X_25892_ clknet_leaf_15_clk _00765_ net8622 VGND VGND VPWR VPWR pid_q.kp\[4\] sky130_fd_sc_hd__dfrtp_1
Xwire1727 _01461_ VGND VGND VPWR VPWR net1727 sky130_fd_sc_hd__buf_1
Xwire1738 _12418_ VGND VGND VPWR VPWR net1738 sky130_fd_sc_hd__buf_1
Xwire1749 net1750 VGND VGND VPWR VPWR net1749 sky130_fd_sc_hd__buf_1
X_24843_ _04534_ _04654_ net4897 _04642_ VGND VGND VPWR VPWR _00723_ sky130_fd_sc_hd__a2bb2o_1
X_24774_ net7980 _04601_ VGND VGND VPWR VPWR _04602_ sky130_fd_sc_hd__xor2_1
X_21986_ _01992_ _01993_ _01990_ VGND VGND VPWR VPWR _01994_ sky130_fd_sc_hd__a21oi_1
Xmax_length7135 net7136 VGND VGND VPWR VPWR net7135 sky130_fd_sc_hd__buf_1
X_23725_ net4587 net4963 VGND VGND VPWR VPWR _03591_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length7157 matmul0.sin\[3\] VGND VGND VPWR VPWR net7157 sky130_fd_sc_hd__clkbuf_1
X_20937_ _00939_ _00940_ VGND VGND VPWR VPWR _00953_ sky130_fd_sc_hd__xor2_1
XFILLER_0_96_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23656_ _03518_ _03522_ VGND VGND VPWR VPWR _03523_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20868_ _00881_ net3836 _00883_ VGND VGND VPWR VPWR _00884_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_154_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length6478 net6475 VGND VGND VPWR VPWR net6478 sky130_fd_sc_hd__buf_1
XFILLER_0_113_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22607_ _02579_ _02580_ net3770 VGND VGND VPWR VPWR _02581_ sky130_fd_sc_hd__and3b_1
XFILLER_0_119_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23587_ _03357_ _03358_ _03454_ VGND VGND VPWR VPWR _03455_ sky130_fd_sc_hd__a21o_1
XFILLER_0_165_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20799_ _00810_ _00814_ VGND VGND VPWR VPWR _00815_ sky130_fd_sc_hd__nand2_1
XFILLER_0_180_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13340_ _05520_ _05522_ _05518_ VGND VGND VPWR VPWR _05613_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25326_ clknet_leaf_79_clk _00209_ net8491 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.f\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22538_ net9117 net1700 _02531_ VGND VGND VPWR VPWR _00541_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13271_ _05543_ net1136 net1137 VGND VGND VPWR VPWR _05544_ sky130_fd_sc_hd__a21bo_1
X_25257_ clknet_leaf_70_clk _00140_ net8457 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.b\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_22469_ net1169 _02344_ net2060 VGND VGND VPWR VPWR _02470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5010 net4999 VGND VGND VPWR VPWR net5010 sky130_fd_sc_hd__clkbuf_1
X_15010_ _07082_ _07083_ VGND VGND VPWR VPWR _07084_ sky130_fd_sc_hd__or2_1
X_24208_ net3040 _03973_ _04068_ VGND VGND VPWR VPWR _04069_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_122_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5032 net5034 VGND VGND VPWR VPWR net5032 sky130_fd_sc_hd__clkbuf_1
X_25188_ clknet_leaf_62_clk _00077_ net8671 VGND VGND VPWR VPWR matmul0.a_in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire5054 net5055 VGND VGND VPWR VPWR net5054 sky130_fd_sc_hd__buf_1
Xwire5065 net5066 VGND VGND VPWR VPWR net5065 sky130_fd_sc_hd__buf_1
Xwire4320 net4318 VGND VGND VPWR VPWR net4320 sky130_fd_sc_hd__buf_1
Xwire5076 net5072 VGND VGND VPWR VPWR net5076 sky130_fd_sc_hd__clkbuf_1
X_24139_ _03994_ _04000_ VGND VGND VPWR VPWR _04001_ sky130_fd_sc_hd__xnor2_2
Xwire5087 net5088 VGND VGND VPWR VPWR net5087 sky130_fd_sc_hd__buf_1
Xwire4342 net4343 VGND VGND VPWR VPWR net4342 sky130_fd_sc_hd__clkbuf_1
Xwire5098 net5102 VGND VGND VPWR VPWR net5098 sky130_fd_sc_hd__clkbuf_1
Xwire4353 net4352 VGND VGND VPWR VPWR net4353 sky130_fd_sc_hd__clkbuf_1
Xwire4375 net4368 VGND VGND VPWR VPWR net4375 sky130_fd_sc_hd__buf_1
Xwire3641 _06533_ VGND VGND VPWR VPWR net3641 sky130_fd_sc_hd__buf_1
Xwire4386 net4387 VGND VGND VPWR VPWR net4386 sky130_fd_sc_hd__clkbuf_1
X_16961_ _08850_ VGND VGND VPWR VPWR _08924_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_60_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3652 net3653 VGND VGND VPWR VPWR net3652 sky130_fd_sc_hd__clkbuf_1
Xwire4397 net4398 VGND VGND VPWR VPWR net4397 sky130_fd_sc_hd__clkbuf_1
Xwire3663 net3664 VGND VGND VPWR VPWR net3663 sky130_fd_sc_hd__clkbuf_1
Xwire3674 _05709_ VGND VGND VPWR VPWR net3674 sky130_fd_sc_hd__buf_1
X_18700_ net2588 net6785 VGND VGND VPWR VPWR _10546_ sky130_fd_sc_hd__nor2_1
Xwire3685 net3686 VGND VGND VPWR VPWR net3685 sky130_fd_sc_hd__buf_1
Xwire2940 net2941 VGND VGND VPWR VPWR net2940 sky130_fd_sc_hd__clkbuf_1
X_15912_ _07852_ _07854_ _07980_ VGND VGND VPWR VPWR _07981_ sky130_fd_sc_hd__a21o_1
Xwire2951 net2952 VGND VGND VPWR VPWR net2951 sky130_fd_sc_hd__clkbuf_1
Xwire3696 _04886_ VGND VGND VPWR VPWR net3696 sky130_fd_sc_hd__buf_1
X_19680_ net6220 net3195 net3162 _11466_ VGND VGND VPWR VPWR _11516_ sky130_fd_sc_hd__or4_1
X_16892_ cordic0.slte0.opA\[17\] _08855_ VGND VGND VPWR VPWR _08856_ sky130_fd_sc_hd__or2_1
Xwire2962 net2963 VGND VGND VPWR VPWR net2962 sky130_fd_sc_hd__clkbuf_1
Xwire2984 net2985 VGND VGND VPWR VPWR net2984 sky130_fd_sc_hd__buf_1
X_18631_ net6827 net3966 VGND VGND VPWR VPWR _10478_ sky130_fd_sc_hd__or2_1
Xwire2995 net2996 VGND VGND VPWR VPWR net2995 sky130_fd_sc_hd__clkbuf_1
X_15843_ _07911_ _07912_ VGND VGND VPWR VPWR _07913_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18562_ _10328_ _10346_ _10394_ VGND VGND VPWR VPWR _10410_ sky130_fd_sc_hd__a21o_1
X_12986_ _05257_ _05258_ VGND VGND VPWR VPWR _05259_ sky130_fd_sc_hd__xor2_1
X_15774_ net2761 _07840_ _07842_ net2640 VGND VGND VPWR VPWR _07844_ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17513_ _09315_ _09395_ net3271 VGND VGND VPWR VPWR _09399_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_111_Left_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length8381 net8382 VGND VGND VPWR VPWR net8381 sky130_fd_sc_hd__buf_1
X_14725_ _06824_ _06863_ VGND VGND VPWR VPWR _06864_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18493_ _10342_ VGND VGND VPWR VPWR _10343_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17444_ _09340_ VGND VGND VPWR VPWR _00392_ sky130_fd_sc_hd__clkbuf_1
X_14656_ net8965 _06801_ _06812_ VGND VGND VPWR VPWR _00132_ sky130_fd_sc_hd__a21o_1
XFILLER_0_156_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13607_ _05875_ _05876_ VGND VGND VPWR VPWR _05877_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17375_ _09195_ VGND VGND VPWR VPWR _09286_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14587_ net7214 net5198 VGND VGND VPWR VPWR _06762_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_40_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19114_ _10940_ _10949_ _10950_ VGND VGND VPWR VPWR _10951_ sky130_fd_sc_hd__nand3_1
X_16326_ net2772 net2204 VGND VGND VPWR VPWR _08389_ sky130_fd_sc_hd__nand2_1
X_13538_ net7722 net1313 VGND VGND VPWR VPWR _05809_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19045_ net6261 net6245 VGND VGND VPWR VPWR _10882_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13469_ net1131 _05588_ _05581_ VGND VGND VPWR VPWR _05742_ sky130_fd_sc_hd__o21a_1
X_16257_ net2246 _08040_ VGND VGND VPWR VPWR _08321_ sky130_fd_sc_hd__nor2_1
XFILLER_0_180_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout6194 net6214 VGND VGND VPWR VPWR net6194 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_120_Left_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15208_ _07246_ _07247_ VGND VGND VPWR VPWR _07282_ sky130_fd_sc_hd__xnor2_1
Xfanout5471 net5483 VGND VGND VPWR VPWR net5471 sky130_fd_sc_hd__clkbuf_1
X_16188_ net2211 net2215 VGND VGND VPWR VPWR _08253_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15139_ _07202_ _07203_ _07212_ VGND VGND VPWR VPWR _07213_ sky130_fd_sc_hd__or3_1
XFILLER_0_121_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19947_ _11777_ _11778_ VGND VGND VPWR VPWR _11779_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19878_ _11708_ _11710_ VGND VGND VPWR VPWR _11711_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18829_ net6868 net3920 VGND VGND VPWR VPWR _10672_ sky130_fd_sc_hd__xnor2_1
X_21840_ _01847_ _01848_ VGND VGND VPWR VPWR _01849_ sky130_fd_sc_hd__xor2_1
XFILLER_0_172_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21771_ net5857 net5376 VGND VGND VPWR VPWR _01781_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23510_ net934 _03378_ VGND VGND VPWR VPWR _03379_ sky130_fd_sc_hd__xnor2_2
X_20722_ net6035 _12481_ VGND VGND VPWR VPWR _12494_ sky130_fd_sc_hd__nor2_1
XFILLER_0_176_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24490_ _04343_ _04346_ VGND VGND VPWR VPWR _04347_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_176_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8619 net8617 VGND VGND VPWR VPWR net8619 sky130_fd_sc_hd__clkbuf_2
X_23441_ pid_q.curr_int\[0\] pid_q.prev_int\[0\] VGND VGND VPWR VPWR _03311_ sky130_fd_sc_hd__xor2_1
Xmax_length4317 net4314 VGND VGND VPWR VPWR net4317 sky130_fd_sc_hd__buf_1
XFILLER_0_46_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20653_ net1394 _12430_ VGND VGND VPWR VPWR _12431_ sky130_fd_sc_hd__xor2_1
XFILLER_0_135_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7907 net7908 VGND VGND VPWR VPWR net7907 sky130_fd_sc_hd__buf_1
Xwire309 net310 VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__clkbuf_1
Xmax_length3605 net3606 VGND VGND VPWR VPWR net3605 sky130_fd_sc_hd__buf_1
XFILLER_0_162_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7929 svm0.periodTop\[1\] VGND VGND VPWR VPWR net7929 sky130_fd_sc_hd__buf_1
X_23372_ net4721 net4886 VGND VGND VPWR VPWR _03242_ sky130_fd_sc_hd__nand2_1
X_20584_ net1745 _12342_ net1742 VGND VGND VPWR VPWR _12367_ sky130_fd_sc_hd__or3_2
XFILLER_0_73_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25111_ _04852_ VGND VGND VPWR VPWR _04853_ sky130_fd_sc_hd__buf_1
XFILLER_0_6_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22323_ net336 _02326_ VGND VGND VPWR VPWR _02327_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_190_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25042_ net331 net1630 _04792_ net9174 _04793_ VGND VGND VPWR VPWR _00783_ sky130_fd_sc_hd__a221o_1
XFILLER_0_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22254_ _02256_ _02257_ VGND VGND VPWR VPWR _02259_ sky130_fd_sc_hd__or2_1
XFILLER_0_143_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21205_ net761 net760 _01220_ VGND VGND VPWR VPWR _01221_ sky130_fd_sc_hd__a21o_1
X_22185_ _02059_ _02161_ VGND VGND VPWR VPWR _02190_ sky130_fd_sc_hd__nor2_1
X_21136_ _01150_ _01151_ VGND VGND VPWR VPWR _01152_ sky130_fd_sc_hd__xnor2_1
Xwire2203 _08677_ VGND VGND VPWR VPWR net2203 sky130_fd_sc_hd__clkbuf_1
Xwire2214 _07900_ VGND VGND VPWR VPWR net2214 sky130_fd_sc_hd__buf_1
Xwire2225 net2226 VGND VGND VPWR VPWR net2225 sky130_fd_sc_hd__buf_1
Xwire2236 net2237 VGND VGND VPWR VPWR net2236 sky130_fd_sc_hd__clkbuf_1
X_21067_ _01079_ _01082_ VGND VGND VPWR VPWR _01083_ sky130_fd_sc_hd__xnor2_2
Xwire1502 net1503 VGND VGND VPWR VPWR net1502 sky130_fd_sc_hd__clkbuf_1
Xwire2247 net2248 VGND VGND VPWR VPWR net2247 sky130_fd_sc_hd__clkbuf_1
Xwire2258 _06980_ VGND VGND VPWR VPWR net2258 sky130_fd_sc_hd__clkbuf_1
Xwire1513 net1514 VGND VGND VPWR VPWR net1513 sky130_fd_sc_hd__buf_1
Xwire2269 net2270 VGND VGND VPWR VPWR net2269 sky130_fd_sc_hd__clkbuf_1
Xwire1524 _07956_ VGND VGND VPWR VPWR net1524 sky130_fd_sc_hd__clkbuf_1
Xwire1535 _07766_ VGND VGND VPWR VPWR net1535 sky130_fd_sc_hd__buf_1
Xwire1546 _07244_ VGND VGND VPWR VPWR net1546 sky130_fd_sc_hd__clkbuf_1
X_20018_ _11788_ _11810_ _11847_ VGND VGND VPWR VPWR _11848_ sky130_fd_sc_hd__o21ai_4
X_25875_ clknet_leaf_15_clk _00748_ net8618 VGND VGND VPWR VPWR pid_q.ki\[3\] sky130_fd_sc_hd__dfrtp_1
Xwire1557 net1558 VGND VGND VPWR VPWR net1557 sky130_fd_sc_hd__clkbuf_1
Xwire1568 net1569 VGND VGND VPWR VPWR net1568 sky130_fd_sc_hd__buf_1
Xwire1579 net1580 VGND VGND VPWR VPWR net1579 sky130_fd_sc_hd__buf_1
X_12840_ net1957 _05111_ VGND VGND VPWR VPWR _05113_ sky130_fd_sc_hd__or2_1
X_24826_ net7480 net1010 net2416 VGND VGND VPWR VPWR _04646_ sky130_fd_sc_hd__a21o_1
X_12771_ _04927_ _04933_ net7800 net1615 VGND VGND VPWR VPWR _05044_ sky130_fd_sc_hd__o211a_1
X_24757_ net7996 _04580_ _04581_ net2009 VGND VGND VPWR VPWR _04587_ sky130_fd_sc_hd__a31o_1
X_21969_ _01975_ _01976_ VGND VGND VPWR VPWR _01977_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14510_ net7282 net5254 VGND VGND VPWR VPWR _06691_ sky130_fd_sc_hd__xor2_1
Xmax_length6242 net6240 VGND VGND VPWR VPWR net6242 sky130_fd_sc_hd__clkbuf_1
X_23708_ net7503 _03573_ _03574_ VGND VGND VPWR VPWR _03575_ sky130_fd_sc_hd__and3_1
X_15490_ net1274 net1875 VGND VGND VPWR VPWR _07563_ sky130_fd_sc_hd__or2_1
X_24688_ net9107 net1648 _04526_ VGND VGND VPWR VPWR _00696_ sky130_fd_sc_hd__a21o_1
XFILLER_0_167_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23639_ _03432_ _03437_ _03430_ VGND VGND VPWR VPWR _03506_ sky130_fd_sc_hd__o21a_1
X_14441_ net5210 net1293 net2889 net4407 _06634_ VGND VGND VPWR VPWR _06635_ sky130_fd_sc_hd__a221o_1
XFILLER_0_126_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length4840 net4829 VGND VGND VPWR VPWR net4840 sky130_fd_sc_hd__clkbuf_1
Xmax_length5585 net5580 VGND VGND VPWR VPWR net5585 sky130_fd_sc_hd__buf_1
X_14372_ net8295 _06575_ VGND VGND VPWR VPWR _06582_ sky130_fd_sc_hd__and2_1
Xwire810 _12245_ VGND VGND VPWR VPWR net810 sky130_fd_sc_hd__clkbuf_1
X_17160_ _09098_ _09112_ VGND VGND VPWR VPWR _09113_ sky130_fd_sc_hd__or2_1
Xmax_length5596 net5597 VGND VGND VPWR VPWR net5596 sky130_fd_sc_hd__buf_1
Xwire821 _09470_ VGND VGND VPWR VPWR net821 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire843 _05626_ VGND VGND VPWR VPWR net843 sky130_fd_sc_hd__clkbuf_2
X_13323_ net7774 _04960_ _05507_ _05506_ VGND VGND VPWR VPWR _05596_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16111_ _08094_ _08095_ _08176_ VGND VGND VPWR VPWR _08177_ sky130_fd_sc_hd__o21a_1
Xmax_length4895 net4896 VGND VGND VPWR VPWR net4895 sky130_fd_sc_hd__clkbuf_1
Xwire854 _03858_ VGND VGND VPWR VPWR net854 sky130_fd_sc_hd__buf_1
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25309_ clknet_leaf_76_clk _00192_ net8462 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.e\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire865 _12173_ VGND VGND VPWR VPWR net865 sky130_fd_sc_hd__buf_1
X_17091_ net6981 net1551 VGND VGND VPWR VPWR _09049_ sky130_fd_sc_hd__nor2_1
Xwire876 _09519_ VGND VGND VPWR VPWR net876 sky130_fd_sc_hd__clkbuf_1
Xwire887 _07777_ VGND VGND VPWR VPWR net887 sky130_fd_sc_hd__buf_1
X_13254_ net2301 net2297 VGND VGND VPWR VPWR _05527_ sky130_fd_sc_hd__nor2_1
X_16042_ net1515 _08108_ VGND VGND VPWR VPWR _08109_ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13185_ net7650 net2339 net1967 VGND VGND VPWR VPWR _05458_ sky130_fd_sc_hd__and3_1
XFILLER_0_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4150 net4151 VGND VGND VPWR VPWR net4150 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19801_ net6151 net2104 _11582_ VGND VGND VPWR VPWR _11635_ sky130_fd_sc_hd__or3_1
Xwire4161 net4162 VGND VGND VPWR VPWR net4161 sky130_fd_sc_hd__buf_1
Xwire4172 _07002_ VGND VGND VPWR VPWR net4172 sky130_fd_sc_hd__buf_1
X_17993_ net6940 _09843_ VGND VGND VPWR VPWR _09844_ sky130_fd_sc_hd__nand2_1
Xwire4183 _06994_ VGND VGND VPWR VPWR net4183 sky130_fd_sc_hd__clkbuf_1
Xwire4194 _06983_ VGND VGND VPWR VPWR net4194 sky130_fd_sc_hd__buf_1
Xwire3460 net3463 VGND VGND VPWR VPWR net3460 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_159_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19732_ net3881 net6099 _11449_ VGND VGND VPWR VPWR _11567_ sky130_fd_sc_hd__or3_1
X_16944_ net2177 _08907_ VGND VGND VPWR VPWR _08908_ sky130_fd_sc_hd__xor2_1
Xwire3471 net3472 VGND VGND VPWR VPWR net3471 sky130_fd_sc_hd__buf_1
XFILLER_0_19_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3493 net3494 VGND VGND VPWR VPWR net3493 sky130_fd_sc_hd__clkbuf_1
Xwire2770 net2771 VGND VGND VPWR VPWR net2770 sky130_fd_sc_hd__clkbuf_1
X_19663_ _11494_ _11498_ VGND VGND VPWR VPWR _11499_ sky130_fd_sc_hd__and2b_1
Xwire2781 _07140_ VGND VGND VPWR VPWR net2781 sky130_fd_sc_hd__buf_1
X_16875_ net7134 net1551 VGND VGND VPWR VPWR _08840_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2792 net2793 VGND VGND VPWR VPWR net2792 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18614_ net1196 _10452_ net814 VGND VGND VPWR VPWR _10461_ sky130_fd_sc_hd__o21a_1
X_15826_ net2660 VGND VGND VPWR VPWR _07896_ sky130_fd_sc_hd__buf_1
X_19594_ _11289_ VGND VGND VPWR VPWR _11431_ sky130_fd_sc_hd__buf_1
XFILLER_0_149_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18545_ _10384_ _10393_ VGND VGND VPWR VPWR _10394_ sky130_fd_sc_hd__xnor2_1
X_15757_ _07826_ _07827_ VGND VGND VPWR VPWR _07828_ sky130_fd_sc_hd__nand2_1
X_12969_ net1140 net1004 VGND VGND VPWR VPWR _05242_ sky130_fd_sc_hd__xor2_1
XFILLER_0_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14708_ net7456 net1908 VGND VGND VPWR VPWR _06851_ sky130_fd_sc_hd__nand2_1
X_18476_ _10322_ net1205 VGND VGND VPWR VPWR _10326_ sky130_fd_sc_hd__xor2_1
X_15688_ net3537 VGND VGND VPWR VPWR _07759_ sky130_fd_sc_hd__buf_1
XFILLER_0_142_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17427_ _09278_ _09325_ net668 VGND VGND VPWR VPWR _09327_ sky130_fd_sc_hd__o21ai_1
X_14639_ net8960 net2879 _06803_ VGND VGND VPWR VPWR _00124_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17358_ net7377 net669 VGND VGND VPWR VPWR _09271_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16309_ _08297_ _08299_ _08245_ VGND VGND VPWR VPWR _08372_ sky130_fd_sc_hd__a21bo_1
X_17289_ net6669 net1796 VGND VGND VPWR VPWR _09204_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19028_ net2528 _10832_ _10795_ net2530 net3214 VGND VGND VPWR VPWR _10865_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_140_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23990_ _03852_ _03764_ _03853_ VGND VGND VPWR VPWR _03854_ sky130_fd_sc_hd__a21o_1
X_22941_ net5327 pid_d.curr_int\[13\] _02829_ VGND VGND VPWR VPWR _02830_ sky130_fd_sc_hd__a21oi_1
X_25660_ clknet_leaf_24_clk _00533_ net8584 VGND VGND VPWR VPWR pid_d.curr_int\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_97_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22872_ _02768_ VGND VGND VPWR VPWR _00638_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24611_ _04464_ _04465_ _04412_ VGND VGND VPWR VPWR _04466_ sky130_fd_sc_hd__mux2_1
X_21823_ _01066_ net5645 VGND VGND VPWR VPWR _01832_ sky130_fd_sc_hd__nand2_2
X_25591_ clknet_leaf_91_clk _00464_ net8423 VGND VGND VPWR VPWR cordic0.cos\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_174_Right_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24542_ _04372_ _04375_ VGND VGND VPWR VPWR _04398_ sky130_fd_sc_hd__nand2_1
X_21754_ net5801 net5431 VGND VGND VPWR VPWR _01764_ sky130_fd_sc_hd__nand2_1
XFILLER_0_176_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20705_ net3139 _12477_ _12478_ VGND VGND VPWR VPWR _00516_ sky130_fd_sc_hd__a21oi_1
X_24473_ net7524 VGND VGND VPWR VPWR _04330_ sky130_fd_sc_hd__inv_2
Xwire8416 net8417 VGND VGND VPWR VPWR net8416 sky130_fd_sc_hd__clkbuf_1
X_21685_ _01689_ _01694_ VGND VGND VPWR VPWR _01696_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length4114 net4115 VGND VGND VPWR VPWR net4114 sky130_fd_sc_hd__clkbuf_1
Xwire7704 net7700 VGND VGND VPWR VPWR net7704 sky130_fd_sc_hd__buf_1
XFILLER_0_11_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8449 net8445 VGND VGND VPWR VPWR net8449 sky130_fd_sc_hd__buf_1
X_23424_ _03282_ _03293_ VGND VGND VPWR VPWR _03294_ sky130_fd_sc_hd__xnor2_1
Xwire7715 net7716 VGND VGND VPWR VPWR net7715 sky130_fd_sc_hd__buf_1
X_20636_ _12414_ _12415_ net6164 VGND VGND VPWR VPWR _12416_ sky130_fd_sc_hd__mux2_1
Xfanout6919 net6929 VGND VGND VPWR VPWR net6919 sky130_fd_sc_hd__clkbuf_2
Xwire7726 net7727 VGND VGND VPWR VPWR net7726 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7737 net7738 VGND VGND VPWR VPWR net7737 sky130_fd_sc_hd__buf_1
XFILLER_0_190_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7748 net7749 VGND VGND VPWR VPWR net7748 sky130_fd_sc_hd__clkbuf_1
Xwire7759 net7760 VGND VGND VPWR VPWR net7759 sky130_fd_sc_hd__buf_1
X_23355_ _02949_ _02951_ _03224_ VGND VGND VPWR VPWR _03225_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length2712 net2714 VGND VGND VPWR VPWR net2712 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_150_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20567_ net6470 net3927 VGND VGND VPWR VPWR _12351_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22306_ net1704 net1703 _02221_ VGND VGND VPWR VPWR _02310_ sky130_fd_sc_hd__a21bo_1
X_23286_ _03151_ _03155_ VGND VGND VPWR VPWR _03156_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20498_ net2183 _12284_ net3359 VGND VGND VPWR VPWR _12286_ sky130_fd_sc_hd__a21oi_1
X_25025_ net4457 net1631 net2394 _04778_ VGND VGND VPWR VPWR _00781_ sky130_fd_sc_hd__a22o_1
Xmax_length2789 _07138_ VGND VGND VPWR VPWR net2789 sky130_fd_sc_hd__buf_1
X_22237_ net756 _02241_ VGND VGND VPWR VPWR _02242_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_131_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22168_ net5967 VGND VGND VPWR VPWR _02174_ sky130_fd_sc_hd__inv_2
Xwire2000 net2001 VGND VGND VPWR VPWR net2000 sky130_fd_sc_hd__clkbuf_2
Xwire2011 net2012 VGND VGND VPWR VPWR net2011 sky130_fd_sc_hd__buf_1
XFILLER_0_100_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2022 net2023 VGND VGND VPWR VPWR net2022 sky130_fd_sc_hd__buf_1
X_21119_ net5585 VGND VGND VPWR VPWR _01135_ sky130_fd_sc_hd__inv_2
Xwire2033 net2034 VGND VGND VPWR VPWR net2033 sky130_fd_sc_hd__buf_1
X_22099_ net4353 _02104_ _02105_ VGND VGND VPWR VPWR _02106_ sky130_fd_sc_hd__and3_1
Xwire2044 net2045 VGND VGND VPWR VPWR net2044 sky130_fd_sc_hd__buf_1
X_14990_ net4213 net4211 net4175 net4173 VGND VGND VPWR VPWR _07064_ sky130_fd_sc_hd__o22a_1
Xwire1310 _05753_ VGND VGND VPWR VPWR net1310 sky130_fd_sc_hd__buf_1
Xwire2055 net2056 VGND VGND VPWR VPWR net2055 sky130_fd_sc_hd__buf_1
Xwire1321 net1322 VGND VGND VPWR VPWR net1321 sky130_fd_sc_hd__clkbuf_1
X_13941_ net837 net907 VGND VGND VPWR VPWR _06207_ sky130_fd_sc_hd__nand2_1
Xwire1332 _05294_ VGND VGND VPWR VPWR net1332 sky130_fd_sc_hd__clkbuf_2
Xwire2077 net2078 VGND VGND VPWR VPWR net2077 sky130_fd_sc_hd__clkbuf_2
X_25927_ clknet_leaf_1_clk _00800_ net8574 VGND VGND VPWR VPWR pid_d.prev_int\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1343 net1344 VGND VGND VPWR VPWR net1343 sky130_fd_sc_hd__clkbuf_2
Xwire2088 _12271_ VGND VGND VPWR VPWR net2088 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1354 net1355 VGND VGND VPWR VPWR net1354 sky130_fd_sc_hd__buf_1
Xwire2099 _11591_ VGND VGND VPWR VPWR net2099 sky130_fd_sc_hd__buf_1
XFILLER_0_191_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1365 net1366 VGND VGND VPWR VPWR net1365 sky130_fd_sc_hd__buf_1
Xwire1376 _04508_ VGND VGND VPWR VPWR net1376 sky130_fd_sc_hd__buf_1
X_16660_ matmul0.matmul_stage_inst.mult2\[6\] matmul0.matmul_stage_inst.mult1\[6\]
+ VGND VGND VPWR VPWR _08695_ sky130_fd_sc_hd__xor2_1
Xwire1387 _03280_ VGND VGND VPWR VPWR net1387 sky130_fd_sc_hd__clkbuf_1
X_25858_ clknet_leaf_16_clk _00731_ net8619 VGND VGND VPWR VPWR pid_q.mult0.a\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13872_ _06067_ _06138_ VGND VGND VPWR VPWR _06139_ sky130_fd_sc_hd__nor2_1
Xwire1398 net1400 VGND VGND VPWR VPWR net1398 sky130_fd_sc_hd__buf_1
X_15611_ net6542 matmul0.matmul_stage_inst.c\[15\] matmul0.matmul_stage_inst.b\[15\]
+ net6615 VGND VGND VPWR VPWR _07683_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24809_ net9151 net1644 _04542_ net227 VGND VGND VPWR VPWR _00711_ sky130_fd_sc_hd__a22o_1
X_12823_ net7727 net2978 net2336 VGND VGND VPWR VPWR _05096_ sky130_fd_sc_hd__and3_1
X_16591_ matmul0.matmul_stage_inst.mult2\[6\] net359 net2616 VGND VGND VPWR VPWR _08643_
+ sky130_fd_sc_hd__mux2_1
X_25789_ clknet_leaf_64_clk _00662_ net8672 VGND VGND VPWR VPWR matmul0.beta_pass\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18330_ _10164_ _10180_ VGND VGND VPWR VPWR _10181_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_141_Right_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15542_ net3456 net3554 VGND VGND VPWR VPWR _07615_ sky130_fd_sc_hd__nor2_1
X_12754_ net1154 _04996_ _04995_ VGND VGND VPWR VPWR _05027_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_96_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18261_ net3247 _10111_ VGND VGND VPWR VPWR _10112_ sky130_fd_sc_hd__xnor2_1
X_12685_ net5255 _04856_ net4277 _04889_ svm0.vC\[7\] VGND VGND VPWR VPWR _04958_
+ sky130_fd_sc_hd__a32oi_1
X_15473_ net1875 _07544_ _07546_ net1274 VGND VGND VPWR VPWR _07547_ sky130_fd_sc_hd__o211a_1
Xmax_length6083 net6080 VGND VGND VPWR VPWR net6083 sky130_fd_sc_hd__clkbuf_1
Xfanout8866 net8870 VGND VGND VPWR VPWR net8866 sky130_fd_sc_hd__buf_1
XFILLER_0_126_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length5360 pid_d.out\[7\] VGND VGND VPWR VPWR net5360 sky130_fd_sc_hd__buf_1
Xmax_length5371 pid_d.out_valid VGND VGND VPWR VPWR net5371 sky130_fd_sc_hd__clkbuf_1
X_17212_ _09148_ _09151_ _09146_ VGND VGND VPWR VPWR _09161_ sky130_fd_sc_hd__a21o_1
X_14424_ net8127 net3633 VGND VGND VPWR VPWR _06622_ sky130_fd_sc_hd__and2_1
Xmax_length5382 net5383 VGND VGND VPWR VPWR net5382 sky130_fd_sc_hd__clkbuf_1
Xwire8950 net8951 VGND VGND VPWR VPWR net8950 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout8899 net8907 VGND VGND VPWR VPWR net8899 sky130_fd_sc_hd__buf_1
X_18192_ net6927 net6945 VGND VGND VPWR VPWR _10043_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17143_ net4047 VGND VGND VPWR VPWR _09097_ sky130_fd_sc_hd__buf_1
Xwire640 net641 VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__buf_1
X_14355_ _06568_ VGND VGND VPWR VPWR _00075_ sky130_fd_sc_hd__clkbuf_1
Xwire651 _03181_ VGND VGND VPWR VPWR net651 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire662 _10267_ VGND VGND VPWR VPWR net662 sky130_fd_sc_hd__clkbuf_1
Xwire673 _08075_ VGND VGND VPWR VPWR net673 sky130_fd_sc_hd__buf_1
X_13306_ net7650 net2350 net2346 VGND VGND VPWR VPWR _05579_ sky130_fd_sc_hd__and3_1
Xwire684 _05305_ VGND VGND VPWR VPWR net684 sky130_fd_sc_hd__buf_1
X_14286_ net75 _06518_ _06519_ net7820 VGND VGND VPWR VPWR _00055_ sky130_fd_sc_hd__a22o_1
X_17074_ net6494 VGND VGND VPWR VPWR _09032_ sky130_fd_sc_hd__inv_2
Xmax_length3991 _09641_ VGND VGND VPWR VPWR net3991 sky130_fd_sc_hd__clkbuf_1
Xwire695 _04016_ VGND VGND VPWR VPWR net695 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13237_ net7740 net1353 _05451_ _05452_ VGND VGND VPWR VPWR _05510_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16025_ _08016_ net673 VGND VGND VPWR VPWR _08092_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13168_ _05440_ VGND VGND VPWR VPWR _05441_ sky130_fd_sc_hd__dlymetal6s2s_1
X_13099_ _05257_ _05258_ _05371_ VGND VGND VPWR VPWR _05372_ sky130_fd_sc_hd__o21a_1
X_17976_ net3245 net1779 VGND VGND VPWR VPWR _09827_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3290 net3295 VGND VGND VPWR VPWR net3290 sky130_fd_sc_hd__buf_1
X_19715_ _11548_ _11550_ VGND VGND VPWR VPWR _11551_ sky130_fd_sc_hd__xnor2_1
X_16927_ cordic0.slte0.opA\[3\] net6419 VGND VGND VPWR VPWR _08891_ sky130_fd_sc_hd__and2b_1
X_19646_ _11482_ VGND VGND VPWR VPWR _11483_ sky130_fd_sc_hd__inv_2
X_16858_ net6277 net6216 net6498 VGND VGND VPWR VPWR _08823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15809_ _07768_ net1530 VGND VGND VPWR VPWR _07879_ sky130_fd_sc_hd__nand2_1
X_19577_ _11327_ net1419 net1751 VGND VGND VPWR VPWR _11414_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_177_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16789_ _08784_ VGND VGND VPWR VPWR _00293_ sky130_fd_sc_hd__clkbuf_1
X_18528_ net1765 _10376_ VGND VGND VPWR VPWR _10377_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18459_ _10221_ net2541 VGND VGND VPWR VPWR _10309_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21470_ net5814 net5482 VGND VGND VPWR VPWR _01483_ sky130_fd_sc_hd__nand2_1
X_20421_ _12174_ _12192_ net3313 VGND VGND VPWR VPWR _12217_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5609 net5610 VGND VGND VPWR VPWR net5609 sky130_fd_sc_hd__buf_1
X_23140_ net5140 net4648 VGND VGND VPWR VPWR _03010_ sky130_fd_sc_hd__nand2_1
X_20352_ cordic0.slte0.opA\[5\] net2280 _12152_ VGND VGND VPWR VPWR _12154_ sky130_fd_sc_hd__or3_1
Xwire4908 net4909 VGND VGND VPWR VPWR net4908 sky130_fd_sc_hd__buf_1
XFILLER_0_30_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4919 net4916 VGND VGND VPWR VPWR net4919 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_144_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23071_ net5068 net4608 VGND VGND VPWR VPWR _02941_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20283_ cordic0.slte0.opA\[0\] net2091 VGND VGND VPWR VPWR _12089_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22022_ _02025_ _02028_ VGND VGND VPWR VPWR _02029_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold14 svm0.vC\[11\] VGND VGND VPWR VPWR net8967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 matmul0.matmul_stage_inst.d\[10\] VGND VGND VPWR VPWR net8978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 matmul0.matmul_stage_inst.a\[6\] VGND VGND VPWR VPWR net8989 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 net151 VGND VGND VPWR VPWR net9000 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 pid_q.target\[11\] VGND VGND VPWR VPWR net9011 sky130_fd_sc_hd__dlygate4sd3_1
X_23973_ net795 _03836_ VGND VGND VPWR VPWR _03837_ sky130_fd_sc_hd__xnor2_1
Xhold69 pid_d.curr_int\[7\] VGND VGND VPWR VPWR net9022 sky130_fd_sc_hd__dlygate4sd3_1
X_25712_ clknet_leaf_9_clk _00585_ net8552 VGND VGND VPWR VPWR pid_d.mult0.a\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_22924_ _02813_ _02814_ VGND VGND VPWR VPWR _02815_ sky130_fd_sc_hd__and2_1
X_25643_ clknet_leaf_102_clk _00516_ net8366 VGND VGND VPWR VPWR cordic0.vec\[0\]\[15\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_97_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22855_ net5364 net5980 VGND VGND VPWR VPWR _02753_ sky130_fd_sc_hd__xor2_1
XFILLER_0_168_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21806_ net4358 _01814_ _01815_ VGND VGND VPWR VPWR _01816_ sky130_fd_sc_hd__and3_1
X_22786_ pid_d.kp\[5\] _02672_ net1680 VGND VGND VPWR VPWR _02701_ sky130_fd_sc_hd__mux2_1
X_25574_ clknet_leaf_97_clk _00447_ net8398 VGND VGND VPWR VPWR cordic0.sin\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24525_ _04373_ _04381_ VGND VGND VPWR VPWR _04382_ sky130_fd_sc_hd__xnor2_1
X_21737_ _01660_ _01670_ _01665_ VGND VGND VPWR VPWR _01747_ sky130_fd_sc_hd__a21bo_1
Xwire8202 net8203 VGND VGND VPWR VPWR net8202 sky130_fd_sc_hd__clkbuf_1
Xwire8213 net8214 VGND VGND VPWR VPWR net8213 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8224 net30 VGND VGND VPWR VPWR net8224 sky130_fd_sc_hd__clkbuf_1
Xwire8235 net8236 VGND VGND VPWR VPWR net8235 sky130_fd_sc_hd__clkbuf_1
Xfanout6705 svm0.counter\[9\] VGND VGND VPWR VPWR net6705 sky130_fd_sc_hd__buf_1
Xwire8246 net8247 VGND VGND VPWR VPWR net8246 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7512 net7513 VGND VGND VPWR VPWR net7512 sky130_fd_sc_hd__buf_1
X_24456_ net928 _04313_ VGND VGND VPWR VPWR _04314_ sky130_fd_sc_hd__nand2b_2
X_21668_ _01562_ _01564_ VGND VGND VPWR VPWR _01679_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8257 net8258 VGND VGND VPWR VPWR net8257 sky130_fd_sc_hd__clkbuf_1
Xwire7523 net7524 VGND VGND VPWR VPWR net7523 sky130_fd_sc_hd__buf_1
Xwire8268 net8269 VGND VGND VPWR VPWR net8268 sky130_fd_sc_hd__clkbuf_1
Xwire7534 pid_d.iterate_enable VGND VGND VPWR VPWR net7534 sky130_fd_sc_hd__clkbuf_1
Xwire8279 net24 VGND VGND VPWR VPWR net8279 sky130_fd_sc_hd__clkbuf_1
Xmax_length3232 _10063_ VGND VGND VPWR VPWR net3232 sky130_fd_sc_hd__buf_1
Xwire6800 net6801 VGND VGND VPWR VPWR net6800 sky130_fd_sc_hd__clkbuf_1
X_23407_ net2427 _03276_ VGND VGND VPWR VPWR _03277_ sky130_fd_sc_hd__nor2_1
Xwire7545 cordic0.in_valid VGND VGND VPWR VPWR net7545 sky130_fd_sc_hd__clkbuf_1
X_20619_ _12391_ net707 _12399_ VGND VGND VPWR VPWR _12400_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24387_ _04238_ _04245_ VGND VGND VPWR VPWR _04246_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6811 net6807 VGND VGND VPWR VPWR net6811 sky130_fd_sc_hd__clkbuf_2
Xwire7556 net7557 VGND VGND VPWR VPWR net7556 sky130_fd_sc_hd__clkbuf_1
Xwire6822 net6819 VGND VGND VPWR VPWR net6822 sky130_fd_sc_hd__buf_1
XFILLER_0_85_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7567 matmul0.b_in\[7\] VGND VGND VPWR VPWR net7567 sky130_fd_sc_hd__clkbuf_1
X_21599_ net5383 _01607_ _01610_ net5897 VGND VGND VPWR VPWR _01611_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7578 net7579 VGND VGND VPWR VPWR net7578 sky130_fd_sc_hd__clkbuf_1
X_14140_ _06349_ net834 _06400_ VGND VGND VPWR VPWR _06401_ sky130_fd_sc_hd__o21a_1
Xwire6844 net6846 VGND VGND VPWR VPWR net6844 sky130_fd_sc_hd__buf_1
X_23338_ net5022 net4638 VGND VGND VPWR VPWR _03208_ sky130_fd_sc_hd__nand2_2
XFILLER_0_104_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7589 net7590 VGND VGND VPWR VPWR net7589 sky130_fd_sc_hd__clkbuf_1
Xwire6855 net6854 VGND VGND VPWR VPWR net6855 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_160_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6877 net6876 VGND VGND VPWR VPWR net6877 sky130_fd_sc_hd__buf_2
Xwire6888 net6889 VGND VGND VPWR VPWR net6888 sky130_fd_sc_hd__clkbuf_1
X_14071_ _06221_ _06174_ _06333_ net7625 VGND VGND VPWR VPWR _06334_ sky130_fd_sc_hd__o22a_1
Xmax_length2586 _09164_ VGND VGND VPWR VPWR net2586 sky130_fd_sc_hd__buf_1
X_23269_ _03133_ _03136_ _03138_ VGND VGND VPWR VPWR _03139_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_120_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13022_ net7933 _05290_ net1592 _05294_ VGND VGND VPWR VPWR _05295_ sky130_fd_sc_hd__a31o_1
X_25008_ _04762_ _04763_ VGND VGND VPWR VPWR _04764_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17830_ _09679_ _09680_ VGND VGND VPWR VPWR _09681_ sky130_fd_sc_hd__or2b_1
X_17761_ _09603_ _09611_ VGND VGND VPWR VPWR _09612_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_83_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14973_ net4191 net4185 net4162 net4158 VGND VGND VPWR VPWR _07047_ sky130_fd_sc_hd__o22a_1
XFILLER_0_195_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1140 net1141 VGND VGND VPWR VPWR net1140 sky130_fd_sc_hd__clkbuf_2
X_19500_ _11267_ _11268_ _11035_ VGND VGND VPWR VPWR _11337_ sky130_fd_sc_hd__a21o_1
Xwire1151 net1152 VGND VGND VPWR VPWR net1151 sky130_fd_sc_hd__dlymetal6s2s_1
X_16712_ _08739_ VGND VGND VPWR VPWR _00261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1162 _03708_ VGND VGND VPWR VPWR net1162 sky130_fd_sc_hd__buf_1
X_13924_ _06093_ _06094_ net7704 net1307 VGND VGND VPWR VPWR _06190_ sky130_fd_sc_hd__o211a_1
X_17692_ net1791 _09543_ _09549_ _09551_ _09571_ VGND VGND VPWR VPWR _09572_ sky130_fd_sc_hd__a41o_1
Xwire1173 _01687_ VGND VGND VPWR VPWR net1173 sky130_fd_sc_hd__buf_1
Xwire1184 _01020_ VGND VGND VPWR VPWR net1184 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19431_ net6154 net6140 VGND VGND VPWR VPWR _11268_ sky130_fd_sc_hd__or2b_1
Xwire1195 _10497_ VGND VGND VPWR VPWR net1195 sky130_fd_sc_hd__buf_1
X_16643_ matmul0.matmul_stage_inst.mult2\[3\] VGND VGND VPWR VPWR _08680_ sky130_fd_sc_hd__inv_2
X_13855_ _06053_ _06054_ _06121_ VGND VGND VPWR VPWR _06122_ sky130_fd_sc_hd__a21o_1
XFILLER_0_159_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12806_ _05072_ _05078_ VGND VGND VPWR VPWR _05079_ sky130_fd_sc_hd__xor2_2
X_19362_ _11195_ _11152_ _11188_ VGND VGND VPWR VPWR _11199_ sky130_fd_sc_hd__and3_1
X_16574_ _08547_ _08589_ _08590_ VGND VGND VPWR VPWR _08633_ sky130_fd_sc_hd__o21a_1
X_13786_ net7641 net2332 net2327 VGND VGND VPWR VPWR _06054_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18313_ net7126 _10160_ _10163_ VGND VGND VPWR VPWR _10164_ sky130_fd_sc_hd__a21o_1
X_15525_ net4083 net4081 VGND VGND VPWR VPWR _07598_ sky130_fd_sc_hd__or2_1
X_12737_ _04982_ _05009_ VGND VGND VPWR VPWR _05010_ sky130_fd_sc_hd__xnor2_2
X_19293_ net3884 net3901 _11124_ _11129_ VGND VGND VPWR VPWR _11130_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_84_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18244_ net3956 _10039_ _10094_ VGND VGND VPWR VPWR _10095_ sky130_fd_sc_hd__a21boi_1
X_15456_ _07527_ _07529_ VGND VGND VPWR VPWR _07530_ sky130_fd_sc_hd__xnor2_1
X_12668_ _04916_ _04940_ VGND VGND VPWR VPWR _04941_ sky130_fd_sc_hd__xnor2_2
Xfanout8696 net8702 VGND VGND VPWR VPWR net8696 sky130_fd_sc_hd__buf_1
XFILLER_0_167_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14407_ net4233 VGND VGND VPWR VPWR _06609_ sky130_fd_sc_hd__clkbuf_1
Xwire8780 net8778 VGND VGND VPWR VPWR net8780 sky130_fd_sc_hd__buf_1
XFILLER_0_114_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18175_ _10025_ _09822_ VGND VGND VPWR VPWR _10026_ sky130_fd_sc_hd__nand2_1
Xwire8791 net8790 VGND VGND VPWR VPWR net8791 sky130_fd_sc_hd__buf_1
XFILLER_0_5_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15387_ _07459_ net1116 _07460_ VGND VGND VPWR VPWR _07461_ sky130_fd_sc_hd__o21ai_1
X_12599_ _04878_ VGND VGND VPWR VPWR _00004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17126_ net3344 _08931_ net2593 VGND VGND VPWR VPWR _09081_ sky130_fd_sc_hd__mux2_1
Xwire470 _03566_ VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__clkbuf_1
X_14338_ _06555_ matmul0.a_in\[4\] net902 VGND VGND VPWR VPWR _06556_ sky130_fd_sc_hd__mux2_1
Xwire481 net482 VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__clkbuf_1
Xwire492 _08234_ VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__buf_1
XFILLER_0_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17057_ net7039 _09014_ _09015_ _08994_ VGND VGND VPWR VPWR _09016_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14269_ net62 net2931 net2278 net9060 VGND VGND VPWR VPWR _00042_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16008_ _08016_ net673 VGND VGND VPWR VPWR _08076_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17959_ _09696_ _09604_ VGND VGND VPWR VPWR _09810_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20970_ _00984_ _00985_ VGND VGND VPWR VPWR _00986_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_174_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_189_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19629_ net6178 net6269 VGND VGND VPWR VPWR _11466_ sky130_fd_sc_hd__xnor2_2
Xmax_length6808 net6809 VGND VGND VPWR VPWR net6808 sky130_fd_sc_hd__buf_1
X_22640_ net3114 net3076 VGND VGND VPWR VPWR _02605_ sky130_fd_sc_hd__nand2_1
XFILLER_0_177_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22571_ net9050 net2043 net3093 net3092 VGND VGND VPWR VPWR _00553_ sky130_fd_sc_hd__a22o_1
XFILLER_0_180_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_60_clk clknet_4_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_35_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24310_ _04045_ _04119_ _04168_ _04169_ VGND VGND VPWR VPWR _04170_ sky130_fd_sc_hd__a31o_1
XFILLER_0_75_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21522_ net5971 _01430_ _01534_ VGND VGND VPWR VPWR _01535_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_134_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25290_ clknet_leaf_77_clk _00173_ net8436 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.d\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24241_ _04097_ net852 VGND VGND VPWR VPWR _04102_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21453_ net5807 net5490 VGND VGND VPWR VPWR _01466_ sky130_fd_sc_hd__nand2_1
Xwire6107 net6108 VGND VGND VPWR VPWR net6107 sky130_fd_sc_hd__buf_1
XFILLER_0_17_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6129 net6130 VGND VGND VPWR VPWR net6129 sky130_fd_sc_hd__buf_1
X_20404_ cordic0.slte0.opA\[9\] net1915 _12200_ VGND VGND VPWR VPWR _12202_ sky130_fd_sc_hd__or3_1
XFILLER_0_32_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24172_ _04031_ _04032_ VGND VGND VPWR VPWR _04034_ sky130_fd_sc_hd__or2_1
Xwire5417 net5418 VGND VGND VPWR VPWR net5417 sky130_fd_sc_hd__clkbuf_1
X_21384_ _01276_ net1390 _01397_ VGND VGND VPWR VPWR _01398_ sky130_fd_sc_hd__a21o_1
XFILLER_0_189_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5428 net5429 VGND VGND VPWR VPWR net5428 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5439 net5443 VGND VGND VPWR VPWR net5439 sky130_fd_sc_hd__buf_1
X_23123_ _02991_ _02992_ VGND VGND VPWR VPWR _02993_ sky130_fd_sc_hd__xnor2_2
Xwire4705 net4706 VGND VGND VPWR VPWR net4705 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20335_ net951 _12125_ cordic0.slte0.opA\[3\] VGND VGND VPWR VPWR _12138_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4716 net4717 VGND VGND VPWR VPWR net4716 sky130_fd_sc_hd__buf_1
Xwire4727 net4728 VGND VGND VPWR VPWR net4727 sky130_fd_sc_hd__buf_1
Xwire4738 net4739 VGND VGND VPWR VPWR net4738 sky130_fd_sc_hd__buf_1
Xwire4749 net4750 VGND VGND VPWR VPWR net4749 sky130_fd_sc_hd__buf_1
X_23054_ net4742 net4772 _02923_ VGND VGND VPWR VPWR _02924_ sky130_fd_sc_hd__o21ai_1
X_20266_ net4 _12076_ VGND VGND VPWR VPWR _12077_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22005_ _02010_ _02011_ VGND VGND VPWR VPWR _02013_ sky130_fd_sc_hd__or2_1
Xinput104 pid_d_data[1] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_1
X_20197_ net6042 net6000 _12021_ net6063 net6024 VGND VGND VPWR VPWR _12022_ sky130_fd_sc_hd__o221a_1
Xinput115 pid_q_addr[10] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_1
Xinput126 pid_q_addr[6] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_1
Xinput137 pid_q_data[1] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_1
Xinput148 valid VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_1
Xmax_length8711 net8708 VGND VGND VPWR VPWR net8711 sky130_fd_sc_hd__clkbuf_2
X_23956_ net4488 _03819_ VGND VGND VPWR VPWR _03820_ sky130_fd_sc_hd__nand2_1
Xmax_length8766 net8763 VGND VGND VPWR VPWR net8766 sky130_fd_sc_hd__clkbuf_1
X_22907_ pid_d.out\[10\] net2466 _02799_ net4329 VGND VGND VPWR VPWR _02800_ sky130_fd_sc_hd__a22o_1
X_23887_ net1163 _03647_ _03751_ VGND VGND VPWR VPWR _03752_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length8799 net8800 VGND VGND VPWR VPWR net8799 sky130_fd_sc_hd__clkbuf_1
X_13640_ _05908_ _05909_ VGND VGND VPWR VPWR _05910_ sky130_fd_sc_hd__xnor2_1
X_25626_ clknet_leaf_117_clk _00499_ net8337 VGND VGND VPWR VPWR cordic0.slte0.opA\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22838_ pid_d.out\[3\] net5982 VGND VGND VPWR VPWR _02738_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_195_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13571_ _05840_ _05841_ VGND VGND VPWR VPWR _05842_ sky130_fd_sc_hd__or2b_1
XFILLER_0_137_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25557_ clknet_leaf_117_clk _00430_ net8332 VGND VGND VPWR VPWR cordic0.gm0.iter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22769_ pid_d.ki\[14\] _02690_ net2039 VGND VGND VPWR VPWR _02691_ sky130_fd_sc_hd__mux2_1
Xwire8010 net8011 VGND VGND VPWR VPWR net8010 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_51_clk clknet_4_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_52_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8021 pid_q.target\[3\] VGND VGND VPWR VPWR net8021 sky130_fd_sc_hd__clkbuf_1
X_15310_ _07382_ _07383_ VGND VGND VPWR VPWR _07384_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_186_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8032 net8033 VGND VGND VPWR VPWR net8032 sky130_fd_sc_hd__clkbuf_1
X_24508_ _04355_ _04364_ VGND VGND VPWR VPWR _04365_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16290_ _08249_ net1251 net1508 VGND VGND VPWR VPWR _08354_ sky130_fd_sc_hd__a21bo_1
X_25488_ clknet_leaf_48_clk _00368_ net8761 VGND VGND VPWR VPWR svm0.tA\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8043 net8044 VGND VGND VPWR VPWR net8043 sky130_fd_sc_hd__buf_1
Xfanout6524 net6529 VGND VGND VPWR VPWR net6524 sky130_fd_sc_hd__clkbuf_1
Xwire8065 net8066 VGND VGND VPWR VPWR net8065 sky130_fd_sc_hd__clkbuf_1
Xwire7320 net7321 VGND VGND VPWR VPWR net7320 sky130_fd_sc_hd__buf_1
Xwire8076 net8077 VGND VGND VPWR VPWR net8076 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15241_ _07302_ _07314_ VGND VGND VPWR VPWR _07315_ sky130_fd_sc_hd__xnor2_2
Xfanout6535 net6545 VGND VGND VPWR VPWR net6535 sky130_fd_sc_hd__buf_1
Xwire7331 net7332 VGND VGND VPWR VPWR net7331 sky130_fd_sc_hd__clkbuf_1
Xwire8087 net8088 VGND VGND VPWR VPWR net8087 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24439_ _04296_ net4918 net4896 _04287_ VGND VGND VPWR VPWR _04297_ sky130_fd_sc_hd__a211o_1
Xwire7342 net7351 VGND VGND VPWR VPWR net7342 sky130_fd_sc_hd__clkbuf_1
Xwire7353 net7354 VGND VGND VPWR VPWR net7353 sky130_fd_sc_hd__buf_1
Xwire8098 net95 VGND VGND VPWR VPWR net8098 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7364 net7365 VGND VGND VPWR VPWR net7364 sky130_fd_sc_hd__buf_1
Xwire6630 net6631 VGND VGND VPWR VPWR net6630 sky130_fd_sc_hd__buf_1
X_15172_ net3576 net3572 net4213 net4211 VGND VGND VPWR VPWR _07246_ sky130_fd_sc_hd__o22a_1
Xwire7386 net7387 VGND VGND VPWR VPWR net7386 sky130_fd_sc_hd__clkbuf_1
Xwire6652 net6653 VGND VGND VPWR VPWR net6652 sky130_fd_sc_hd__clkbuf_1
Xfanout5856 net5864 VGND VGND VPWR VPWR net5856 sky130_fd_sc_hd__buf_1
Xmax_length3084 net3085 VGND VGND VPWR VPWR net3084 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2350 net2351 VGND VGND VPWR VPWR net2350 sky130_fd_sc_hd__buf_1
XFILLER_0_50_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5867 net5875 VGND VGND VPWR VPWR net5867 sky130_fd_sc_hd__buf_1
X_14123_ _06340_ VGND VGND VPWR VPWR _06385_ sky130_fd_sc_hd__inv_2
Xwire6674 net6675 VGND VGND VPWR VPWR net6674 sky130_fd_sc_hd__clkbuf_1
Xfanout5878 net5885 VGND VGND VPWR VPWR net5878 sky130_fd_sc_hd__buf_1
X_19980_ _11764_ _11810_ VGND VGND VPWR VPWR _11811_ sky130_fd_sc_hd__xnor2_1
Xwire5940 net5936 VGND VGND VPWR VPWR net5940 sky130_fd_sc_hd__buf_1
Xwire6696 svm0.counter\[13\] VGND VGND VPWR VPWR net6696 sky130_fd_sc_hd__clkbuf_1
Xmax_length2383 net2384 VGND VGND VPWR VPWR net2383 sky130_fd_sc_hd__clkbuf_1
Xwire5951 net5952 VGND VGND VPWR VPWR net5951 sky130_fd_sc_hd__buf_1
XFILLER_0_162_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5973 pid_d.curr_error\[0\] VGND VGND VPWR VPWR net5973 sky130_fd_sc_hd__clkbuf_2
X_18931_ _06500_ VGND VGND VPWR VPWR _10770_ sky130_fd_sc_hd__buf_1
Xwire5984 net5985 VGND VGND VPWR VPWR net5984 sky130_fd_sc_hd__clkbuf_2
X_14054_ _06316_ _06317_ VGND VGND VPWR VPWR _06318_ sky130_fd_sc_hd__nor2_1
Xwire5995 net5996 VGND VGND VPWR VPWR net5995 sky130_fd_sc_hd__buf_1
X_13005_ _05264_ _05277_ VGND VGND VPWR VPWR _05278_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18862_ _10703_ _10680_ net1428 VGND VGND VPWR VPWR _10704_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17813_ net6974 net6925 VGND VGND VPWR VPWR _09664_ sky130_fd_sc_hd__nand2_1
X_18793_ _10582_ _10583_ net3983 VGND VGND VPWR VPWR _10637_ sky130_fd_sc_hd__mux2_1
X_17744_ net5370 _06525_ _09596_ net6443 VGND VGND VPWR VPWR _00437_ sky130_fd_sc_hd__a22o_1
X_14956_ net6559 net6587 matmul0.matmul_stage_inst.e\[7\] VGND VGND VPWR VPWR _07030_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_178_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13907_ net3686 net2968 VGND VGND VPWR VPWR _06173_ sky130_fd_sc_hd__nand2_1
X_17675_ svm0.tA\[3\] _09554_ _09243_ VGND VGND VPWR VPWR _09555_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14887_ _06961_ VGND VGND VPWR VPWR _00214_ sky130_fd_sc_hd__clkbuf_1
X_19414_ _11103_ _11244_ _11247_ _11249_ _11250_ VGND VGND VPWR VPWR _11251_ sky130_fd_sc_hd__o32a_1
X_16626_ matmul0.matmul_stage_inst.mult2\[1\] matmul0.matmul_stage_inst.mult1\[1\]
+ VGND VGND VPWR VPWR _08665_ sky130_fd_sc_hd__nand2_1
X_13838_ _06096_ _06104_ VGND VGND VPWR VPWR _06105_ sky130_fd_sc_hd__xnor2_2
X_19345_ _10803_ _11181_ VGND VGND VPWR VPWR _11182_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16557_ _08612_ net1242 VGND VGND VPWR VPWR _08616_ sky130_fd_sc_hd__xnor2_1
X_13769_ net7700 net1943 net2292 VGND VGND VPWR VPWR _06037_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_42_clk clknet_4_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_57_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15508_ net2677 _07580_ VGND VGND VPWR VPWR _07581_ sky130_fd_sc_hd__xnor2_1
X_19276_ _10909_ _11112_ net872 VGND VGND VPWR VPWR _11113_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16488_ _08501_ _08537_ _08538_ VGND VGND VPWR VPWR _08548_ sky130_fd_sc_hd__a21o_1
Xfanout8471 net8476 VGND VGND VPWR VPWR net8471 sky130_fd_sc_hd__buf_1
XFILLER_0_127_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18227_ net7094 _10077_ _09809_ VGND VGND VPWR VPWR _10078_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15439_ _07372_ _07373_ _07512_ VGND VGND VPWR VPWR _07513_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18158_ _10003_ _10005_ net1212 VGND VGND VPWR VPWR _10009_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17109_ net1818 _09065_ net8049 VGND VGND VPWR VPWR _09066_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18089_ net2548 _09939_ VGND VGND VPWR VPWR _09940_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_159_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20120_ _11946_ _11947_ VGND VGND VPWR VPWR _11948_ sky130_fd_sc_hd__and2_1
Xclkbuf_4_3__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_4_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20051_ net6077 _11490_ VGND VGND VPWR VPWR _11880_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1909 _06846_ VGND VGND VPWR VPWR net1909 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23810_ _03673_ _03674_ VGND VGND VPWR VPWR _03675_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_175_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24790_ _04614_ _04615_ VGND VGND VPWR VPWR _04616_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_178_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23741_ net5120 net3744 _03606_ VGND VGND VPWR VPWR _03607_ sky130_fd_sc_hd__a21o_1
X_20953_ net5635 net5613 net5797 VGND VGND VPWR VPWR _00969_ sky130_fd_sc_hd__and3b_1
Xmax_length7328 matmul0.alpha_pass\[4\] VGND VGND VPWR VPWR net7328 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23672_ _03537_ _03538_ VGND VGND VPWR VPWR _03539_ sky130_fd_sc_hd__or2b_1
X_20884_ _00896_ _00899_ VGND VGND VPWR VPWR _00900_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_177_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25411_ clknet_leaf_80_clk _00294_ net8494 VGND VGND VPWR VPWR matmul0.a\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_192_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22623_ net7203 _02590_ VGND VGND VPWR VPWR _02593_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_33_clk clknet_4_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_193_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22554_ net8988 net2049 _02539_ VGND VGND VPWR VPWR _00549_ sky130_fd_sc_hd__a21o_1
X_25342_ clknet_leaf_83_clk _00225_ net8714 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21505_ _01515_ net947 VGND VGND VPWR VPWR _01518_ sky130_fd_sc_hd__xor2_1
XFILLER_0_133_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22485_ net5671 _02354_ _02482_ _02483_ _02485_ VGND VGND VPWR VPWR _02486_ sky130_fd_sc_hd__a32o_1
XFILLER_0_134_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25273_ clknet_leaf_93_clk _00156_ net8449 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.c\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24224_ _04081_ _04084_ VGND VGND VPWR VPWR _04085_ sky130_fd_sc_hd__xnor2_1
X_21436_ net5685 net5608 VGND VGND VPWR VPWR _01449_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_15_Left_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5214 net5215 VGND VGND VPWR VPWR net5214 sky130_fd_sc_hd__buf_1
Xwire5225 net5226 VGND VGND VPWR VPWR net5225 sky130_fd_sc_hd__clkbuf_1
X_24155_ _03922_ _03931_ VGND VGND VPWR VPWR _04017_ sky130_fd_sc_hd__nor2_1
Xwire5236 net5237 VGND VGND VPWR VPWR net5236 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4502 net4498 VGND VGND VPWR VPWR net4502 sky130_fd_sc_hd__buf_1
Xwire5247 net5248 VGND VGND VPWR VPWR net5247 sky130_fd_sc_hd__clkbuf_2
X_21367_ net5416 net5922 VGND VGND VPWR VPWR _01381_ sky130_fd_sc_hd__nand2_1
Xwire4513 net4507 VGND VGND VPWR VPWR net4513 sky130_fd_sc_hd__buf_1
XFILLER_0_31_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5258 matmul0.beta_pass\[7\] VGND VGND VPWR VPWR net5258 sky130_fd_sc_hd__clkbuf_1
Xwire4524 net4517 VGND VGND VPWR VPWR net4524 sky130_fd_sc_hd__buf_1
Xwire5269 net5270 VGND VGND VPWR VPWR net5269 sky130_fd_sc_hd__buf_1
XFILLER_0_43_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23106_ _02974_ _02975_ VGND VGND VPWR VPWR _02976_ sky130_fd_sc_hd__nand2_1
Xwire4535 net4536 VGND VGND VPWR VPWR net4535 sky130_fd_sc_hd__buf_1
X_20318_ net4037 _12098_ _12120_ _12121_ net6459 VGND VGND VPWR VPWR _12122_ sky130_fd_sc_hd__a221oi_1
Xwire4546 net4547 VGND VGND VPWR VPWR net4546 sky130_fd_sc_hd__buf_1
X_24086_ pid_q.prev_error\[7\] pid_q.curr_error\[7\] VGND VGND VPWR VPWR _03949_ sky130_fd_sc_hd__xnor2_1
Xwire3801 net3802 VGND VGND VPWR VPWR net3801 sky130_fd_sc_hd__clkbuf_1
Xwire4557 net4558 VGND VGND VPWR VPWR net4557 sky130_fd_sc_hd__clkbuf_1
X_21298_ _01304_ _01312_ VGND VGND VPWR VPWR _01313_ sky130_fd_sc_hd__xnor2_2
Xwire3812 net3813 VGND VGND VPWR VPWR net3812 sky130_fd_sc_hd__buf_1
Xwire3823 net3824 VGND VGND VPWR VPWR net3823 sky130_fd_sc_hd__clkbuf_2
Xwire4579 net4580 VGND VGND VPWR VPWR net4579 sky130_fd_sc_hd__buf_1
Xwire3834 net3835 VGND VGND VPWR VPWR net3834 sky130_fd_sc_hd__clkbuf_1
X_23037_ _02905_ _02906_ VGND VGND VPWR VPWR _02907_ sky130_fd_sc_hd__nand2_1
Xwire3845 _12298_ VGND VGND VPWR VPWR net3845 sky130_fd_sc_hd__clkbuf_1
X_20249_ _12063_ cordic0.slte0.opB\[10\] net2532 VGND VGND VPWR VPWR _12064_ sky130_fd_sc_hd__mux2_1
Xwire3856 _11559_ VGND VGND VPWR VPWR net3856 sky130_fd_sc_hd__buf_2
Xwire3867 net3868 VGND VGND VPWR VPWR net3867 sky130_fd_sc_hd__clkbuf_1
Xwire3878 net3879 VGND VGND VPWR VPWR net3878 sky130_fd_sc_hd__buf_1
Xwire3889 _10882_ VGND VGND VPWR VPWR net3889 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14810_ net7442 net7170 net3628 VGND VGND VPWR VPWR _06922_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_24_Left_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15790_ net987 _07859_ VGND VGND VPWR VPWR _07860_ sky130_fd_sc_hd__xnor2_1
X_24988_ pid_q.kp\[13\] _04728_ _04734_ VGND VGND VPWR VPWR _04749_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14741_ _06873_ _06874_ net7448 VGND VGND VPWR VPWR _06875_ sky130_fd_sc_hd__o21ai_1
X_23939_ _03795_ _03802_ VGND VGND VPWR VPWR _03803_ sky130_fd_sc_hd__xnor2_1
Xmax_length8563 net8561 VGND VGND VPWR VPWR net8563 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_58_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17460_ _09281_ _09349_ _09353_ VGND VGND VPWR VPWR _09354_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_98_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14672_ _06817_ net3620 VGND VGND VPWR VPWR _06824_ sky130_fd_sc_hd__nor2_1
Xmax_length7884 net7885 VGND VGND VPWR VPWR net7884 sky130_fd_sc_hd__clkbuf_1
X_16411_ net1507 _08472_ VGND VGND VPWR VPWR _08473_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_2_3_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3_0_clk sky130_fd_sc_hd__clkbuf_8
X_13623_ _05889_ _05891_ net911 VGND VGND VPWR VPWR _05893_ sky130_fd_sc_hd__a21o_1
X_25609_ clknet_leaf_105_clk _00482_ net8356 VGND VGND VPWR VPWR cordic0.domain\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_17391_ _09295_ net614 _09296_ _09298_ VGND VGND VPWR VPWR _00381_ sky130_fd_sc_hd__a31o_1
XFILLER_0_55_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_24_clk clknet_4_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_16
X_19130_ net3216 _10808_ net3215 VGND VGND VPWR VPWR _10967_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_66_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16342_ _08402_ _08404_ VGND VGND VPWR VPWR _08405_ sky130_fd_sc_hd__and2_1
X_13554_ net7655 net1982 net2360 VGND VGND VPWR VPWR _05825_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19061_ net6352 VGND VGND VPWR VPWR _10898_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_33_Left_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout7066 net7077 VGND VGND VPWR VPWR net7066 sky130_fd_sc_hd__buf_1
X_16273_ _08276_ _08281_ _08336_ VGND VGND VPWR VPWR _08337_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_180_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13485_ _05743_ _05757_ VGND VGND VPWR VPWR _05758_ sky130_fd_sc_hd__xnor2_1
X_18012_ net7082 _09617_ VGND VGND VPWR VPWR _09863_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout5620 pid_d.mult0.a\[2\] VGND VGND VPWR VPWR net5620 sky130_fd_sc_hd__buf_1
X_15224_ _07278_ _07280_ _07295_ _07297_ VGND VGND VPWR VPWR _07298_ sky130_fd_sc_hd__a22o_1
Xwire7161 matmul0.sin\[1\] VGND VGND VPWR VPWR net7161 sky130_fd_sc_hd__buf_1
Xwire7172 net7173 VGND VGND VPWR VPWR net7172 sky130_fd_sc_hd__buf_1
Xwire7183 matmul0.a\[0\] VGND VGND VPWR VPWR net7183 sky130_fd_sc_hd__clkbuf_1
Xwire7194 net7195 VGND VGND VPWR VPWR net7194 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire6471 net6472 VGND VGND VPWR VPWR net6471 sky130_fd_sc_hd__buf_1
X_15155_ _07227_ _07228_ VGND VGND VPWR VPWR _07229_ sky130_fd_sc_hd__xor2_2
XFILLER_0_50_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6482 net6481 VGND VGND VPWR VPWR net6482 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_196_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6493 net6495 VGND VGND VPWR VPWR net6493 sky130_fd_sc_hd__buf_1
XFILLER_0_1_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14106_ _06323_ _06352_ _06367_ VGND VGND VPWR VPWR _06368_ sky130_fd_sc_hd__a21oi_4
Xwire5770 net5771 VGND VGND VPWR VPWR net5770 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5781 net5782 VGND VGND VPWR VPWR net5781 sky130_fd_sc_hd__clkbuf_1
X_19963_ net6094 _11755_ _11758_ VGND VGND VPWR VPWR _11794_ sky130_fd_sc_hd__nor3_1
X_15086_ net2790 _07154_ _07155_ _07147_ _07159_ VGND VGND VPWR VPWR _07160_ sky130_fd_sc_hd__o32a_1
Xfanout4996 net5008 VGND VGND VPWR VPWR net4996 sky130_fd_sc_hd__buf_1
XFILLER_0_38_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14037_ net7663 net2955 net3674 VGND VGND VPWR VPWR _06301_ sky130_fd_sc_hd__and3_1
X_18914_ net6828 net6876 VGND VGND VPWR VPWR _10754_ sky130_fd_sc_hd__nor2_1
X_19894_ _11667_ _11716_ _11720_ _11723_ _11726_ VGND VGND VPWR VPWR _11727_ sky130_fd_sc_hd__o32a_1
X_18845_ _10629_ _10647_ VGND VGND VPWR VPWR _10688_ sky130_fd_sc_hd__nor2_1
XFILLER_0_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18776_ _10601_ _10602_ net764 VGND VGND VPWR VPWR _10620_ sky130_fd_sc_hd__a21bo_1
X_15988_ net3449 _07838_ VGND VGND VPWR VPWR _08056_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17727_ _09586_ VGND VGND VPWR VPWR _00430_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_4_11__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_4_11__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_14939_ net6619 net6644 net7384 VGND VGND VPWR VPWR _07013_ sky130_fd_sc_hd__o21a_1
XFILLER_0_145_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17658_ _09534_ _09535_ _09536_ _09537_ VGND VGND VPWR VPWR _09538_ sky130_fd_sc_hd__and4b_1
XFILLER_0_159_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16609_ _08654_ VGND VGND VPWR VPWR _00243_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17589_ net2154 net1794 net1460 net820 VGND VGND VPWR VPWR _09471_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_15_clk clknet_4_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_18_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19328_ net6263 _11163_ net3871 VGND VGND VPWR VPWR _11165_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19259_ _10869_ _11095_ VGND VGND VPWR VPWR _11096_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22270_ net381 _02273_ VGND VGND VPWR VPWR _02274_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold100 pid_q.target\[6\] VGND VGND VPWR VPWR net9053 sky130_fd_sc_hd__dlygate4sd3_1
X_21221_ _00938_ _00968_ VGND VGND VPWR VPWR _01237_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold111 cordic0.sin\[6\] VGND VGND VPWR VPWR net9064 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 cordic0.sin\[4\] VGND VGND VPWR VPWR net9075 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 matmul0.op_in\[1\] VGND VGND VPWR VPWR net9086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 svm0.vC\[15\] VGND VGND VPWR VPWR net9097 sky130_fd_sc_hd__dlygate4sd3_1
X_21152_ net5618 net5937 VGND VGND VPWR VPWR _01168_ sky130_fd_sc_hd__nand2_1
Xhold155 svm0.tA\[1\] VGND VGND VPWR VPWR net9108 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3108 net3109 VGND VGND VPWR VPWR net3108 sky130_fd_sc_hd__buf_1
Xwire3119 net3120 VGND VGND VPWR VPWR net3119 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold166 pid_d.prev_error\[8\] VGND VGND VPWR VPWR net9119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 matmul0.matmul_stage_inst.b\[11\] VGND VGND VPWR VPWR net9130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 svm0.tB\[12\] VGND VGND VPWR VPWR net9141 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20103_ _11928_ _11920_ _11930_ VGND VGND VPWR VPWR _11931_ sky130_fd_sc_hd__o21ai_1
Xhold199 svm0.tC\[0\] VGND VGND VPWR VPWR net9152 sky130_fd_sc_hd__dlygate4sd3_1
X_21083_ net5879 _01097_ _01098_ VGND VGND VPWR VPWR _01099_ sky130_fd_sc_hd__a21bo_1
Xwire2418 net2419 VGND VGND VPWR VPWR net2418 sky130_fd_sc_hd__clkbuf_1
Xwire2429 _03205_ VGND VGND VPWR VPWR net2429 sky130_fd_sc_hd__buf_1
X_24911_ net3730 net2011 _04700_ net114 VGND VGND VPWR VPWR _04701_ sky130_fd_sc_hd__a22o_1
XFILLER_0_186_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20034_ net6013 net6028 VGND VGND VPWR VPWR _11864_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1706 net1707 VGND VGND VPWR VPWR net1706 sky130_fd_sc_hd__clkbuf_2
X_25891_ clknet_leaf_16_clk _00764_ net8622 VGND VGND VPWR VPWR pid_q.kp\[3\] sky130_fd_sc_hd__dfrtp_1
Xwire1717 _01887_ VGND VGND VPWR VPWR net1717 sky130_fd_sc_hd__buf_1
Xwire1728 _01388_ VGND VGND VPWR VPWR net1728 sky130_fd_sc_hd__buf_1
Xwire1739 _12408_ VGND VGND VPWR VPWR net1739 sky130_fd_sc_hd__buf_1
X_24842_ net7479 net457 _04184_ VGND VGND VPWR VPWR _04654_ sky130_fd_sc_hd__a21oi_1
X_24773_ _04599_ _04600_ net1988 VGND VGND VPWR VPWR _04601_ sky130_fd_sc_hd__o21ai_1
X_21985_ net2068 _01885_ VGND VGND VPWR VPWR _01993_ sky130_fd_sc_hd__nand2_1
X_23724_ net4562 net4997 VGND VGND VPWR VPWR _03590_ sky130_fd_sc_hd__nand2_1
Xmax_length7147 net7143 VGND VGND VPWR VPWR net7147 sky130_fd_sc_hd__buf_1
X_20936_ _00949_ _00951_ VGND VGND VPWR VPWR _00952_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23655_ _03520_ _03521_ VGND VGND VPWR VPWR _03522_ sky130_fd_sc_hd__xnor2_2
X_20867_ net5627 net5775 VGND VGND VPWR VPWR _00883_ sky130_fd_sc_hd__nand2_1
XFILLER_0_194_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22606_ net7250 _02576_ VGND VGND VPWR VPWR _02580_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23586_ _03357_ _03358_ _03359_ VGND VGND VPWR VPWR _03454_ sky130_fd_sc_hd__o21a_1
XFILLER_0_107_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20798_ _12541_ _12546_ _00813_ VGND VGND VPWR VPWR _00814_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_153_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25325_ clknet_leaf_79_clk _00208_ net8491 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.f\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22537_ net5968 net2381 net2047 VGND VGND VPWR VPWR _02531_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13270_ _05441_ _05444_ VGND VGND VPWR VPWR _05543_ sky130_fd_sc_hd__xor2_1
XFILLER_0_63_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25256_ clknet_leaf_71_clk _00139_ net8457 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.b\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_22468_ _02344_ _02446_ net1169 VGND VGND VPWR VPWR _02469_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5000 net5001 VGND VGND VPWR VPWR net5000 sky130_fd_sc_hd__buf_1
Xwire5022 net5023 VGND VGND VPWR VPWR net5022 sky130_fd_sc_hd__buf_1
X_24207_ net3040 _03973_ _03968_ VGND VGND VPWR VPWR _04068_ sky130_fd_sc_hd__a21bo_1
Xwire5033 net5034 VGND VGND VPWR VPWR net5033 sky130_fd_sc_hd__clkbuf_1
X_21419_ _01428_ _01429_ _01431_ VGND VGND VPWR VPWR _01433_ sky130_fd_sc_hd__and3_1
X_22399_ pid_d.prev_error\[13\] net5965 _02262_ _02391_ VGND VGND VPWR VPWR _02401_
+ sky130_fd_sc_hd__a2bb2o_1
X_25187_ clknet_leaf_63_clk _00076_ net8667 VGND VGND VPWR VPWR matmul0.a_in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire5044 net5045 VGND VGND VPWR VPWR net5044 sky130_fd_sc_hd__clkbuf_1
Xwire5055 net5043 VGND VGND VPWR VPWR net5055 sky130_fd_sc_hd__clkbuf_1
Xwire4310 _04862_ VGND VGND VPWR VPWR net4310 sky130_fd_sc_hd__buf_1
Xwire5066 net5061 VGND VGND VPWR VPWR net5066 sky130_fd_sc_hd__buf_1
Xwire4321 net4322 VGND VGND VPWR VPWR net4321 sky130_fd_sc_hd__clkbuf_1
Xwire5077 net5078 VGND VGND VPWR VPWR net5077 sky130_fd_sc_hd__buf_1
X_24138_ _03998_ _03999_ VGND VGND VPWR VPWR _04000_ sky130_fd_sc_hd__and2b_1
Xwire4332 net4333 VGND VGND VPWR VPWR net4332 sky130_fd_sc_hd__clkbuf_1
Xwire4343 net4344 VGND VGND VPWR VPWR net4343 sky130_fd_sc_hd__clkbuf_1
Xwire5088 net5089 VGND VGND VPWR VPWR net5088 sky130_fd_sc_hd__buf_1
Xwire5099 net5100 VGND VGND VPWR VPWR net5099 sky130_fd_sc_hd__buf_1
Xwire4354 net4355 VGND VGND VPWR VPWR net4354 sky130_fd_sc_hd__buf_1
Xwire4365 net4366 VGND VGND VPWR VPWR net4365 sky130_fd_sc_hd__buf_1
Xwire3620 net3621 VGND VGND VPWR VPWR net3620 sky130_fd_sc_hd__buf_1
Xwire4376 net4377 VGND VGND VPWR VPWR net4376 sky130_fd_sc_hd__clkbuf_1
Xwire3631 net3632 VGND VGND VPWR VPWR net3631 sky130_fd_sc_hd__buf_1
X_16960_ net7129 net2177 _08919_ _08922_ _08838_ VGND VGND VPWR VPWR _08923_ sky130_fd_sc_hd__a32o_1
X_24069_ _03922_ _03931_ VGND VGND VPWR VPWR _03932_ sky130_fd_sc_hd__nand2_1
Xwire4387 net4388 VGND VGND VPWR VPWR net4387 sky130_fd_sc_hd__clkbuf_1
Xwire3653 net3654 VGND VGND VPWR VPWR net3653 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4398 net4399 VGND VGND VPWR VPWR net4398 sky130_fd_sc_hd__clkbuf_1
Xwire3664 net3665 VGND VGND VPWR VPWR net3664 sky130_fd_sc_hd__clkbuf_1
Xwire2930 _06514_ VGND VGND VPWR VPWR net2930 sky130_fd_sc_hd__buf_1
X_15911_ _07852_ _07854_ _07850_ VGND VGND VPWR VPWR _07980_ sky130_fd_sc_hd__o21a_1
Xwire3675 _05616_ VGND VGND VPWR VPWR net3675 sky130_fd_sc_hd__buf_1
Xwire3686 net3687 VGND VGND VPWR VPWR net3686 sky130_fd_sc_hd__buf_1
XFILLER_0_21_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16891_ _08852_ _08853_ _08854_ VGND VGND VPWR VPWR _08855_ sky130_fd_sc_hd__a21oi_1
Xwire2941 _06501_ VGND VGND VPWR VPWR net2941 sky130_fd_sc_hd__clkbuf_1
Xwire2952 net2953 VGND VGND VPWR VPWR net2952 sky130_fd_sc_hd__clkbuf_1
Xwire3697 _04884_ VGND VGND VPWR VPWR net3697 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_188_Right_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2963 _05285_ VGND VGND VPWR VPWR net2963 sky130_fd_sc_hd__buf_1
XFILLER_0_194_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18630_ net2131 _10476_ VGND VGND VPWR VPWR _10477_ sky130_fd_sc_hd__xnor2_1
X_15842_ _07804_ _07815_ _07813_ VGND VGND VPWR VPWR _07912_ sky130_fd_sc_hd__o21a_1
Xwire2985 net2986 VGND VGND VPWR VPWR net2985 sky130_fd_sc_hd__clkbuf_1
Xwire2996 net2997 VGND VGND VPWR VPWR net2996 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18561_ _10384_ net1436 _10408_ VGND VGND VPWR VPWR _10409_ sky130_fd_sc_hd__o21ba_1
X_15773_ net3396 VGND VGND VPWR VPWR _07843_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12985_ net7715 net2344 net2341 VGND VGND VPWR VPWR _05258_ sky130_fd_sc_hd__and3_1
X_17512_ net3271 net2571 _09396_ _09398_ VGND VGND VPWR VPWR _00402_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14724_ net3613 net7148 _06860_ VGND VGND VPWR VPWR _06863_ sky130_fd_sc_hd__a21o_1
X_18492_ _06500_ net1787 VGND VGND VPWR VPWR _10342_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17443_ _09337_ _09338_ _09339_ VGND VGND VPWR VPWR _09340_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14655_ net7439 net7170 net2874 VGND VGND VPWR VPWR _06812_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13606_ net7746 net1942 net2291 VGND VGND VPWR VPWR _05876_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17374_ svm0.delta\[3\] _09283_ _09284_ VGND VGND VPWR VPWR _09285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14586_ net7233 net5207 VGND VGND VPWR VPWR _06761_ sky130_fd_sc_hd__nor2_1
X_19113_ _10947_ _10948_ net3189 _10945_ VGND VGND VPWR VPWR _10950_ sky130_fd_sc_hd__a211o_1
X_16325_ net2783 net3402 VGND VGND VPWR VPWR _08388_ sky130_fd_sc_hd__nand2_1
X_13537_ _05743_ _05757_ _05807_ VGND VGND VPWR VPWR _05808_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19044_ net6296 net3891 _10880_ VGND VGND VPWR VPWR _10881_ sky130_fd_sc_hd__a21oi_1
Xfanout6151 net6160 VGND VGND VPWR VPWR net6151 sky130_fd_sc_hd__clkbuf_2
X_16256_ net2746 net3415 VGND VGND VPWR VPWR _08320_ sky130_fd_sc_hd__nor2_1
X_13468_ net998 _05740_ VGND VGND VPWR VPWR _05741_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15207_ net3462 net3529 VGND VGND VPWR VPWR _07281_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16187_ _08196_ _08250_ _08251_ VGND VGND VPWR VPWR _08252_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13399_ _05663_ net581 _05661_ net583 VGND VGND VPWR VPWR _05672_ sky130_fd_sc_hd__or4b_1
XFILLER_0_3_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15138_ net1889 _07211_ VGND VGND VPWR VPWR _07212_ sky130_fd_sc_hd__or2b_1
XFILLER_0_26_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout4771 net4780 VGND VGND VPWR VPWR net4771 sky130_fd_sc_hd__dlymetal6s2s_1
X_19946_ _11774_ _11776_ VGND VGND VPWR VPWR _11778_ sky130_fd_sc_hd__or2_1
X_15069_ net6622 net6639 net7383 VGND VGND VPWR VPWR _07143_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_4_clk clknet_4_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_156_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19877_ _11709_ VGND VGND VPWR VPWR _11710_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_155_Right_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18828_ _10668_ _10670_ net6921 VGND VGND VPWR VPWR _10671_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_156_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18759_ net421 _10565_ VGND VGND VPWR VPWR _10604_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21770_ _01779_ _01695_ _01696_ VGND VGND VPWR VPWR _01780_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_194_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20721_ _08915_ _12482_ _12492_ VGND VGND VPWR VPWR _12493_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length5019 net5020 VGND VGND VPWR VPWR net5019 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8609 net8608 VGND VGND VPWR VPWR net8609 sky130_fd_sc_hd__buf_1
X_23440_ _03308_ _03309_ VGND VGND VPWR VPWR _03310_ sky130_fd_sc_hd__nor2_1
X_20652_ net1077 _12429_ VGND VGND VPWR VPWR _12430_ sky130_fd_sc_hd__nand2_1
XFILLER_0_175_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7908 net7909 VGND VGND VPWR VPWR net7908 sky130_fd_sc_hd__buf_1
X_23371_ net4863 net4741 VGND VGND VPWR VPWR _03241_ sky130_fd_sc_hd__nand2_1
Xwire7919 net7920 VGND VGND VPWR VPWR net7919 sky130_fd_sc_hd__buf_1
X_20583_ net1740 VGND VGND VPWR VPWR _12366_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25110_ _04851_ VGND VGND VPWR VPWR _04852_ sky130_fd_sc_hd__clkbuf_2
X_22322_ _02324_ _02325_ VGND VGND VPWR VPWR _02326_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25041_ pid_q.out\[6\] net1995 _04791_ VGND VGND VPWR VPWR _04793_ sky130_fd_sc_hd__nor3_1
X_22253_ _02256_ _02257_ VGND VGND VPWR VPWR _02258_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21204_ net808 _01078_ VGND VGND VPWR VPWR _01220_ sky130_fd_sc_hd__and2_1
X_22184_ _02159_ _02188_ VGND VGND VPWR VPWR _02189_ sky130_fd_sc_hd__nand2_1
X_21135_ net5603 net5932 VGND VGND VPWR VPWR _01151_ sky130_fd_sc_hd__nand2_2
Xwire2204 _08258_ VGND VGND VPWR VPWR net2204 sky130_fd_sc_hd__clkbuf_2
Xwire2215 _07898_ VGND VGND VPWR VPWR net2215 sky130_fd_sc_hd__buf_1
Xwire2226 _07788_ VGND VGND VPWR VPWR net2226 sky130_fd_sc_hd__clkbuf_1
X_21066_ _01080_ _01081_ VGND VGND VPWR VPWR _01082_ sky130_fd_sc_hd__xor2_1
Xwire1503 net1504 VGND VGND VPWR VPWR net1503 sky130_fd_sc_hd__clkbuf_1
Xwire2259 _06875_ VGND VGND VPWR VPWR net2259 sky130_fd_sc_hd__clkbuf_1
X_20017_ _11788_ _11810_ _11764_ VGND VGND VPWR VPWR _11847_ sky130_fd_sc_hd__a21bo_1
Xwire1525 net1526 VGND VGND VPWR VPWR net1525 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_122_Right_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1536 _07751_ VGND VGND VPWR VPWR net1536 sky130_fd_sc_hd__buf_1
X_25874_ clknet_leaf_14_clk _00747_ net8621 VGND VGND VPWR VPWR pid_q.ki\[2\] sky130_fd_sc_hd__dfrtp_1
Xwire1547 _06849_ VGND VGND VPWR VPWR net1547 sky130_fd_sc_hd__clkbuf_1
Xwire1558 net1559 VGND VGND VPWR VPWR net1558 sky130_fd_sc_hd__buf_1
Xwire1569 net1570 VGND VGND VPWR VPWR net1569 sky130_fd_sc_hd__clkbuf_1
X_24825_ net5117 _04642_ net2000 net927 VGND VGND VPWR VPWR _00714_ sky130_fd_sc_hd__a22o_1
X_24756_ _04580_ _04581_ net7996 VGND VGND VPWR VPWR _04586_ sky130_fd_sc_hd__a21o_1
X_12770_ _05039_ _05042_ VGND VGND VPWR VPWR _05043_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_90_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21968_ net2065 _01876_ VGND VGND VPWR VPWR _01976_ sky130_fd_sc_hd__nand2_1
Xmax_length6221 net6222 VGND VGND VPWR VPWR net6221 sky130_fd_sc_hd__clkbuf_1
X_23707_ _03571_ _03572_ VGND VGND VPWR VPWR _03574_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20919_ _00877_ _00934_ VGND VGND VPWR VPWR _00935_ sky130_fd_sc_hd__xnor2_1
X_24687_ pid_q.curr_error\[15\] net3020 net1646 VGND VGND VPWR VPWR _04526_ sky130_fd_sc_hd__and3_1
Xmax_length6265 net6266 VGND VGND VPWR VPWR net6265 sky130_fd_sc_hd__buf_1
X_21899_ net5968 VGND VGND VPWR VPWR _01908_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length6276 net6275 VGND VGND VPWR VPWR net6276 sky130_fd_sc_hd__buf_1
X_14440_ net8186 net3631 VGND VGND VPWR VPWR _06634_ sky130_fd_sc_hd__and2_1
X_23638_ _03417_ _03419_ _03504_ VGND VGND VPWR VPWR _03505_ sky130_fd_sc_hd__o21ai_1
Xmax_length6287 net6289 VGND VGND VPWR VPWR net6287 sky130_fd_sc_hd__buf_1
Xmax_length5553 net5548 VGND VGND VPWR VPWR net5553 sky130_fd_sc_hd__buf_1
XFILLER_0_182_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire800 net801 VGND VGND VPWR VPWR net800 sky130_fd_sc_hd__buf_1
X_14371_ _06581_ VGND VGND VPWR VPWR _00078_ sky130_fd_sc_hd__clkbuf_1
X_23569_ _03433_ _03436_ VGND VGND VPWR VPWR _03437_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_153_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire811 _12196_ VGND VGND VPWR VPWR net811 sky130_fd_sc_hd__buf_1
XFILLER_0_107_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire822 _09100_ VGND VGND VPWR VPWR net822 sky130_fd_sc_hd__buf_1
XFILLER_0_37_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire833 _06410_ VGND VGND VPWR VPWR net833 sky130_fd_sc_hd__dlymetal6s2s_1
X_16110_ _08094_ _08095_ _08096_ VGND VGND VPWR VPWR _08176_ sky130_fd_sc_hd__a21o_1
X_13322_ _05591_ _05594_ VGND VGND VPWR VPWR _05595_ sky130_fd_sc_hd__xnor2_1
X_25308_ clknet_leaf_72_clk _00191_ net8469 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.e\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire844 _05603_ VGND VGND VPWR VPWR net844 sky130_fd_sc_hd__buf_1
X_17090_ net1829 _09047_ net8050 VGND VGND VPWR VPWR _09048_ sky130_fd_sc_hd__o21ai_1
Xwire855 _03639_ VGND VGND VPWR VPWR net855 sky130_fd_sc_hd__buf_1
XFILLER_0_40_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire866 _12026_ VGND VGND VPWR VPWR net866 sky130_fd_sc_hd__buf_1
Xwire877 _09467_ VGND VGND VPWR VPWR net877 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16041_ _07841_ net1260 _08107_ VGND VGND VPWR VPWR _08108_ sky130_fd_sc_hd__o21a_1
XFILLER_0_150_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13253_ _05413_ _05414_ _05525_ VGND VGND VPWR VPWR _05526_ sky130_fd_sc_hd__o21a_1
Xwire888 _07669_ VGND VGND VPWR VPWR net888 sky130_fd_sc_hd__dlymetal6s2s_1
X_25239_ clknet_leaf_68_clk _00122_ net8454 VGND VGND VPWR VPWR matmul0.op\[0\] sky130_fd_sc_hd__dfrtp_1
Xwire899 _06572_ VGND VGND VPWR VPWR net899 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_150_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13184_ net7672 _05216_ VGND VGND VPWR VPWR _05457_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4140 net4141 VGND VGND VPWR VPWR net4140 sky130_fd_sc_hd__clkbuf_2
X_19800_ _11632_ _11633_ net6170 VGND VGND VPWR VPWR _11634_ sky130_fd_sc_hd__mux2_1
Xwire4151 net4152 VGND VGND VPWR VPWR net4151 sky130_fd_sc_hd__buf_1
Xwire4162 net4163 VGND VGND VPWR VPWR net4162 sky130_fd_sc_hd__buf_1
X_17992_ net6967 net7084 net7034 VGND VGND VPWR VPWR _09843_ sky130_fd_sc_hd__and3_2
Xwire4173 net4174 VGND VGND VPWR VPWR net4173 sky130_fd_sc_hd__buf_1
XFILLER_0_20_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3450 _07230_ VGND VGND VPWR VPWR net3450 sky130_fd_sc_hd__buf_1
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16943_ net1828 _08906_ VGND VGND VPWR VPWR _08907_ sky130_fd_sc_hd__nand2_1
X_19731_ net6030 _11508_ VGND VGND VPWR VPWR _11566_ sky130_fd_sc_hd__nand2_1
Xwire3461 net3462 VGND VGND VPWR VPWR net3461 sky130_fd_sc_hd__clkbuf_1
Xwire3472 net3473 VGND VGND VPWR VPWR net3472 sky130_fd_sc_hd__clkbuf_1
Xwire3483 _07150_ VGND VGND VPWR VPWR net3483 sky130_fd_sc_hd__buf_1
Xwire3494 _07118_ VGND VGND VPWR VPWR net3494 sky130_fd_sc_hd__buf_1
Xwire2760 _07190_ VGND VGND VPWR VPWR net2760 sky130_fd_sc_hd__buf_1
X_16874_ net1829 net1828 net8069 VGND VGND VPWR VPWR _08839_ sky130_fd_sc_hd__o21ai_1
X_19662_ _11492_ _11497_ _11493_ net3135 VGND VGND VPWR VPWR _11498_ sky130_fd_sc_hd__o22a_1
Xwire2771 _07153_ VGND VGND VPWR VPWR net2771 sky130_fd_sc_hd__clkbuf_1
Xwire2782 _07140_ VGND VGND VPWR VPWR net2782 sky130_fd_sc_hd__buf_1
XFILLER_0_189_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2793 _07134_ VGND VGND VPWR VPWR net2793 sky130_fd_sc_hd__clkbuf_1
X_15825_ net1529 net1850 VGND VGND VPWR VPWR _07895_ sky130_fd_sc_hd__nand2_1
X_18613_ net2134 _10459_ _10460_ net1203 net8966 VGND VGND VPWR VPWR _00442_ sky130_fd_sc_hd__a32o_1
XFILLER_0_95_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19593_ _11289_ net2106 VGND VGND VPWR VPWR _11430_ sky130_fd_sc_hd__or2_1
XFILLER_0_189_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15756_ _07824_ _07825_ _07823_ VGND VGND VPWR VPWR _07827_ sky130_fd_sc_hd__o21ai_1
X_18544_ _10386_ net1436 VGND VGND VPWR VPWR _10393_ sky130_fd_sc_hd__xnor2_1
X_12968_ net1140 net1004 VGND VGND VPWR VPWR _05241_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14707_ net7149 _06847_ VGND VGND VPWR VPWR _06850_ sky130_fd_sc_hd__or2_1
XFILLER_0_169_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18475_ net1774 _10323_ _10324_ VGND VGND VPWR VPWR _10325_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15687_ _07749_ _07757_ VGND VGND VPWR VPWR _07758_ sky130_fd_sc_hd__xnor2_1
X_12899_ net7715 net2978 net2335 VGND VGND VPWR VPWR _05172_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17426_ _09270_ _09325_ VGND VGND VPWR VPWR _09326_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14638_ net7437 matmul0.cos\[0\] net2878 VGND VGND VPWR VPWR _06803_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17357_ net3276 _09269_ VGND VGND VPWR VPWR _09270_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14569_ _06738_ _06744_ _06745_ VGND VGND VPWR VPWR _06746_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_56_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16308_ _08371_ VGND VGND VPWR VPWR _00225_ sky130_fd_sc_hd__clkbuf_1
X_17288_ _09195_ _09202_ VGND VGND VPWR VPWR _09203_ sky130_fd_sc_hd__nand2_1
X_19027_ net3214 net2528 _10832_ _10863_ net2530 VGND VGND VPWR VPWR _10864_ sky130_fd_sc_hd__a32o_1
X_16239_ _08302_ _08303_ VGND VGND VPWR VPWR _08304_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19929_ net6084 net3879 VGND VGND VPWR VPWR _11761_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22940_ net5327 pid_d.curr_int\[13\] _02813_ _02820_ VGND VGND VPWR VPWR _02829_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22871_ net8898 _02767_ VGND VGND VPWR VPWR _02768_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24610_ _04423_ _04463_ _04461_ VGND VGND VPWR VPWR _04465_ sky130_fd_sc_hd__a21oi_1
X_21822_ _01749_ _01751_ _01830_ VGND VGND VPWR VPWR _01831_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_183_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25590_ clknet_leaf_91_clk _00463_ net8425 VGND VGND VPWR VPWR cordic0.cos\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24541_ _04314_ _04372_ VGND VGND VPWR VPWR _04397_ sky130_fd_sc_hd__nor2_1
X_21753_ net5765 net5485 VGND VGND VPWR VPWR _01763_ sky130_fd_sc_hd__and2_1
XFILLER_0_148_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20704_ net6056 net1496 _12476_ VGND VGND VPWR VPWR _12478_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24472_ net2433 VGND VGND VPWR VPWR _04329_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21684_ _01689_ _01694_ VGND VGND VPWR VPWR _01695_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8428 net8426 VGND VGND VPWR VPWR net8428 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_50_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8439 net8440 VGND VGND VPWR VPWR net8439 sky130_fd_sc_hd__clkbuf_2
X_23423_ _03287_ _03292_ VGND VGND VPWR VPWR _03293_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7716 net7711 VGND VGND VPWR VPWR net7716 sky130_fd_sc_hd__buf_1
XFILLER_0_110_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20635_ net1495 _12413_ VGND VGND VPWR VPWR _12415_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7727 net7728 VGND VGND VPWR VPWR net7727 sky130_fd_sc_hd__buf_1
XFILLER_0_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7738 net7739 VGND VGND VPWR VPWR net7738 sky130_fd_sc_hd__buf_1
Xwire7749 net7753 VGND VGND VPWR VPWR net7749 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23354_ _02949_ _02951_ _02950_ VGND VGND VPWR VPWR _03224_ sky130_fd_sc_hd__o21a_1
X_20566_ net3848 _12275_ net2602 VGND VGND VPWR VPWR _12350_ sky130_fd_sc_hd__mux2_1
Xmax_length2713 net2714 VGND VGND VPWR VPWR net2713 sky130_fd_sc_hd__buf_1
XFILLER_0_116_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22305_ net944 _02308_ VGND VGND VPWR VPWR _02309_ sky130_fd_sc_hd__xor2_2
XFILLER_0_132_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23285_ _03152_ _03154_ VGND VGND VPWR VPWR _03155_ sky130_fd_sc_hd__xor2_1
XFILLER_0_131_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20497_ net6350 net1471 VGND VGND VPWR VPWR _12285_ sky130_fd_sc_hd__nand2_1
Xmax_length2779 _07142_ VGND VGND VPWR VPWR net2779 sky130_fd_sc_hd__buf_1
X_25024_ net7471 _04776_ _04777_ net7497 net462 VGND VGND VPWR VPWR _04778_ sky130_fd_sc_hd__a32o_1
X_22236_ _02237_ _02240_ VGND VGND VPWR VPWR _02241_ sky130_fd_sc_hd__xnor2_1
X_22167_ net339 VGND VGND VPWR VPWR _02173_ sky130_fd_sc_hd__inv_2
Xwire2001 _04643_ VGND VGND VPWR VPWR net2001 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2012 net2013 VGND VGND VPWR VPWR net2012 sky130_fd_sc_hd__clkbuf_1
X_21118_ net5564 net5949 net5929 net5911 VGND VGND VPWR VPWR _01134_ sky130_fd_sc_hd__a22o_1
Xwire2023 _04010_ VGND VGND VPWR VPWR net2023 sky130_fd_sc_hd__buf_1
X_22098_ _02102_ _02103_ VGND VGND VPWR VPWR _02105_ sky130_fd_sc_hd__or2_1
Xwire2034 _02715_ VGND VGND VPWR VPWR net2034 sky130_fd_sc_hd__buf_1
Xwire1311 net1312 VGND VGND VPWR VPWR net1311 sky130_fd_sc_hd__buf_1
Xwire2056 net2057 VGND VGND VPWR VPWR net2056 sky130_fd_sc_hd__buf_1
X_13940_ net837 net907 VGND VGND VPWR VPWR _06206_ sky130_fd_sc_hd__nor2_1
Xwire1322 net1323 VGND VGND VPWR VPWR net1322 sky130_fd_sc_hd__buf_1
Xwire2067 _01779_ VGND VGND VPWR VPWR net2067 sky130_fd_sc_hd__buf_2
X_25926_ clknet_leaf_1_clk net9197 net8413 VGND VGND VPWR VPWR pid_d.prev_int\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_21049_ _01031_ _01059_ _01064_ VGND VGND VPWR VPWR _01065_ sky130_fd_sc_hd__a21o_1
Xwire1333 net1334 VGND VGND VPWR VPWR net1333 sky130_fd_sc_hd__buf_1
Xwire2078 _12503_ VGND VGND VPWR VPWR net2078 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1344 net1345 VGND VGND VPWR VPWR net1344 sky130_fd_sc_hd__clkbuf_1
Xwire2089 net2090 VGND VGND VPWR VPWR net2089 sky130_fd_sc_hd__buf_1
Xwire1366 _04543_ VGND VGND VPWR VPWR net1366 sky130_fd_sc_hd__buf_1
X_25857_ clknet_leaf_19_clk _00730_ net8624 VGND VGND VPWR VPWR pid_q.mult0.a\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13871_ net996 _06071_ VGND VGND VPWR VPWR _06138_ sky130_fd_sc_hd__and2b_1
Xwire1388 _02571_ VGND VGND VPWR VPWR net1388 sky130_fd_sc_hd__buf_1
XFILLER_0_97_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1399 net1400 VGND VGND VPWR VPWR net1399 sky130_fd_sc_hd__buf_1
X_15610_ net6542 matmul0.matmul_stage_inst.c\[14\] matmul0.matmul_stage_inst.b\[14\]
+ net6614 VGND VGND VPWR VPWR _07682_ sky130_fd_sc_hd__a22oi_1
X_24808_ _04631_ VGND VGND VPWR VPWR _04632_ sky130_fd_sc_hd__inv_2
X_12822_ net7737 net2345 net2342 VGND VGND VPWR VPWR _05095_ sky130_fd_sc_hd__and3_1
X_16590_ _08642_ VGND VGND VPWR VPWR _00236_ sky130_fd_sc_hd__clkbuf_1
X_25788_ clknet_leaf_63_clk _00661_ net8672 VGND VGND VPWR VPWR matmul0.beta_pass\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15541_ net3532 net3552 VGND VGND VPWR VPWR _07614_ sky130_fd_sc_hd__nor2_1
X_24739_ net8007 _04565_ _04566_ VGND VGND VPWR VPWR _04571_ sky130_fd_sc_hd__and3_1
X_12753_ net1354 VGND VGND VPWR VPWR _05026_ sky130_fd_sc_hd__buf_1
Xmax_length6040 net6035 VGND VGND VPWR VPWR net6040 sky130_fd_sc_hd__clkbuf_1
X_18260_ _10108_ _10110_ VGND VGND VPWR VPWR _10111_ sky130_fd_sc_hd__xnor2_1
X_15472_ _07343_ _07344_ net1542 VGND VGND VPWR VPWR _07546_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12684_ net2976 VGND VGND VPWR VPWR _04957_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length5350 pid_d.out\[10\] VGND VGND VPWR VPWR net5350 sky130_fd_sc_hd__clkbuf_1
X_17211_ _09146_ _09148_ _09151_ net6819 VGND VGND VPWR VPWR _09160_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_7_Left_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14423_ _06621_ VGND VGND VPWR VPWR _00090_ sky130_fd_sc_hd__clkbuf_1
Xwire8940 net8941 VGND VGND VPWR VPWR net8940 sky130_fd_sc_hd__clkbuf_1
X_18191_ _10039_ _10041_ VGND VGND VPWR VPWR _10042_ sky130_fd_sc_hd__xnor2_1
Xwire8951 net8952 VGND VGND VPWR VPWR net8951 sky130_fd_sc_hd__clkbuf_1
Xmax_length5394 net5395 VGND VGND VPWR VPWR net5394 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_112_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17142_ _09095_ VGND VGND VPWR VPWR _09096_ sky130_fd_sc_hd__buf_2
Xwire630 _04595_ VGND VGND VPWR VPWR net630 sky130_fd_sc_hd__clkbuf_1
X_14354_ _06567_ matmul0.a_in\[8\] net905 VGND VGND VPWR VPWR _06568_ sky130_fd_sc_hd__mux2_1
Xwire641 net642 VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__clkbuf_1
Xwire652 _01549_ VGND VGND VPWR VPWR net652 sky130_fd_sc_hd__clkbuf_1
X_13305_ net7619 net2339 net1967 VGND VGND VPWR VPWR _05578_ sky130_fd_sc_hd__and3_1
Xwire663 net664 VGND VGND VPWR VPWR net663 sky130_fd_sc_hd__buf_1
XFILLER_0_24_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire674 _07562_ VGND VGND VPWR VPWR net674 sky130_fd_sc_hd__buf_1
X_17073_ net4062 VGND VGND VPWR VPWR _09031_ sky130_fd_sc_hd__buf_1
X_14285_ net2915 VGND VGND VPWR VPWR _06519_ sky130_fd_sc_hd__clkbuf_2
Xwire685 _04801_ VGND VGND VPWR VPWR net685 sky130_fd_sc_hd__buf_1
Xwire696 _03468_ VGND VGND VPWR VPWR net696 sky130_fd_sc_hd__buf_1
XFILLER_0_122_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16024_ _08016_ net673 VGND VGND VPWR VPWR _08091_ sky130_fd_sc_hd__or2_1
X_13236_ _05505_ _05508_ VGND VGND VPWR VPWR _05509_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_126_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13167_ net7756 net2324 net2320 VGND VGND VPWR VPWR _05440_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13098_ net7728 net1616 _05257_ _05258_ VGND VGND VPWR VPWR _05371_ sky130_fd_sc_hd__a22o_1
X_17975_ net3245 _09825_ net1779 VGND VGND VPWR VPWR _09826_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3280 net3281 VGND VGND VPWR VPWR net3280 sky130_fd_sc_hd__buf_1
Xwire3291 net3292 VGND VGND VPWR VPWR net3291 sky130_fd_sc_hd__buf_1
X_19714_ net570 net3857 VGND VGND VPWR VPWR _11550_ sky130_fd_sc_hd__or2_1
X_16926_ cordic0.slte0.opA\[5\] VGND VGND VPWR VPWR _08890_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2590 _09069_ VGND VGND VPWR VPWR net2590 sky130_fd_sc_hd__clkbuf_1
X_19645_ _11429_ _11480_ VGND VGND VPWR VPWR _11482_ sky130_fd_sc_hd__nor2_1
X_16857_ net6254 net6195 net6498 VGND VGND VPWR VPWR _08822_ sky130_fd_sc_hd__mux2_1
X_15808_ _07869_ _07877_ VGND VGND VPWR VPWR _07878_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19576_ net1416 _11412_ VGND VGND VPWR VPWR _11413_ sky130_fd_sc_hd__xnor2_2
X_16788_ net7585 matmul0.a\[13\] net3372 VGND VGND VPWR VPWR _08784_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15739_ net2672 VGND VGND VPWR VPWR _07810_ sky130_fd_sc_hd__clkbuf_1
X_18527_ net2129 _10375_ VGND VGND VPWR VPWR _10376_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18458_ net1207 _10307_ VGND VGND VPWR VPWR _10308_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17409_ net2575 _09312_ VGND VGND VPWR VPWR _09313_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18389_ net3253 net3267 _10239_ VGND VGND VPWR VPWR _10240_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_117_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20420_ net6467 _12118_ _12175_ VGND VGND VPWR VPWR _12216_ sky130_fd_sc_hd__or3_1
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20351_ net1490 _12152_ net3316 VGND VGND VPWR VPWR _12153_ sky130_fd_sc_hd__a21o_1
X_23070_ net5017 net4655 VGND VGND VPWR VPWR _02940_ sky130_fd_sc_hd__nand2_2
Xwire4909 net4910 VGND VGND VPWR VPWR net4909 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20282_ net9208 _12087_ _12088_ net2091 VGND VGND VPWR VPWR _00483_ sky130_fd_sc_hd__a22o_1
XFILLER_0_178_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22021_ _02026_ _02027_ VGND VGND VPWR VPWR _02028_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold15 cordic0.cos\[3\] VGND VGND VPWR VPWR net8968 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 matmul0.matmul_stage_inst.a\[1\] VGND VGND VPWR VPWR net8979 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 pid_q.target\[14\] VGND VGND VPWR VPWR net8990 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 _00407_ VGND VGND VPWR VPWR net9001 sky130_fd_sc_hd__dlygate4sd3_1
X_23972_ net932 _03835_ VGND VGND VPWR VPWR _03836_ sky130_fd_sc_hd__xnor2_1
Xhold59 pid_d.prev_error\[12\] VGND VGND VPWR VPWR net9012 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length8915 net8916 VGND VGND VPWR VPWR net8915 sky130_fd_sc_hd__clkbuf_1
X_25711_ clknet_leaf_9_clk _00584_ net8552 VGND VGND VPWR VPWR pid_d.mult0.a\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_22923_ net5975 _02812_ VGND VGND VPWR VPWR _02814_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25642_ clknet_leaf_102_clk _00515_ net8366 VGND VGND VPWR VPWR cordic0.vec\[0\]\[14\]
+ sky130_fd_sc_hd__dfstp_1
X_22854_ net5981 _02747_ _02751_ VGND VGND VPWR VPWR _02752_ sky130_fd_sc_hd__o21a_1
XFILLER_0_168_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21805_ _01812_ _01813_ VGND VGND VPWR VPWR _01815_ sky130_fd_sc_hd__or2_1
X_25573_ clknet_leaf_97_clk _00446_ net8398 VGND VGND VPWR VPWR cordic0.sin\[7\] sky130_fd_sc_hd__dfrtp_1
X_22785_ _02700_ VGND VGND VPWR VPWR _00619_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24524_ _04315_ _04374_ _04375_ _04314_ _04380_ VGND VGND VPWR VPWR _04381_ sky130_fd_sc_hd__o221a_1
X_21736_ _01658_ _01685_ _01745_ VGND VGND VPWR VPWR _01746_ sky130_fd_sc_hd__a21o_1
Xwire8203 net33 VGND VGND VPWR VPWR net8203 sky130_fd_sc_hd__clkbuf_1
Xwire8214 net8215 VGND VGND VPWR VPWR net8214 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8225 net8226 VGND VGND VPWR VPWR net8225 sky130_fd_sc_hd__clkbuf_1
Xwire8236 net8237 VGND VGND VPWR VPWR net8236 sky130_fd_sc_hd__clkbuf_1
Xwire7502 net7501 VGND VGND VPWR VPWR net7502 sky130_fd_sc_hd__clkbuf_1
X_24455_ _04227_ net1012 _04312_ VGND VGND VPWR VPWR _04313_ sky130_fd_sc_hd__a21o_1
XFILLER_0_188_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21667_ _01562_ _01564_ VGND VGND VPWR VPWR _01678_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8247 net8248 VGND VGND VPWR VPWR net8247 sky130_fd_sc_hd__clkbuf_1
Xwire7513 net7514 VGND VGND VPWR VPWR net7513 sky130_fd_sc_hd__clkbuf_1
Xwire8258 net8259 VGND VGND VPWR VPWR net8258 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7524 net7521 VGND VGND VPWR VPWR net7524 sky130_fd_sc_hd__clkbuf_2
Xwire8269 net8270 VGND VGND VPWR VPWR net8269 sky130_fd_sc_hd__clkbuf_1
X_23406_ _03272_ _03275_ VGND VGND VPWR VPWR _03276_ sky130_fd_sc_hd__xnor2_1
Xwire7535 net7536 VGND VGND VPWR VPWR net7535 sky130_fd_sc_hd__clkbuf_1
Xwire7546 net7547 VGND VGND VPWR VPWR net7546 sky130_fd_sc_hd__clkbuf_1
X_20618_ net1395 _12398_ VGND VGND VPWR VPWR _12399_ sky130_fd_sc_hd__xor2_1
Xwire6801 net6797 VGND VGND VPWR VPWR net6801 sky130_fd_sc_hd__buf_1
X_24386_ _04243_ _04244_ VGND VGND VPWR VPWR _04245_ sky130_fd_sc_hd__or2b_1
Xwire7557 net7558 VGND VGND VPWR VPWR net7557 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21598_ net5383 net3106 VGND VGND VPWR VPWR _01610_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7568 net7569 VGND VGND VPWR VPWR net7568 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7579 net7580 VGND VGND VPWR VPWR net7579 sky130_fd_sc_hd__clkbuf_1
Xmax_length3266 _09615_ VGND VGND VPWR VPWR net3266 sky130_fd_sc_hd__buf_1
X_23337_ _02933_ _02935_ _03206_ VGND VGND VPWR VPWR _03207_ sky130_fd_sc_hd__a21bo_1
Xmax_length3277 _09268_ VGND VGND VPWR VPWR net3277 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire6845 net6846 VGND VGND VPWR VPWR net6845 sky130_fd_sc_hd__buf_1
XFILLER_0_61_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20549_ _12301_ _12302_ net6326 VGND VGND VPWR VPWR _12334_ sky130_fd_sc_hd__a21oi_1
Xwire6856 net6854 VGND VGND VPWR VPWR net6856 sky130_fd_sc_hd__buf_1
Xmax_length2554 _09720_ VGND VGND VPWR VPWR net2554 sky130_fd_sc_hd__clkbuf_2
X_14070_ _06221_ net1125 VGND VGND VPWR VPWR _06333_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23268_ _03134_ _03137_ _03135_ VGND VGND VPWR VPWR _03138_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_89_Left_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13021_ _05187_ VGND VGND VPWR VPWR _05294_ sky130_fd_sc_hd__buf_1
X_25007_ net4466 net5179 VGND VGND VPWR VPWR _04763_ sky130_fd_sc_hd__xor2_1
X_22219_ _02130_ _02131_ _02129_ VGND VGND VPWR VPWR _02224_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23199_ _03062_ _03067_ _03068_ VGND VGND VPWR VPWR _03069_ sky130_fd_sc_hd__o21a_1
XFILLER_0_195_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14972_ net2839 _07045_ VGND VGND VPWR VPWR _07046_ sky130_fd_sc_hd__nor2_1
X_17760_ _09605_ _09610_ VGND VGND VPWR VPWR _09611_ sky130_fd_sc_hd__xor2_1
Xwire1130 _05640_ VGND VGND VPWR VPWR net1130 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1141 net1142 VGND VGND VPWR VPWR net1141 sky130_fd_sc_hd__clkbuf_1
X_13923_ _06185_ _06188_ VGND VGND VPWR VPWR _06189_ sky130_fd_sc_hd__xnor2_2
Xwire1152 net1153 VGND VGND VPWR VPWR net1152 sky130_fd_sc_hd__clkbuf_1
X_16711_ net7224 _08738_ net6548 VGND VGND VPWR VPWR _08739_ sky130_fd_sc_hd__mux2_1
X_17691_ _09561_ net2565 net964 VGND VGND VPWR VPWR _09571_ sky130_fd_sc_hd__and3_1
Xwire1163 _03643_ VGND VGND VPWR VPWR net1163 sky130_fd_sc_hd__dlymetal6s2s_1
X_25909_ clknet_leaf_29_clk _00782_ net8656 VGND VGND VPWR VPWR pid_q.out\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1174 _01656_ VGND VGND VPWR VPWR net1174 sky130_fd_sc_hd__buf_1
Xwire1185 _01018_ VGND VGND VPWR VPWR net1185 sky130_fd_sc_hd__buf_1
X_19430_ net6070 net6105 VGND VGND VPWR VPWR _11267_ sky130_fd_sc_hd__xor2_2
Xwire1196 _10419_ VGND VGND VPWR VPWR net1196 sky130_fd_sc_hd__buf_1
X_16642_ matmul0.matmul_stage_inst.mult1\[3\] VGND VGND VPWR VPWR _08679_ sky130_fd_sc_hd__inv_2
X_13854_ _06053_ _06054_ net7669 net1312 VGND VGND VPWR VPWR _06121_ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_98_Left_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12805_ _04955_ _05074_ _05076_ _04941_ _05077_ VGND VGND VPWR VPWR _05078_ sky130_fd_sc_hd__a221o_1
X_19361_ _11166_ _11197_ VGND VGND VPWR VPWR _11198_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16573_ _08622_ _08631_ VGND VGND VPWR VPWR _08632_ sky130_fd_sc_hd__xnor2_1
X_13785_ net7636 net2322 net2318 VGND VGND VPWR VPWR _06053_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18312_ net7040 _10161_ _10108_ _10162_ VGND VGND VPWR VPWR _10163_ sky130_fd_sc_hd__a31o_1
X_15524_ _07593_ _07596_ VGND VGND VPWR VPWR _07597_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout8620 net8644 VGND VGND VPWR VPWR net8620 sky130_fd_sc_hd__clkbuf_2
X_12736_ _04980_ _04981_ VGND VGND VPWR VPWR _05009_ sky130_fd_sc_hd__xnor2_1
X_19292_ _11126_ _11128_ net6243 VGND VGND VPWR VPWR _11129_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8653 net8658 VGND VGND VPWR VPWR net8653 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18243_ net6894 net6922 VGND VGND VPWR VPWR _10094_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout8664 net8670 VGND VGND VPWR VPWR net8664 sky130_fd_sc_hd__buf_1
X_15455_ net3412 _07016_ VGND VGND VPWR VPWR _07529_ sky130_fd_sc_hd__nand2_1
Xfanout7930 net7936 VGND VGND VPWR VPWR net7930 sky130_fd_sc_hd__clkbuf_1
X_12667_ _04935_ _04939_ VGND VGND VPWR VPWR _04940_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length5180 pid_q.curr_int\[2\] VGND VGND VPWR VPWR net5180 sky130_fd_sc_hd__dlymetal6s2s_1
X_14406_ net1548 VGND VGND VPWR VPWR _06608_ sky130_fd_sc_hd__buf_1
XFILLER_0_5_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8770 net8771 VGND VGND VPWR VPWR net8770 sky130_fd_sc_hd__buf_1
X_18174_ _09686_ _09787_ _09784_ VGND VGND VPWR VPWR _10025_ sky130_fd_sc_hd__o21a_1
X_15386_ _07459_ net1116 _07430_ VGND VGND VPWR VPWR _07460_ sky130_fd_sc_hd__a21o_1
X_12598_ net7531 net8904 net4389 VGND VGND VPWR VPWR _04878_ sky130_fd_sc_hd__and3_1
X_17125_ net6932 _09079_ _09080_ VGND VGND VPWR VPWR _00333_ sky130_fd_sc_hd__a21bo_1
Xwire460 net461 VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__clkbuf_1
X_14337_ net7320 net1299 net2896 pid_d.out\[4\] _06554_ VGND VGND VPWR VPWR _06555_
+ sky130_fd_sc_hd__a221o_1
Xwire471 _01925_ VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__buf_1
XFILLER_0_40_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire482 net483 VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__clkbuf_1
Xwire493 _08160_ VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__buf_1
X_17056_ net7057 _08977_ VGND VGND VPWR VPWR _09015_ sky130_fd_sc_hd__xnor2_1
X_14268_ net61 net2931 net2278 net9053 VGND VGND VPWR VPWR _00041_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16007_ _08064_ _08074_ VGND VGND VPWR VPWR _08075_ sky130_fd_sc_hd__xnor2_1
X_13219_ net7672 _05216_ _05458_ VGND VGND VPWR VPWR _05492_ sky130_fd_sc_hd__a21o_1
X_14199_ _06456_ _06458_ VGND VGND VPWR VPWR _06459_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17958_ net3952 _09630_ VGND VGND VPWR VPWR _09809_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_164_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16909_ net6373 _08871_ VGND VGND VPWR VPWR _08873_ sky130_fd_sc_hd__nand2_1
X_17889_ net6966 net7005 VGND VGND VPWR VPWR _09740_ sky130_fd_sc_hd__xnor2_1
X_19628_ _11190_ _11191_ net6222 VGND VGND VPWR VPWR _11465_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19559_ net2513 _10938_ VGND VGND VPWR VPWR _11396_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22570_ net3769 _02550_ _02551_ VGND VGND VPWR VPWR _02552_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21521_ net5971 _01428_ _01429_ pid_d.prev_error\[2\] VGND VGND VPWR VPWR _01534_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_173_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24240_ _04097_ net852 VGND VGND VPWR VPWR _04101_ sky130_fd_sc_hd__and2_1
X_21452_ net5616 _00851_ _01349_ _01464_ _01347_ VGND VGND VPWR VPWR _01465_ sky130_fd_sc_hd__o32a_1
Xwire6108 net6104 VGND VGND VPWR VPWR net6108 sky130_fd_sc_hd__buf_1
XFILLER_0_160_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6119 net6121 VGND VGND VPWR VPWR net6119 sky130_fd_sc_hd__clkbuf_2
X_20403_ net1466 _12200_ net3355 VGND VGND VPWR VPWR _12201_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24171_ _04031_ _04032_ VGND VGND VPWR VPWR _04033_ sky130_fd_sc_hd__nand2_1
Xwire5407 net5408 VGND VGND VPWR VPWR net5407 sky130_fd_sc_hd__buf_1
X_21383_ _01276_ net1390 net1391 VGND VGND VPWR VPWR _01397_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_31_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5418 net5413 VGND VGND VPWR VPWR net5418 sky130_fd_sc_hd__buf_1
X_23122_ _02969_ _02970_ VGND VGND VPWR VPWR _02992_ sky130_fd_sc_hd__xnor2_1
X_20334_ _12132_ _12136_ VGND VGND VPWR VPWR _12137_ sky130_fd_sc_hd__xnor2_1
Xwire4717 net4718 VGND VGND VPWR VPWR net4717 sky130_fd_sc_hd__buf_1
XFILLER_0_101_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4739 net4740 VGND VGND VPWR VPWR net4739 sky130_fd_sc_hd__buf_1
X_23053_ net4865 net4772 net4913 VGND VGND VPWR VPWR _02923_ sky130_fd_sc_hd__a21o_1
X_20265_ net3 _12072_ net8121 VGND VGND VPWR VPWR _12076_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22004_ _02010_ _02011_ VGND VGND VPWR VPWR _02012_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20196_ net3145 _11996_ net2580 VGND VGND VPWR VPWR _12021_ sky130_fd_sc_hd__a21oi_1
Xinput105 pid_d_data[2] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_1
Xinput116 pid_q_addr[11] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_1
Xinput127 pid_q_addr[7] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_1
Xinput138 pid_q_data[2] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_1
Xmax_length8701 net8696 VGND VGND VPWR VPWR net8701 sky130_fd_sc_hd__buf_1
X_23955_ net5071 net5036 VGND VGND VPWR VPWR _03819_ sky130_fd_sc_hd__xor2_1
X_22906_ pid_d.out\[10\] _02795_ _02798_ VGND VGND VPWR VPWR _02799_ sky130_fd_sc_hd__mux2_1
X_23886_ net1163 _03647_ _03648_ VGND VGND VPWR VPWR _03751_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_195_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25625_ clknet_leaf_117_clk _00498_ net8332 VGND VGND VPWR VPWR cordic0.slte0.opA\[15\]
+ sky130_fd_sc_hd__dfrtp_2
X_22837_ _02734_ _02736_ VGND VGND VPWR VPWR _02737_ sky130_fd_sc_hd__and2_1
XFILLER_0_183_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13570_ net7895 net1928 _05839_ VGND VGND VPWR VPWR _05841_ sky130_fd_sc_hd__a21o_1
X_25556_ clknet_leaf_77_clk net6619 net8439 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22768_ net4302 net8936 VGND VGND VPWR VPWR _02690_ sky130_fd_sc_hd__and2_1
Xwire8000 net8001 VGND VGND VPWR VPWR net8000 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24507_ _04357_ _04363_ VGND VGND VPWR VPWR _04364_ sky130_fd_sc_hd__xnor2_2
Xwire8022 net8023 VGND VGND VPWR VPWR net8022 sky130_fd_sc_hd__buf_1
X_21719_ _01728_ _01638_ _01729_ VGND VGND VPWR VPWR _01730_ sky130_fd_sc_hd__a21o_1
Xwire8033 pid_q.target\[1\] VGND VGND VPWR VPWR net8033 sky130_fd_sc_hd__clkbuf_1
X_25487_ clknet_leaf_46_clk _00367_ net8780 VGND VGND VPWR VPWR svm0.tA\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22699_ pid_d.ki\[10\] net2446 net3696 pid_d.kp\[10\] VGND VGND VPWR VPWR _02641_
+ sky130_fd_sc_hd__a22o_1
Xwire8044 net8045 VGND VGND VPWR VPWR net8044 sky130_fd_sc_hd__clkbuf_2
Xfanout6503 cordic0.gm0.iter\[1\] VGND VGND VPWR VPWR net6503 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8055 net8056 VGND VGND VPWR VPWR net8055 sky130_fd_sc_hd__buf_1
Xwire7310 net7311 VGND VGND VPWR VPWR net7310 sky130_fd_sc_hd__clkbuf_1
X_15240_ _07306_ net3443 VGND VGND VPWR VPWR _07314_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7321 net7322 VGND VGND VPWR VPWR net7321 sky130_fd_sc_hd__clkbuf_1
X_24438_ net4515 VGND VGND VPWR VPWR _04296_ sky130_fd_sc_hd__inv_2
Xwire8066 net8067 VGND VGND VPWR VPWR net8066 sky130_fd_sc_hd__clkbuf_1
Xwire8077 net8078 VGND VGND VPWR VPWR net8077 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7332 net7333 VGND VGND VPWR VPWR net7332 sky130_fd_sc_hd__buf_1
Xwire8088 net8089 VGND VGND VPWR VPWR net8088 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout6547 net6562 VGND VGND VPWR VPWR net6547 sky130_fd_sc_hd__buf_1
Xwire7343 net7344 VGND VGND VPWR VPWR net7343 sky130_fd_sc_hd__buf_1
Xfanout5802 pid_d.mult0.b\[7\] VGND VGND VPWR VPWR net5802 sky130_fd_sc_hd__buf_1
Xwire8099 net91 VGND VGND VPWR VPWR net8099 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7354 net7355 VGND VGND VPWR VPWR net7354 sky130_fd_sc_hd__clkbuf_1
Xwire7365 net7366 VGND VGND VPWR VPWR net7365 sky130_fd_sc_hd__buf_1
XFILLER_0_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6620 net6621 VGND VGND VPWR VPWR net6620 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire7376 net7377 VGND VGND VPWR VPWR net7376 sky130_fd_sc_hd__buf_1
X_15171_ net4222 net4220 net4206 net4202 VGND VGND VPWR VPWR _07245_ sky130_fd_sc_hd__o22a_1
Xwire6631 net6626 VGND VGND VPWR VPWR net6631 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_151_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24369_ net1655 net1654 _04137_ VGND VGND VPWR VPWR _04228_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6642 net6643 VGND VGND VPWR VPWR net6642 sky130_fd_sc_hd__clkbuf_1
Xwire7387 net7388 VGND VGND VPWR VPWR net7387 sky130_fd_sc_hd__clkbuf_1
Xwire6653 net6654 VGND VGND VPWR VPWR net6653 sky130_fd_sc_hd__clkbuf_1
Xwire7398 net7399 VGND VGND VPWR VPWR net7398 sky130_fd_sc_hd__clkbuf_1
X_14122_ _06382_ _06383_ VGND VGND VPWR VPWR _06384_ sky130_fd_sc_hd__xnor2_1
Xwire6664 net6665 VGND VGND VPWR VPWR net6664 sky130_fd_sc_hd__buf_1
Xwire6675 net6676 VGND VGND VPWR VPWR net6675 sky130_fd_sc_hd__clkbuf_1
Xwire5930 net5928 VGND VGND VPWR VPWR net5930 sky130_fd_sc_hd__buf_1
XFILLER_0_162_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5963 net5958 VGND VGND VPWR VPWR net5963 sky130_fd_sc_hd__buf_1
X_14053_ _06311_ _06314_ VGND VGND VPWR VPWR _06317_ sky130_fd_sc_hd__nor2_1
Xwire5974 pid_d.curr_int\[15\] VGND VGND VPWR VPWR net5974 sky130_fd_sc_hd__buf_1
X_18930_ net9074 net2287 net1450 _10769_ VGND VGND VPWR VPWR _00450_ sky130_fd_sc_hd__a31o_1
Xwire5996 net5997 VGND VGND VPWR VPWR net5996 sky130_fd_sc_hd__buf_1
XFILLER_0_30_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13004_ _05269_ _05276_ VGND VGND VPWR VPWR _05277_ sky130_fd_sc_hd__xnor2_2
X_18861_ _10679_ VGND VGND VPWR VPWR _10703_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17812_ net6856 VGND VGND VPWR VPWR _09663_ sky130_fd_sc_hd__inv_2
X_18792_ net3957 _10632_ _10635_ VGND VGND VPWR VPWR _10636_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_27_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17743_ net6453 net6649 net6449 VGND VGND VPWR VPWR _09596_ sky130_fd_sc_hd__o21ai_1
X_14955_ net6620 net6640 matmul0.matmul_stage_inst.f\[7\] VGND VGND VPWR VPWR _07029_
+ sky130_fd_sc_hd__o21a_1
X_13906_ _06167_ _06171_ VGND VGND VPWR VPWR _06172_ sky130_fd_sc_hd__xnor2_2
X_17674_ net4002 svm0.tA\[2\] _09553_ VGND VGND VPWR VPWR _09554_ sky130_fd_sc_hd__a21o_1
X_14886_ matmul0.b\[15\] matmul0.matmul_stage_inst.f\[15\] net3623 VGND VGND VPWR
+ VPWR _06961_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19413_ _11245_ _11246_ VGND VGND VPWR VPWR _11250_ sky130_fd_sc_hd__nand2_1
X_13837_ _06098_ _06103_ VGND VGND VPWR VPWR _06104_ sky130_fd_sc_hd__xnor2_1
X_16625_ _08664_ VGND VGND VPWR VPWR _00249_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19344_ net6179 net6289 net3890 VGND VGND VPWR VPWR _11181_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16556_ _08258_ _08613_ _08614_ VGND VGND VPWR VPWR _08615_ sky130_fd_sc_hd__and3_1
X_13768_ net7696 net2308 net1953 VGND VGND VPWR VPWR _06036_ sky130_fd_sc_hd__and3_1
XFILLER_0_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12719_ _04990_ _04991_ VGND VGND VPWR VPWR _04992_ sky130_fd_sc_hd__xnor2_1
X_15507_ net4160 net4156 net4105 net4101 VGND VGND VPWR VPWR _07580_ sky130_fd_sc_hd__o22a_1
XFILLER_0_72_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout8450 net8456 VGND VGND VPWR VPWR net8450 sky130_fd_sc_hd__clkbuf_2
X_19275_ _10907_ _10908_ _10862_ VGND VGND VPWR VPWR _11112_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16487_ net208 _08542_ _08543_ VGND VGND VPWR VPWR _08547_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_13699_ net7615 net1338 net1563 net1148 net7654 VGND VGND VPWR VPWR _05968_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_57_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18226_ _10038_ VGND VGND VPWR VPWR _10077_ sky130_fd_sc_hd__inv_2
X_15438_ _07377_ _07511_ _07373_ _07374_ VGND VGND VPWR VPWR _07512_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout7771 svm0.periodTop\[7\] VGND VGND VPWR VPWR net7771 sky130_fd_sc_hd__buf_1
XFILLER_0_142_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18157_ _10003_ _10005_ net1212 VGND VGND VPWR VPWR _10008_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15369_ _07419_ _07442_ VGND VGND VPWR VPWR _07443_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire290 _04327_ VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__clkbuf_1
X_17108_ _09063_ _09064_ VGND VGND VPWR VPWR _09065_ sky130_fd_sc_hd__nor2_1
X_18088_ _09932_ _09938_ VGND VGND VPWR VPWR _09939_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_29_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17039_ net1483 _08980_ _08998_ VGND VGND VPWR VPWR _08999_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20050_ net6058 _11490_ VGND VGND VPWR VPWR _11879_ sky130_fd_sc_hd__nor2_1
XFILLER_0_175_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23740_ net5120 net3744 net5155 VGND VGND VPWR VPWR _03606_ sky130_fd_sc_hd__o21a_1
X_20952_ _00944_ _00963_ _00967_ VGND VGND VPWR VPWR _00968_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_36_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23671_ _03525_ _03536_ VGND VGND VPWR VPWR _03538_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20883_ _00897_ _00898_ VGND VGND VPWR VPWR _00899_ sky130_fd_sc_hd__xnor2_1
X_25410_ clknet_leaf_75_clk _00293_ net8511 VGND VGND VPWR VPWR matmul0.a\[13\] sky130_fd_sc_hd__dfrtp_1
X_22622_ net8993 _02544_ _02546_ net858 VGND VGND VPWR VPWR _00564_ sky130_fd_sc_hd__a22o_1
XFILLER_0_191_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length5938 net5940 VGND VGND VPWR VPWR net5938 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25341_ clknet_leaf_56_clk _00224_ net8723 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_22553_ pid_d.curr_error\[14\] net3018 net2460 VGND VGND VPWR VPWR _02539_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21504_ net1182 net1181 _01516_ VGND VGND VPWR VPWR _01517_ sky130_fd_sc_hd__a21oi_1
X_25272_ clknet_leaf_93_clk _00155_ net8446 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.c\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22484_ net5671 _02484_ net5407 VGND VGND VPWR VPWR _02485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length805 _01816_ VGND VGND VPWR VPWR net805 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24223_ net3040 _04083_ VGND VGND VPWR VPWR _04084_ sky130_fd_sc_hd__xnor2_1
X_21435_ net3807 net5654 VGND VGND VPWR VPWR _01448_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5204 net5205 VGND VGND VPWR VPWR net5204 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5215 net5216 VGND VGND VPWR VPWR net5215 sky130_fd_sc_hd__clkbuf_2
Xwire5226 net5227 VGND VGND VPWR VPWR net5226 sky130_fd_sc_hd__clkbuf_1
X_24154_ _04003_ _04015_ VGND VGND VPWR VPWR _04016_ sky130_fd_sc_hd__xnor2_1
Xwire5237 net5238 VGND VGND VPWR VPWR net5237 sky130_fd_sc_hd__buf_1
X_21366_ net5963 net5382 VGND VGND VPWR VPWR _01380_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_169_Right_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5248 net5249 VGND VGND VPWR VPWR net5248 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5259 net5260 VGND VGND VPWR VPWR net5259 sky130_fd_sc_hd__buf_1
XFILLER_0_114_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23105_ net4948 net4774 VGND VGND VPWR VPWR _02975_ sky130_fd_sc_hd__nand2_1
Xwire4536 net4537 VGND VGND VPWR VPWR net4536 sky130_fd_sc_hd__buf_1
X_20317_ net6515 net1482 _08943_ VGND VGND VPWR VPWR _12121_ sky130_fd_sc_hd__or3_1
Xwire4547 net4549 VGND VGND VPWR VPWR net4547 sky130_fd_sc_hd__clkbuf_1
X_24085_ _03946_ _03854_ _03947_ VGND VGND VPWR VPWR _03948_ sky130_fd_sc_hd__a21o_1
Xwire3802 _01317_ VGND VGND VPWR VPWR net3802 sky130_fd_sc_hd__clkbuf_1
X_21297_ _01306_ _01311_ VGND VGND VPWR VPWR _01312_ sky130_fd_sc_hd__xor2_1
Xwire3813 net3814 VGND VGND VPWR VPWR net3813 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3824 _00977_ VGND VGND VPWR VPWR net3824 sky130_fd_sc_hd__clkbuf_1
X_23036_ _02899_ _02904_ VGND VGND VPWR VPWR _02906_ sky130_fd_sc_hd__or2_1
Xwire3835 _00917_ VGND VGND VPWR VPWR net3835 sky130_fd_sc_hd__clkbuf_1
X_20248_ net15 _12062_ VGND VGND VPWR VPWR _12063_ sky130_fd_sc_hd__xnor2_1
Xwire3846 _12296_ VGND VGND VPWR VPWR net3846 sky130_fd_sc_hd__buf_1
Xwire3857 net3858 VGND VGND VPWR VPWR net3857 sky130_fd_sc_hd__buf_1
X_20179_ _11998_ _11999_ _12002_ _12004_ VGND VGND VPWR VPWR _12005_ sky130_fd_sc_hd__o22a_1
XFILLER_0_157_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24987_ _04748_ VGND VGND VPWR VPWR _00773_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14740_ net7161 net7164 net7158 net7156 net3614 VGND VGND VPWR VPWR _06874_ sky130_fd_sc_hd__o311a_1
XFILLER_0_169_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23938_ _03800_ _03801_ VGND VGND VPWR VPWR _03802_ sky130_fd_sc_hd__and2b_1
XFILLER_0_192_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14671_ net4281 VGND VGND VPWR VPWR _06823_ sky130_fd_sc_hd__buf_1
XFILLER_0_169_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23869_ net1162 _03733_ VGND VGND VPWR VPWR _03734_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_129_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length7874 net7875 VGND VGND VPWR VPWR net7874 sky130_fd_sc_hd__buf_1
X_16410_ _08468_ _08470_ _08471_ VGND VGND VPWR VPWR _08472_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_168_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13622_ _05889_ net911 _05891_ VGND VGND VPWR VPWR _05892_ sky130_fd_sc_hd__and3_1
X_25608_ clknet_leaf_105_clk _00481_ net8358 VGND VGND VPWR VPWR cordic0.domain\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_17390_ net612 _09297_ _09295_ VGND VGND VPWR VPWR _09298_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_183_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16341_ _08325_ net1249 _08403_ VGND VGND VPWR VPWR _08404_ sky130_fd_sc_hd__a21o_1
X_13553_ net7671 net1150 VGND VGND VPWR VPWR _05824_ sky130_fd_sc_hd__nand2_1
X_25539_ clknet_leaf_32_clk _00419_ net8682 VGND VGND VPWR VPWR pid_q.prev_int\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout7012 net7018 VGND VGND VPWR VPWR net7012 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_27_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout7034 net7049 VGND VGND VPWR VPWR net7034 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19060_ _10819_ _10896_ VGND VGND VPWR VPWR _10897_ sky130_fd_sc_hd__xnor2_2
Xfanout6311 net6314 VGND VGND VPWR VPWR net6311 sky130_fd_sc_hd__buf_1
X_16272_ _08276_ _08281_ _08274_ VGND VGND VPWR VPWR _08336_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_82_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13484_ _05748_ _05756_ VGND VGND VPWR VPWR _05757_ sky130_fd_sc_hd__xor2_2
XFILLER_0_89_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6333 net6346 VGND VGND VPWR VPWR net6333 sky130_fd_sc_hd__clkbuf_1
Xwire7140 net7139 VGND VGND VPWR VPWR net7140 sky130_fd_sc_hd__buf_1
Xfanout6344 cordic0.vec\[0\]\[1\] VGND VGND VPWR VPWR net6344 sky130_fd_sc_hd__buf_1
X_18011_ _09636_ _09861_ VGND VGND VPWR VPWR _09862_ sky130_fd_sc_hd__nand2_1
Xfanout7089 net7093 VGND VGND VPWR VPWR net7089 sky130_fd_sc_hd__buf_1
X_15223_ _07292_ net1276 _07296_ VGND VGND VPWR VPWR _07297_ sky130_fd_sc_hd__o21ai_1
Xwire7151 matmul0.sin\[8\] VGND VGND VPWR VPWR net7151 sky130_fd_sc_hd__buf_1
Xwire7162 net7163 VGND VGND VPWR VPWR net7162 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout6377 net6380 VGND VGND VPWR VPWR net6377 sky130_fd_sc_hd__buf_1
Xwire7173 net7174 VGND VGND VPWR VPWR net7173 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7195 net7196 VGND VGND VPWR VPWR net7195 sky130_fd_sc_hd__clkbuf_1
Xwire6461 net6460 VGND VGND VPWR VPWR net6461 sky130_fd_sc_hd__buf_1
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15154_ _07026_ _07028_ net4169 net4164 VGND VGND VPWR VPWR _07228_ sky130_fd_sc_hd__o22a_1
Xfanout4920 net4924 VGND VGND VPWR VPWR net4920 sky130_fd_sc_hd__buf_1
Xwire6472 net6473 VGND VGND VPWR VPWR net6472 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_136_Right_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6483 net6484 VGND VGND VPWR VPWR net6483 sky130_fd_sc_hd__buf_1
X_14105_ _06323_ _06352_ _06354_ VGND VGND VPWR VPWR _06367_ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5760 net5761 VGND VGND VPWR VPWR net5760 sky130_fd_sc_hd__buf_1
Xwire5771 net5772 VGND VGND VPWR VPWR net5771 sky130_fd_sc_hd__clkbuf_1
X_19962_ net3153 _11755_ VGND VGND VPWR VPWR _11793_ sky130_fd_sc_hd__nand2_1
X_15085_ net2778 net2243 _07158_ VGND VGND VPWR VPWR _07159_ sky130_fd_sc_hd__o21ai_1
Xwire5782 net5777 VGND VGND VPWR VPWR net5782 sky130_fd_sc_hd__buf_1
Xwire5793 net5792 VGND VGND VPWR VPWR net5793 sky130_fd_sc_hd__buf_1
X_14036_ net7706 net1315 VGND VGND VPWR VPWR _06300_ sky130_fd_sc_hd__nand2_1
X_18913_ _10123_ _10371_ _10372_ net6832 net6859 VGND VGND VPWR VPWR _10753_ sky130_fd_sc_hd__o221a_1
X_19893_ _11720_ _11721_ _11725_ _11661_ net3858 VGND VGND VPWR VPWR _11726_ sky130_fd_sc_hd__a221oi_1
X_18844_ net2125 VGND VGND VPWR VPWR _10687_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18775_ net764 _10603_ VGND VGND VPWR VPWR _10619_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15987_ net2712 net4071 _08053_ _08054_ VGND VGND VPWR VPWR _08055_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_145_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17726_ net6506 _09585_ net8043 VGND VGND VPWR VPWR _09586_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14938_ _07011_ VGND VGND VPWR VPWR _07012_ sky130_fd_sc_hd__buf_1
XFILLER_0_171_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17657_ net4004 svm0.tA\[13\] VGND VGND VPWR VPWR _09537_ sky130_fd_sc_hd__nand2_1
XFILLER_0_188_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14869_ _06952_ VGND VGND VPWR VPWR _00205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16608_ matmul0.matmul_stage_inst.mult2\[11\] net276 net3471 VGND VGND VPWR VPWR
+ _08654_ sky130_fd_sc_hd__mux2_1
X_17588_ _09420_ _09424_ _09427_ net877 _09469_ VGND VGND VPWR VPWR _09470_ sky130_fd_sc_hd__o311a_1
X_19327_ net6199 net6276 VGND VGND VPWR VPWR _11164_ sky130_fd_sc_hd__nand2_1
X_16539_ net976 net879 _08596_ net1086 VGND VGND VPWR VPWR _08598_ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19258_ _10906_ _10889_ VGND VGND VPWR VPWR _11095_ sky130_fd_sc_hd__xor2_1
XFILLER_0_115_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18209_ net3239 net3238 _10058_ _10059_ VGND VGND VPWR VPWR _10060_ sky130_fd_sc_hd__a22o_1
XFILLER_0_171_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19189_ net6259 net6294 VGND VGND VPWR VPWR _11026_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21220_ _00938_ _00968_ VGND VGND VPWR VPWR _01236_ sky130_fd_sc_hd__nor2_1
Xhold101 svm0.tB\[1\] VGND VGND VPWR VPWR net9054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 matmul0.matmul_stage_inst.d\[9\] VGND VGND VPWR VPWR net9065 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 cordic0.sin\[9\] VGND VGND VPWR VPWR net9076 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_103_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold134 matmul0.matmul_stage_inst.d\[13\] VGND VGND VPWR VPWR net9087 sky130_fd_sc_hd__dlygate4sd3_1
X_21151_ _01153_ _01154_ VGND VGND VPWR VPWR _01167_ sky130_fd_sc_hd__xor2_1
Xhold145 cordic0.sin\[7\] VGND VGND VPWR VPWR net9098 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 pid_d.prev_int\[13\] VGND VGND VPWR VPWR net9109 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3109 net3110 VGND VGND VPWR VPWR net3109 sky130_fd_sc_hd__clkbuf_1
Xhold167 matmul0.matmul_stage_inst.b\[14\] VGND VGND VPWR VPWR net9120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 svm0.tA\[13\] VGND VGND VPWR VPWR net9131 sky130_fd_sc_hd__dlygate4sd3_1
X_20102_ _11911_ net420 VGND VGND VPWR VPWR _11930_ sky130_fd_sc_hd__or2_1
Xhold189 pid_q.prev_error\[8\] VGND VGND VPWR VPWR net9142 sky130_fd_sc_hd__dlygate4sd3_1
X_21082_ net5562 net5879 _01095_ _01068_ VGND VGND VPWR VPWR _01098_ sky130_fd_sc_hd__a211o_1
XFILLER_0_186_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2408 _03985_ VGND VGND VPWR VPWR net2408 sky130_fd_sc_hd__buf_1
XFILLER_0_10_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2419 _03388_ VGND VGND VPWR VPWR net2419 sky130_fd_sc_hd__buf_1
XFILLER_0_42_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24910_ _04699_ VGND VGND VPWR VPWR _04700_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20033_ _11860_ _11862_ VGND VGND VPWR VPWR _11863_ sky130_fd_sc_hd__xnor2_2
X_25890_ clknet_leaf_14_clk _00763_ net8621 VGND VGND VPWR VPWR pid_q.kp\[2\] sky130_fd_sc_hd__dfrtp_1
Xwire1707 _02206_ VGND VGND VPWR VPWR net1707 sky130_fd_sc_hd__clkbuf_1
Xwire1718 _01874_ VGND VGND VPWR VPWR net1718 sky130_fd_sc_hd__buf_1
Xwire1729 _01358_ VGND VGND VPWR VPWR net1729 sky130_fd_sc_hd__buf_1
X_24841_ net4916 net2008 net2001 net508 VGND VGND VPWR VPWR _00722_ sky130_fd_sc_hd__a22o_1
X_24772_ net5220 _04597_ _04598_ VGND VGND VPWR VPWR _04600_ sky130_fd_sc_hd__and3_1
X_21984_ net2068 _01885_ VGND VGND VPWR VPWR _01992_ sky130_fd_sc_hd__or2_1
Xmax_length7104 net7103 VGND VGND VPWR VPWR net7104 sky130_fd_sc_hd__buf_1
XFILLER_0_68_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23723_ net4600 net4942 VGND VGND VPWR VPWR _03589_ sky130_fd_sc_hd__nand2_1
X_20935_ _00903_ _00950_ VGND VGND VPWR VPWR _00951_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23654_ net5094 net4511 VGND VGND VPWR VPWR _03521_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20866_ net5802 VGND VGND VPWR VPWR _00882_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22605_ net7250 _02576_ VGND VGND VPWR VPWR _02579_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23585_ net1670 net1667 _03452_ VGND VGND VPWR VPWR _03453_ sky130_fd_sc_hd__o21ai_2
X_20797_ _00811_ _00812_ VGND VGND VPWR VPWR _00813_ sky130_fd_sc_hd__xor2_1
X_25324_ clknet_leaf_75_clk _00207_ net8464 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.f\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22536_ net9124 net1700 _02530_ VGND VGND VPWR VPWR _00540_ sky130_fd_sc_hd__a21o_1
XFILLER_0_134_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length613 _09282_ VGND VGND VPWR VPWR net613 sky130_fd_sc_hd__buf_1
XFILLER_0_180_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25255_ clknet_leaf_77_clk _00138_ net8437 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.b\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_22467_ net4297 _02463_ _02467_ net4379 VGND VGND VPWR VPWR _02468_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_161_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5001 net5002 VGND VGND VPWR VPWR net5001 sky130_fd_sc_hd__buf_1
X_24206_ _04058_ _04066_ VGND VGND VPWR VPWR _04067_ sky130_fd_sc_hd__xnor2_2
Xwire5012 net5013 VGND VGND VPWR VPWR net5012 sky130_fd_sc_hd__buf_1
X_21418_ _01430_ _01431_ VGND VGND VPWR VPWR _01432_ sky130_fd_sc_hd__nor2_1
Xwire5023 net5025 VGND VGND VPWR VPWR net5023 sky130_fd_sc_hd__buf_1
X_25186_ clknet_leaf_72_clk _00075_ net8662 VGND VGND VPWR VPWR matmul0.a_in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire5034 net5035 VGND VGND VPWR VPWR net5034 sky130_fd_sc_hd__buf_1
XFILLER_0_161_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22398_ _02397_ _02398_ VGND VGND VPWR VPWR _02400_ sky130_fd_sc_hd__nand2_1
Xwire5045 net5046 VGND VGND VPWR VPWR net5045 sky130_fd_sc_hd__clkbuf_1
Xwire4300 net4301 VGND VGND VPWR VPWR net4300 sky130_fd_sc_hd__buf_1
XFILLER_0_60_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4311 net4312 VGND VGND VPWR VPWR net4311 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24137_ _03996_ _03997_ VGND VGND VPWR VPWR _03999_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4322 net4323 VGND VGND VPWR VPWR net4322 sky130_fd_sc_hd__buf_1
X_21349_ _01361_ _01362_ VGND VGND VPWR VPWR _01363_ sky130_fd_sc_hd__xnor2_1
Xwire5078 net5079 VGND VGND VPWR VPWR net5078 sky130_fd_sc_hd__buf_1
Xwire4333 net4331 VGND VGND VPWR VPWR net4333 sky130_fd_sc_hd__buf_1
Xwire5089 net5090 VGND VGND VPWR VPWR net5089 sky130_fd_sc_hd__buf_1
Xwire4344 net4345 VGND VGND VPWR VPWR net4344 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3610 net3611 VGND VGND VPWR VPWR net3610 sky130_fd_sc_hd__clkbuf_2
Xwire4355 net4356 VGND VGND VPWR VPWR net4355 sky130_fd_sc_hd__clkbuf_1
Xwire4366 net4361 VGND VGND VPWR VPWR net4366 sky130_fd_sc_hd__buf_1
Xwire3621 _06823_ VGND VGND VPWR VPWR net3621 sky130_fd_sc_hd__dlymetal6s2s_1
X_24068_ _03930_ VGND VGND VPWR VPWR _03931_ sky130_fd_sc_hd__inv_2
Xwire3632 net3634 VGND VGND VPWR VPWR net3632 sky130_fd_sc_hd__buf_1
Xwire4377 net4378 VGND VGND VPWR VPWR net4377 sky130_fd_sc_hd__clkbuf_1
Xwire3643 net3644 VGND VGND VPWR VPWR net3643 sky130_fd_sc_hd__buf_1
Xwire3654 net3655 VGND VGND VPWR VPWR net3654 sky130_fd_sc_hd__clkbuf_1
Xwire4399 pid_q.out\[14\] VGND VGND VPWR VPWR net4399 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23019_ _02875_ _02888_ VGND VGND VPWR VPWR _02889_ sky130_fd_sc_hd__xnor2_2
Xwire2920 net2921 VGND VGND VPWR VPWR net2920 sky130_fd_sc_hd__clkbuf_1
Xwire3665 _06510_ VGND VGND VPWR VPWR net3665 sky130_fd_sc_hd__clkbuf_1
X_15910_ _07871_ _07876_ _07978_ VGND VGND VPWR VPWR _07979_ sky130_fd_sc_hd__o21a_1
Xwire2931 _06511_ VGND VGND VPWR VPWR net2931 sky130_fd_sc_hd__buf_2
XFILLER_0_194_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3687 _05053_ VGND VGND VPWR VPWR net3687 sky130_fd_sc_hd__buf_1
X_16890_ net6390 net6368 VGND VGND VPWR VPWR _08854_ sky130_fd_sc_hd__and2b_1
Xwire2942 net2943 VGND VGND VPWR VPWR net2942 sky130_fd_sc_hd__buf_1
Xwire2953 net2954 VGND VGND VPWR VPWR net2953 sky130_fd_sc_hd__clkbuf_1
Xwire2964 net2965 VGND VGND VPWR VPWR net2964 sky130_fd_sc_hd__buf_1
Xwire2975 _04958_ VGND VGND VPWR VPWR net2975 sky130_fd_sc_hd__buf_1
X_15841_ _07802_ _07817_ _07910_ VGND VGND VPWR VPWR _07911_ sky130_fd_sc_hd__o21ai_2
Xwire2986 net2987 VGND VGND VPWR VPWR net2986 sky130_fd_sc_hd__buf_1
Xwire2997 net2998 VGND VGND VPWR VPWR net2997 sky130_fd_sc_hd__buf_1
XFILLER_0_188_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18560_ _10384_ net1436 _10386_ VGND VGND VPWR VPWR _10408_ sky130_fd_sc_hd__a21boi_1
X_12984_ net7688 net2977 net2335 VGND VGND VPWR VPWR _05257_ sky130_fd_sc_hd__and3_1
X_15772_ net2700 _07841_ VGND VGND VPWR VPWR _07842_ sky130_fd_sc_hd__nand2_1
X_17511_ net3271 _09397_ VGND VGND VPWR VPWR _09398_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14723_ net4224 VGND VGND VPWR VPWR _06862_ sky130_fd_sc_hd__clkbuf_1
X_18491_ _10334_ _10340_ VGND VGND VPWR VPWR _10341_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17442_ net6738 VGND VGND VPWR VPWR _09339_ sky130_fd_sc_hd__inv_2
X_14654_ net8970 _06801_ _06811_ VGND VGND VPWR VPWR _00131_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13605_ net7723 net2307 net1952 VGND VGND VPWR VPWR _05875_ sky130_fd_sc_hd__and3_1
XFILLER_0_145_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17373_ net7377 svm0.delta\[1\] net6743 VGND VGND VPWR VPWR _09284_ sky130_fd_sc_hd__or3_1
X_14585_ _06753_ _06758_ _06759_ VGND VGND VPWR VPWR _06760_ sky130_fd_sc_hd__o21a_1
XFILLER_0_184_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19112_ net3189 _10945_ _10947_ _10948_ VGND VGND VPWR VPWR _10949_ sky130_fd_sc_hd__o211ai_1
X_13536_ _05743_ _05757_ _05741_ VGND VGND VPWR VPWR _05807_ sky130_fd_sc_hd__o21ba_1
X_16324_ net2791 net2639 VGND VGND VPWR VPWR _08387_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19043_ net6187 net6229 VGND VGND VPWR VPWR _10880_ sky130_fd_sc_hd__xor2_2
X_16255_ net2751 net2643 VGND VGND VPWR VPWR _08319_ sky130_fd_sc_hd__nor2_2
X_13467_ net912 net997 VGND VGND VPWR VPWR _05740_ sky130_fd_sc_hd__xor2_1
XFILLER_0_153_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15206_ _07253_ _07279_ VGND VGND VPWR VPWR _07280_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_140_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout6185 net6191 VGND VGND VPWR VPWR net6185 sky130_fd_sc_hd__buf_1
XFILLER_0_3_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16186_ net3492 net2645 net3522 net1849 VGND VGND VPWR VPWR _08251_ sky130_fd_sc_hd__and4_1
X_13398_ _05669_ _05670_ _05661_ VGND VGND VPWR VPWR _05671_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15137_ net1894 _07181_ _07210_ VGND VGND VPWR VPWR _07211_ sky130_fd_sc_hd__a21o_1
Xfanout4761 pid_q.mult0.a\[1\] VGND VGND VPWR VPWR net4761 sky130_fd_sc_hd__clkbuf_1
Xwire5590 net5591 VGND VGND VPWR VPWR net5590 sky130_fd_sc_hd__clkbuf_1
X_15068_ net3486 VGND VGND VPWR VPWR _07142_ sky130_fd_sc_hd__buf_1
X_19945_ _11774_ _11776_ VGND VGND VPWR VPWR _11777_ sky130_fd_sc_hd__nand2_1
X_14019_ _06234_ _06242_ net835 VGND VGND VPWR VPWR _06283_ sky130_fd_sc_hd__o21a_1
X_19876_ _11705_ _11707_ VGND VGND VPWR VPWR _11709_ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18827_ _10276_ _10638_ _10669_ net6855 VGND VGND VPWR VPWR _10670_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18758_ _10601_ _10602_ VGND VGND VPWR VPWR _10603_ sky130_fd_sc_hd__and2_1
XFILLER_0_172_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17709_ pid_q.prev_int\[0\] net1218 net1452 net5184 VGND VGND VPWR VPWR _00414_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18689_ net6877 net6896 net6975 VGND VGND VPWR VPWR _10535_ sky130_fd_sc_hd__mux2_1
X_20720_ net6023 _12481_ VGND VGND VPWR VPWR _12492_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20651_ net1738 _12419_ VGND VGND VPWR VPWR _12429_ sky130_fd_sc_hd__or2_1
XFILLER_0_191_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7909 net7910 VGND VGND VPWR VPWR net7909 sky130_fd_sc_hd__buf_1
XFILLER_0_74_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23370_ _03232_ _03234_ _03239_ VGND VGND VPWR VPWR _03240_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20582_ net2594 _12363_ _12364_ _09008_ _12353_ VGND VGND VPWR VPWR _12365_ sky130_fd_sc_hd__o221a_1
XFILLER_0_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22321_ _02279_ net552 VGND VGND VPWR VPWR _02325_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25040_ net1628 _04791_ net2147 VGND VGND VPWR VPWR _04792_ sky130_fd_sc_hd__a21o_1
X_22252_ pid_d.prev_error\[11\] net5966 VGND VGND VPWR VPWR _02257_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21203_ _01114_ _01116_ _01218_ VGND VGND VPWR VPWR _01219_ sky130_fd_sc_hd__a21oi_1
X_22183_ _02162_ net859 VGND VGND VPWR VPWR _02188_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_52_Left_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21134_ net5583 net5952 VGND VGND VPWR VPWR _01150_ sky130_fd_sc_hd__nand2_1
Xclkbuf_2_2_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2_0_clk sky130_fd_sc_hd__clkbuf_8
Xwire2216 _07896_ VGND VGND VPWR VPWR net2216 sky130_fd_sc_hd__clkbuf_1
Xwire2227 _07607_ VGND VGND VPWR VPWR net2227 sky130_fd_sc_hd__buf_1
X_21065_ net5564 net5929 VGND VGND VPWR VPWR _01081_ sky130_fd_sc_hd__nand2_1
Xwire2238 net2241 VGND VGND VPWR VPWR net2238 sky130_fd_sc_hd__buf_1
Xwire1504 net1505 VGND VGND VPWR VPWR net1504 sky130_fd_sc_hd__buf_1
Xwire2249 _07130_ VGND VGND VPWR VPWR net2249 sky130_fd_sc_hd__buf_1
Xwire1515 _08106_ VGND VGND VPWR VPWR net1515 sky130_fd_sc_hd__clkbuf_2
X_20016_ _11812_ _11845_ _11816_ VGND VGND VPWR VPWR _11846_ sky130_fd_sc_hd__o21ai_4
Xwire1526 _07950_ VGND VGND VPWR VPWR net1526 sky130_fd_sc_hd__buf_1
X_25873_ clknet_leaf_17_clk _00746_ net8626 VGND VGND VPWR VPWR pid_q.ki\[1\] sky130_fd_sc_hd__dfrtp_1
Xwire1537 _07678_ VGND VGND VPWR VPWR net1537 sky130_fd_sc_hd__buf_1
Xwire1548 net1550 VGND VGND VPWR VPWR net1548 sky130_fd_sc_hd__buf_1
Xwire1559 _06509_ VGND VGND VPWR VPWR net1559 sky130_fd_sc_hd__buf_1
X_24824_ net7482 net1011 net2419 VGND VGND VPWR VPWR _04645_ sky130_fd_sc_hd__a21o_1
XFILLER_0_193_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24755_ pid_q.curr_error\[7\] net1369 net1366 net737 VGND VGND VPWR VPWR _00704_
+ sky130_fd_sc_hd__a22o_1
X_21967_ net2065 _01876_ VGND VGND VPWR VPWR _01975_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_61_Left_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length6211 net6206 VGND VGND VPWR VPWR net6211 sky130_fd_sc_hd__clkbuf_1
X_23706_ _03571_ _03572_ VGND VGND VPWR VPWR _03573_ sky130_fd_sc_hd__nand2_1
X_20918_ _00931_ _00933_ VGND VGND VPWR VPWR _00934_ sky130_fd_sc_hd__xor2_1
X_24686_ net9067 _04507_ _04525_ VGND VGND VPWR VPWR _00695_ sky130_fd_sc_hd__a21o_1
XFILLER_0_167_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21898_ _01827_ _01906_ VGND VGND VPWR VPWR _01907_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23637_ _03417_ _03419_ _03415_ VGND VGND VPWR VPWR _03504_ sky130_fd_sc_hd__a21bo_1
X_20849_ _12526_ _12528_ VGND VGND VPWR VPWR _00865_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14370_ _06580_ matmul0.a_in\[11\] net899 VGND VGND VPWR VPWR _06581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23568_ _03434_ _03435_ VGND VGND VPWR VPWR _03436_ sky130_fd_sc_hd__xnor2_1
Xwire801 _02595_ VGND VGND VPWR VPWR net801 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4864 net4865 VGND VGND VPWR VPWR net4864 sky130_fd_sc_hd__buf_1
XFILLER_0_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire812 net813 VGND VGND VPWR VPWR net812 sky130_fd_sc_hd__clkbuf_1
X_13321_ _05592_ _05593_ VGND VGND VPWR VPWR _05594_ sky130_fd_sc_hd__xor2_1
X_25307_ clknet_leaf_71_clk _00190_ net8461 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.e\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire823 net824 VGND VGND VPWR VPWR net823 sky130_fd_sc_hd__buf_1
Xwire834 _06373_ VGND VGND VPWR VPWR net834 sky130_fd_sc_hd__buf_1
X_22519_ _02518_ VGND VGND VPWR VPWR _02519_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire845 _05576_ VGND VGND VPWR VPWR net845 sky130_fd_sc_hd__buf_1
X_23499_ _03363_ _03367_ VGND VGND VPWR VPWR _03368_ sky130_fd_sc_hd__xnor2_2
Xwire856 net857 VGND VGND VPWR VPWR net856 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire867 _12012_ VGND VGND VPWR VPWR net867 sky130_fd_sc_hd__buf_1
X_16040_ _07929_ net1260 net2700 VGND VGND VPWR VPWR _08107_ sky130_fd_sc_hd__a21o_1
X_25238_ clknet_leaf_32_clk net2384 net8683 VGND VGND VPWR VPWR pid_q.state\[5\] sky130_fd_sc_hd__dfrtp_1
X_13252_ net7879 net1948 _05413_ _05414_ VGND VGND VPWR VPWR _05525_ sky130_fd_sc_hd__a22o_1
Xwire878 _08940_ VGND VGND VPWR VPWR net878 sky130_fd_sc_hd__buf_1
XFILLER_0_49_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire889 _07592_ VGND VGND VPWR VPWR net889 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_70_Left_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25169_ clknet_leaf_54_clk _00058_ net8729 VGND VGND VPWR VPWR svm0.periodTop\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13183_ _05366_ _05367_ _05455_ VGND VGND VPWR VPWR _05456_ sky130_fd_sc_hd__o21a_1
Xwire4130 net4131 VGND VGND VPWR VPWR net4130 sky130_fd_sc_hd__buf_1
Xwire4141 net4142 VGND VGND VPWR VPWR net4141 sky130_fd_sc_hd__clkbuf_1
Xwire4152 _07014_ VGND VGND VPWR VPWR net4152 sky130_fd_sc_hd__clkbuf_1
X_17991_ _09673_ _09776_ _09841_ VGND VGND VPWR VPWR _09842_ sky130_fd_sc_hd__a21o_1
Xwire4163 _07009_ VGND VGND VPWR VPWR net4163 sky130_fd_sc_hd__buf_1
XFILLER_0_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4174 _07000_ VGND VGND VPWR VPWR net4174 sky130_fd_sc_hd__buf_1
Xwire3440 net3441 VGND VGND VPWR VPWR net3440 sky130_fd_sc_hd__buf_1
Xwire4185 net4187 VGND VGND VPWR VPWR net4185 sky130_fd_sc_hd__buf_1
X_19730_ _11508_ _11562_ _11503_ VGND VGND VPWR VPWR _11565_ sky130_fd_sc_hd__a21oi_1
Xwire3451 net3452 VGND VGND VPWR VPWR net3451 sky130_fd_sc_hd__buf_1
XFILLER_0_159_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16942_ net7138 net1506 VGND VGND VPWR VPWR _08906_ sky130_fd_sc_hd__xnor2_1
Xwire4196 _06982_ VGND VGND VPWR VPWR net4196 sky130_fd_sc_hd__buf_1
Xwire3462 _07189_ VGND VGND VPWR VPWR net3462 sky130_fd_sc_hd__buf_1
Xwire3484 net3485 VGND VGND VPWR VPWR net3484 sky130_fd_sc_hd__clkbuf_1
Xwire3495 _07107_ VGND VGND VPWR VPWR net3495 sky130_fd_sc_hd__buf_1
Xwire2750 net2751 VGND VGND VPWR VPWR net2750 sky130_fd_sc_hd__dlymetal6s2s_1
X_19661_ net6045 _11495_ _11496_ VGND VGND VPWR VPWR _11497_ sky130_fd_sc_hd__a21oi_1
Xwire2761 net2762 VGND VGND VPWR VPWR net2761 sky130_fd_sc_hd__dlymetal6s2s_1
X_16873_ net2189 _08837_ net6460 VGND VGND VPWR VPWR _08838_ sky130_fd_sc_hd__mux2_1
Xwire2772 net2773 VGND VGND VPWR VPWR net2772 sky130_fd_sc_hd__buf_2
Xwire2783 net2784 VGND VGND VPWR VPWR net2783 sky130_fd_sc_hd__buf_1
Xwire2794 net2795 VGND VGND VPWR VPWR net2794 sky130_fd_sc_hd__buf_1
X_18612_ net6377 net422 _10458_ VGND VGND VPWR VPWR _10460_ sky130_fd_sc_hd__nand3_1
X_15824_ _07794_ _07796_ _07893_ VGND VGND VPWR VPWR _07894_ sky130_fd_sc_hd__a21oi_2
X_19592_ _11373_ _11427_ _11428_ VGND VGND VPWR VPWR _11429_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18543_ net3925 _10389_ _10390_ _10391_ VGND VGND VPWR VPWR _10392_ sky130_fd_sc_hd__a211oi_1
X_12967_ _05227_ _05228_ _05235_ _05239_ VGND VGND VPWR VPWR _05240_ sky130_fd_sc_hd__a211o_1
X_15755_ _07823_ _07824_ _07825_ VGND VGND VPWR VPWR _07826_ sky130_fd_sc_hd__or3_1
XFILLER_0_59_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14706_ net9039 net2862 net2262 net1547 VGND VGND VPWR VPWR _00145_ sky130_fd_sc_hd__a22o_1
X_18474_ _10243_ net1773 VGND VGND VPWR VPWR _10324_ sky130_fd_sc_hd__and2b_1
XFILLER_0_129_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12898_ net7727 net2344 net2341 VGND VGND VPWR VPWR _05171_ sky130_fd_sc_hd__and3_1
X_15686_ net1536 _07756_ VGND VGND VPWR VPWR _07757_ sky130_fd_sc_hd__xor2_1
XFILLER_0_185_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17425_ svm0.delta\[12\] net6742 _09320_ VGND VGND VPWR VPWR _09325_ sky130_fd_sc_hd__or3_1
XFILLER_0_158_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14637_ net3697 VGND VGND VPWR VPWR _06802_ sky130_fd_sc_hd__buf_1
XFILLER_0_142_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17356_ svm0.rising net771 net1796 VGND VGND VPWR VPWR _09269_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14568_ net5223 net3640 _06731_ _06730_ net7260 VGND VGND VPWR VPWR _06745_ sky130_fd_sc_hd__o32a_1
XFILLER_0_172_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16307_ matmul0.matmul_stage_inst.mult1\[10\] net247 net3478 VGND VGND VPWR VPWR
+ _08371_ sky130_fd_sc_hd__mux2_1
X_13519_ _05701_ _05702_ net7814 net1586 VGND VGND VPWR VPWR _05790_ sky130_fd_sc_hd__o211a_1
X_17287_ net6700 net6684 net6688 _09201_ VGND VGND VPWR VPWR _09202_ sky130_fd_sc_hd__or4_1
X_14499_ _06680_ _06681_ VGND VGND VPWR VPWR _06682_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19026_ net2528 _10832_ net3214 VGND VGND VPWR VPWR _10863_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16238_ net491 _08301_ VGND VGND VPWR VPWR _08303_ sky130_fd_sc_hd__or2_1
XFILLER_0_180_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16169_ net386 _08159_ _08158_ VGND VGND VPWR VPWR _08235_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_167_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19928_ _11755_ _11759_ VGND VGND VPWR VPWR _11760_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19859_ _11686_ _11691_ VGND VGND VPWR VPWR _11692_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_183_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22870_ net5363 _02766_ net3066 VGND VGND VPWR VPWR _02767_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21821_ _01749_ _01751_ _01750_ VGND VGND VPWR VPWR _01830_ sky130_fd_sc_hd__o21a_1
XFILLER_0_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24540_ _04264_ _04374_ _04375_ VGND VGND VPWR VPWR _04396_ sky130_fd_sc_hd__a21bo_1
X_21752_ _01753_ _01761_ VGND VGND VPWR VPWR _01762_ sky130_fd_sc_hd__xnor2_1
X_20703_ _12142_ _12476_ net8060 VGND VGND VPWR VPWR _12477_ sky130_fd_sc_hd__o21ai_1
X_24471_ net5175 net3757 net2433 _04328_ VGND VGND VPWR VPWR _00677_ sky130_fd_sc_hd__a22o_1
X_21683_ _01690_ _01693_ VGND VGND VPWR VPWR _01694_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8407 net8405 VGND VGND VPWR VPWR net8407 sky130_fd_sc_hd__buf_1
XFILLER_0_148_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8418 net8419 VGND VGND VPWR VPWR net8418 sky130_fd_sc_hd__buf_1
XFILLER_0_148_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23422_ _03289_ _03291_ VGND VGND VPWR VPWR _03292_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7706 net7707 VGND VGND VPWR VPWR net7706 sky130_fd_sc_hd__buf_1
X_20634_ net2190 _12413_ net8054 VGND VGND VPWR VPWR _12414_ sky130_fd_sc_hd__o21a_1
Xwire7728 net7733 VGND VGND VPWR VPWR net7728 sky130_fd_sc_hd__buf_1
XFILLER_0_11_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3415 net3416 VGND VGND VPWR VPWR net3415 sky130_fd_sc_hd__buf_1
Xwire7739 net7740 VGND VGND VPWR VPWR net7739 sky130_fd_sc_hd__clkbuf_1
X_23353_ _02940_ _02942_ _03222_ VGND VGND VPWR VPWR _03223_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_46_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20565_ _12333_ _12336_ _12344_ net2516 VGND VGND VPWR VPWR _12349_ sky130_fd_sc_hd__a31o_1
Xmax_length3448 net3449 VGND VGND VPWR VPWR net3448 sky130_fd_sc_hd__buf_1
XFILLER_0_190_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3459 net3460 VGND VGND VPWR VPWR net3459 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22304_ net5380 net2051 VGND VGND VPWR VPWR _02308_ sky130_fd_sc_hd__nand2_1
X_23284_ _03107_ _03110_ _03153_ VGND VGND VPWR VPWR _03154_ sky130_fd_sc_hd__a21o_1
X_20496_ net2086 _12283_ VGND VGND VPWR VPWR _12284_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25023_ _04774_ _04775_ VGND VGND VPWR VPWR _04777_ sky130_fd_sc_hd__or2_1
X_22235_ net2058 net943 VGND VGND VPWR VPWR _02240_ sky130_fd_sc_hd__xnor2_2
X_22166_ _02115_ _02171_ VGND VGND VPWR VPWR _02172_ sky130_fd_sc_hd__xnor2_1
Xwire2002 net2003 VGND VGND VPWR VPWR net2002 sky130_fd_sc_hd__clkbuf_1
X_21117_ _01130_ _01132_ VGND VGND VPWR VPWR _01133_ sky130_fd_sc_hd__and2b_1
Xwire2013 net2014 VGND VGND VPWR VPWR net2013 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2024 net2025 VGND VGND VPWR VPWR net2024 sky130_fd_sc_hd__buf_2
X_22097_ _02102_ _02103_ VGND VGND VPWR VPWR _02104_ sky130_fd_sc_hd__nand2_1
Xwire2035 net2036 VGND VGND VPWR VPWR net2035 sky130_fd_sc_hd__buf_1
Xwire1312 _05730_ VGND VGND VPWR VPWR net1312 sky130_fd_sc_hd__buf_1
Xwire2057 net2058 VGND VGND VPWR VPWR net2057 sky130_fd_sc_hd__clkbuf_2
X_25925_ clknet_leaf_1_clk _00798_ net8404 VGND VGND VPWR VPWR pid_d.prev_int\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_21048_ _01060_ _01063_ _01058_ VGND VGND VPWR VPWR _01064_ sky130_fd_sc_hd__mux2_1
Xwire1323 net1324 VGND VGND VPWR VPWR net1323 sky130_fd_sc_hd__buf_1
Xwire1334 net1335 VGND VGND VPWR VPWR net1334 sky130_fd_sc_hd__clkbuf_1
Xwire2079 net2080 VGND VGND VPWR VPWR net2079 sky130_fd_sc_hd__clkbuf_2
Xwire1345 _04967_ VGND VGND VPWR VPWR net1345 sky130_fd_sc_hd__clkbuf_1
Xwire1356 _04902_ VGND VGND VPWR VPWR net1356 sky130_fd_sc_hd__buf_1
X_13870_ _06091_ _06136_ VGND VGND VPWR VPWR _06137_ sky130_fd_sc_hd__xnor2_2
X_25856_ clknet_leaf_19_clk _00729_ net8624 VGND VGND VPWR VPWR pid_q.mult0.a\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1367 _04543_ VGND VGND VPWR VPWR net1367 sky130_fd_sc_hd__buf_1
Xwire1378 _04508_ VGND VGND VPWR VPWR net1378 sky130_fd_sc_hd__buf_1
Xwire1389 _02121_ VGND VGND VPWR VPWR net1389 sky130_fd_sc_hd__buf_1
X_12821_ net7759 _04919_ VGND VGND VPWR VPWR _05094_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24807_ _04628_ _04630_ VGND VGND VPWR VPWR _04631_ sky130_fd_sc_hd__xnor2_1
X_22999_ net7524 net7500 net7464 _02868_ net8865 VGND VGND VPWR VPWR _02869_ sky130_fd_sc_hd__o311a_1
X_25787_ clknet_leaf_64_clk _00660_ net8663 VGND VGND VPWR VPWR matmul0.beta_pass\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_12752_ net1155 _05024_ VGND VGND VPWR VPWR _05025_ sky130_fd_sc_hd__nand2_1
X_15540_ net2806 net3557 VGND VGND VPWR VPWR _07613_ sky130_fd_sc_hd__nor2_2
X_24738_ net5265 VGND VGND VPWR VPWR _04570_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15471_ net1875 _07544_ VGND VGND VPWR VPWR _07545_ sky130_fd_sc_hd__and2_1
X_24669_ pid_q.curr_error\[6\] net2383 net1373 VGND VGND VPWR VPWR _04517_ sky130_fd_sc_hd__and3_1
X_12683_ net7283 _04856_ net4278 VGND VGND VPWR VPWR _04956_ sky130_fd_sc_hd__nand3_1
X_17210_ _09159_ VGND VGND VPWR VPWR _00339_ sky130_fd_sc_hd__clkbuf_1
X_14422_ _06620_ matmul0.b_in\[7\] net895 VGND VGND VPWR VPWR _06621_ sky130_fd_sc_hd__mux2_1
Xwire8930 net8931 VGND VGND VPWR VPWR net8930 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18190_ net6892 _10040_ VGND VGND VPWR VPWR _10041_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_71_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8941 net8942 VGND VGND VPWR VPWR net8941 sky130_fd_sc_hd__clkbuf_1
Xwire8952 net100 VGND VGND VPWR VPWR net8952 sky130_fd_sc_hd__clkbuf_1
Xmax_length5384 net5385 VGND VGND VPWR VPWR net5384 sky130_fd_sc_hd__buf_1
XFILLER_0_126_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17141_ net6484 net3325 VGND VGND VPWR VPWR _09095_ sky130_fd_sc_hd__nor2_1
X_14353_ net7280 _06522_ net2900 net5355 _06566_ VGND VGND VPWR VPWR _06567_ sky130_fd_sc_hd__a221o_1
Xwire620 _08714_ VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__clkbuf_1
Xwire631 net632 VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__buf_1
Xwire642 net643 VGND VGND VPWR VPWR net642 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13304_ net7640 net1972 net1969 VGND VGND VPWR VPWR _05577_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire653 net654 VGND VGND VPWR VPWR net653 sky130_fd_sc_hd__buf_1
X_17072_ net3332 _09028_ net3342 _09029_ VGND VGND VPWR VPWR _09030_ sky130_fd_sc_hd__a22o_1
Xwire664 net665 VGND VGND VPWR VPWR net664 sky130_fd_sc_hd__clkbuf_1
X_14284_ net3649 VGND VGND VPWR VPWR _06518_ sky130_fd_sc_hd__clkbuf_2
Xwire675 _07555_ VGND VGND VPWR VPWR net675 sky130_fd_sc_hd__buf_1
Xmax_length3971 _09696_ VGND VGND VPWR VPWR net3971 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire686 net687 VGND VGND VPWR VPWR net686 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire697 _03174_ VGND VGND VPWR VPWR net697 sky130_fd_sc_hd__clkbuf_1
X_13235_ _05506_ _05507_ VGND VGND VPWR VPWR _05508_ sky130_fd_sc_hd__xnor2_1
X_16023_ net425 _08088_ _08089_ _08081_ VGND VGND VPWR VPWR _08090_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_126_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13166_ _05436_ _05437_ _05434_ _05435_ VGND VGND VPWR VPWR _05439_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_62_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13097_ _05366_ _05369_ VGND VGND VPWR VPWR _05370_ sky130_fd_sc_hd__xnor2_1
X_17974_ net3977 _09664_ VGND VGND VPWR VPWR _09825_ sky130_fd_sc_hd__or2_1
Xwire3270 _09575_ VGND VGND VPWR VPWR net3270 sky130_fd_sc_hd__buf_1
X_19713_ net6382 net6386 VGND VGND VPWR VPWR _11549_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_108_Left_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16925_ net6418 _08884_ net6419 _08885_ _08888_ VGND VGND VPWR VPWR _08889_ sky130_fd_sc_hd__o221a_1
Xwire3281 net3283 VGND VGND VPWR VPWR net3281 sky130_fd_sc_hd__buf_1
Xwire3292 net3293 VGND VGND VPWR VPWR net3292 sky130_fd_sc_hd__buf_1
Xwire2580 net2581 VGND VGND VPWR VPWR net2580 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2591 net2594 VGND VGND VPWR VPWR net2591 sky130_fd_sc_hd__clkbuf_1
X_19644_ _11429_ _11480_ VGND VGND VPWR VPWR _11481_ sky130_fd_sc_hd__nand2_1
X_16856_ net6092 net6061 net6501 VGND VGND VPWR VPWR _08821_ sky130_fd_sc_hd__mux2_1
X_15807_ _07871_ _07876_ VGND VGND VPWR VPWR _07877_ sky130_fd_sc_hd__xor2_1
Xwire1890 net1891 VGND VGND VPWR VPWR net1890 sky130_fd_sc_hd__clkbuf_1
X_19575_ _11408_ _11411_ VGND VGND VPWR VPWR _11412_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16787_ _08783_ VGND VGND VPWR VPWR _00292_ sky130_fd_sc_hd__clkbuf_1
X_13999_ _06260_ _06263_ VGND VGND VPWR VPWR _06264_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18526_ net6833 _10370_ _10373_ _10374_ VGND VGND VPWR VPWR _10375_ sky130_fd_sc_hd__a31o_1
XFILLER_0_153_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15738_ _07647_ _07649_ _07808_ VGND VGND VPWR VPWR _07809_ sky130_fd_sc_hd__o21a_1
XFILLER_0_87_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18457_ net1766 net1440 VGND VGND VPWR VPWR _10307_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15669_ matmul0.matmul_stage_inst.mult1\[2\] net433 net2678 VGND VGND VPWR VPWR _07741_
+ sky130_fd_sc_hd__mux2_1
X_17408_ svm0.delta\[9\] _09308_ VGND VGND VPWR VPWR _09312_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_117_Left_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18388_ net3986 net7014 net7098 VGND VGND VPWR VPWR _10239_ sky130_fd_sc_hd__and3_1
XFILLER_0_172_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17339_ _09213_ _09251_ _09252_ VGND VGND VPWR VPWR _09253_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20350_ _12150_ _12151_ VGND VGND VPWR VPWR _12152_ sky130_fd_sc_hd__or2b_1
XFILLER_0_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19009_ net6292 net6313 VGND VGND VPWR VPWR _10846_ sky130_fd_sc_hd__or2_1
XFILLER_0_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20281_ cordic0.slte0.opA\[0\] net1556 VGND VGND VPWR VPWR _12088_ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22020_ net5513 net5669 VGND VGND VPWR VPWR _02027_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_126_Left_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold16 matmul0.matmul_stage_inst.a\[4\] VGND VGND VPWR VPWR net8969 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold27 matmul0.matmul_stage_inst.b\[0\] VGND VGND VPWR VPWR net8980 sky130_fd_sc_hd__dlygate4sd3_1
X_23971_ net1161 _03834_ VGND VGND VPWR VPWR _03835_ sky130_fd_sc_hd__xnor2_2
Xhold38 matmul0.matmul_stage_inst.b\[13\] VGND VGND VPWR VPWR net8991 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold49 matmul0.matmul_stage_inst.d\[6\] VGND VGND VPWR VPWR net9002 sky130_fd_sc_hd__dlygate4sd3_1
X_25710_ clknet_leaf_9_clk _00583_ net8552 VGND VGND VPWR VPWR pid_d.mult0.a\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_22922_ net5975 _02812_ VGND VGND VPWR VPWR _02813_ sky130_fd_sc_hd__or2_1
X_25641_ clknet_leaf_103_clk _00514_ net8376 VGND VGND VPWR VPWR cordic0.vec\[0\]\[13\]
+ sky130_fd_sc_hd__dfstp_1
X_22853_ net5981 _02747_ pid_d.out\[4\] VGND VGND VPWR VPWR _02751_ sky130_fd_sc_hd__a21o_1
X_21804_ _01812_ _01813_ VGND VGND VPWR VPWR _01814_ sky130_fd_sc_hd__nand2_1
X_25572_ clknet_leaf_97_clk _00445_ net8398 VGND VGND VPWR VPWR cordic0.sin\[6\] sky130_fd_sc_hd__dfrtp_1
X_22784_ pid_d.kp\[4\] _02670_ net1680 VGND VGND VPWR VPWR _02700_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24523_ _04378_ _04379_ _04267_ VGND VGND VPWR VPWR _04380_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_135_Left_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21735_ _01658_ _01685_ _01672_ VGND VGND VPWR VPWR _01745_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_164_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8204 net8205 VGND VGND VPWR VPWR net8204 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8215 net8216 VGND VGND VPWR VPWR net8215 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24454_ _04227_ net1012 _04199_ VGND VGND VPWR VPWR _04312_ sky130_fd_sc_hd__o21ba_1
Xwire8226 net8227 VGND VGND VPWR VPWR net8226 sky130_fd_sc_hd__clkbuf_1
X_21666_ _01673_ _01676_ VGND VGND VPWR VPWR _01677_ sky130_fd_sc_hd__xnor2_2
Xwire8237 net8238 VGND VGND VPWR VPWR net8237 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7503 net7504 VGND VGND VPWR VPWR net7503 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8248 net8249 VGND VGND VPWR VPWR net8248 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7514 net7515 VGND VGND VPWR VPWR net7514 sky130_fd_sc_hd__clkbuf_1
Xwire8259 net8260 VGND VGND VPWR VPWR net8259 sky130_fd_sc_hd__clkbuf_1
Xfanout6718 svm0.counter\[6\] VGND VGND VPWR VPWR net6718 sky130_fd_sc_hd__buf_1
X_23405_ _03273_ _03274_ VGND VGND VPWR VPWR _03275_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_164_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20617_ net1226 _12397_ VGND VGND VPWR VPWR _12398_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24385_ _04240_ net929 VGND VGND VPWR VPWR _04244_ sky130_fd_sc_hd__nand2_1
Xwire7536 net7537 VGND VGND VPWR VPWR net7536 sky130_fd_sc_hd__clkbuf_1
Xwire7547 svm0.vC\[11\] VGND VGND VPWR VPWR net7547 sky130_fd_sc_hd__clkbuf_1
X_21597_ net3806 _01608_ VGND VGND VPWR VPWR _01609_ sky130_fd_sc_hd__and2_1
Xwire7558 matmul0.b_in\[14\] VGND VGND VPWR VPWR net7558 sky130_fd_sc_hd__clkbuf_1
Xmax_length2500 net2501 VGND VGND VPWR VPWR net2500 sky130_fd_sc_hd__buf_1
Xwire6813 net6814 VGND VGND VPWR VPWR net6813 sky130_fd_sc_hd__buf_1
Xwire6824 net6819 VGND VGND VPWR VPWR net6824 sky130_fd_sc_hd__buf_1
Xwire7569 net7570 VGND VGND VPWR VPWR net7569 sky130_fd_sc_hd__clkbuf_1
X_23336_ _02933_ _02935_ _02934_ VGND VGND VPWR VPWR _03206_ sky130_fd_sc_hd__o21ai_1
Xwire6835 net6836 VGND VGND VPWR VPWR net6835 sky130_fd_sc_hd__clkbuf_1
X_20548_ _12325_ _12327_ _12328_ _12332_ VGND VGND VPWR VPWR _12333_ sky130_fd_sc_hd__nand4_2
Xwire6846 net6847 VGND VGND VPWR VPWR net6846 sky130_fd_sc_hd__buf_1
Xmax_length3289 _09157_ VGND VGND VPWR VPWR net3289 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire6868 net6869 VGND VGND VPWR VPWR net6868 sky130_fd_sc_hd__buf_1
X_23267_ _03026_ _03033_ VGND VGND VPWR VPWR _03137_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20479_ net3854 net3853 net3852 net3851 net3335 net4060 VGND VGND VPWR VPWR _12268_
+ sky130_fd_sc_hd__mux4_1
X_13020_ net1948 VGND VGND VPWR VPWR _05293_ sky130_fd_sc_hd__clkbuf_1
X_25006_ _04760_ _04761_ VGND VGND VPWR VPWR _04762_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22218_ _02128_ _02133_ _02222_ VGND VGND VPWR VPWR _02223_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_144_Left_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23198_ _03064_ _03066_ VGND VGND VPWR VPWR _03068_ sky130_fd_sc_hd__nand2_1
X_22149_ net1708 VGND VGND VPWR VPWR _02155_ sky130_fd_sc_hd__inv_2
X_14971_ net2834 net3555 net3553 net3545 VGND VGND VPWR VPWR _07045_ sky130_fd_sc_hd__o22a_1
Xwire1120 _06405_ VGND VGND VPWR VPWR net1120 sky130_fd_sc_hd__buf_1
Xwire1131 _05583_ VGND VGND VPWR VPWR net1131 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_22_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16710_ _08736_ _08737_ VGND VGND VPWR VPWR _08738_ sky130_fd_sc_hd__xnor2_1
X_13922_ _06186_ _06187_ VGND VGND VPWR VPWR _06188_ sky130_fd_sc_hd__xnor2_1
Xwire1142 _05193_ VGND VGND VPWR VPWR net1142 sky130_fd_sc_hd__clkbuf_1
X_25908_ clknet_leaf_33_clk _00781_ net8691 VGND VGND VPWR VPWR pid_q.out\[4\] sky130_fd_sc_hd__dfrtp_1
X_17690_ _09537_ _09569_ _09524_ _09523_ _09522_ VGND VGND VPWR VPWR _09570_ sky130_fd_sc_hd__a2111o_1
Xwire1153 _05026_ VGND VGND VPWR VPWR net1153 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1164 _03615_ VGND VGND VPWR VPWR net1164 sky130_fd_sc_hd__buf_1
Xwire1175 net1176 VGND VGND VPWR VPWR net1175 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1186 _00929_ VGND VGND VPWR VPWR net1186 sky130_fd_sc_hd__buf_1
X_16641_ _08678_ VGND VGND VPWR VPWR _00251_ sky130_fd_sc_hd__clkbuf_1
X_13853_ _06115_ _06119_ VGND VGND VPWR VPWR _06120_ sky130_fd_sc_hd__xnor2_1
X_25839_ clknet_leaf_31_clk _00712_ net8684 VGND VGND VPWR VPWR pid_q.curr_error\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1197 net1198 VGND VGND VPWR VPWR net1197 sky130_fd_sc_hd__buf_1
XFILLER_0_53_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12804_ _04955_ _04941_ _05075_ VGND VGND VPWR VPWR _05077_ sky130_fd_sc_hd__nor3_1
X_19360_ _11156_ _11160_ VGND VGND VPWR VPWR _11197_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_153_Left_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16572_ _08626_ _08627_ _08630_ VGND VGND VPWR VPWR _08631_ sky130_fd_sc_hd__or3_1
X_13784_ net7665 net1312 VGND VGND VPWR VPWR _06052_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18311_ net7046 _09675_ _10108_ VGND VGND VPWR VPWR _10162_ sky130_fd_sc_hd__nor3_1
X_15523_ _07594_ _07595_ VGND VGND VPWR VPWR _07596_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12735_ _05005_ _05006_ _05007_ VGND VGND VPWR VPWR _05008_ sky130_fd_sc_hd__o21a_1
X_19291_ net2515 net3213 _10941_ net6291 VGND VGND VPWR VPWR _11128_ sky130_fd_sc_hd__o211ai_1
X_18242_ _10090_ net1777 VGND VGND VPWR VPWR _10093_ sky130_fd_sc_hd__nand2_1
X_12666_ _04936_ _04937_ _04938_ VGND VGND VPWR VPWR _04939_ sky130_fd_sc_hd__a21oi_2
X_15454_ net4175 net4173 VGND VGND VPWR VPWR _07528_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout7942 svm0.periodTop\[0\] VGND VGND VPWR VPWR net7942 sky130_fd_sc_hd__clkbuf_1
Xfanout8687 net8695 VGND VGND VPWR VPWR net8687 sky130_fd_sc_hd__buf_1
XFILLER_0_143_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14405_ _06607_ VGND VGND VPWR VPWR _00086_ sky130_fd_sc_hd__clkbuf_1
X_18173_ _09688_ _09780_ _09781_ VGND VGND VPWR VPWR _10024_ sky130_fd_sc_hd__o21ai_1
Xwire8771 net8772 VGND VGND VPWR VPWR net8771 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_25_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15385_ _07140_ net2251 net2740 VGND VGND VPWR VPWR _07459_ sky130_fd_sc_hd__and3_1
X_12597_ _04877_ VGND VGND VPWR VPWR _00001_ sky130_fd_sc_hd__inv_2
Xwire8782 net8781 VGND VGND VPWR VPWR net8782 sky130_fd_sc_hd__buf_1
XFILLER_0_154_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8793 net8794 VGND VGND VPWR VPWR net8793 sky130_fd_sc_hd__clkbuf_1
X_17124_ net6936 net1819 _09078_ VGND VGND VPWR VPWR _09080_ sky130_fd_sc_hd__or3_1
Xwire450 _06021_ VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14336_ net8243 net3642 VGND VGND VPWR VPWR _06554_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire472 net473 VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire483 net484 VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__clkbuf_1
Xwire494 net495 VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__clkbuf_1
X_14267_ net60 _06511_ _06515_ net9014 VGND VGND VPWR VPWR _00040_ sky130_fd_sc_hd__a22o_1
X_17055_ net2171 _09013_ VGND VGND VPWR VPWR _09014_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_64_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13218_ net1946 _05490_ VGND VGND VPWR VPWR _05491_ sky130_fd_sc_hd__xor2_2
XFILLER_0_122_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16006_ _08066_ _08073_ VGND VGND VPWR VPWR _08074_ sky130_fd_sc_hd__xnor2_1
X_14198_ _06401_ _06419_ _06457_ VGND VGND VPWR VPWR _06458_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13149_ net7909 net2956 net4254 VGND VGND VPWR VPWR _05422_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17957_ net7082 net7108 VGND VGND VPWR VPWR _09808_ sky130_fd_sc_hd__nand2_1
X_16908_ net6373 _08871_ VGND VGND VPWR VPWR _08872_ sky130_fd_sc_hd__nor2_1
X_17888_ _09092_ net3242 _09738_ VGND VGND VPWR VPWR _09739_ sky130_fd_sc_hd__or3_1
XFILLER_0_164_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19627_ net3186 _10923_ _11401_ _11461_ _11463_ VGND VGND VPWR VPWR _11464_ sky130_fd_sc_hd__o311a_1
XFILLER_0_73_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16839_ _08810_ VGND VGND VPWR VPWR _00317_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19558_ net6274 _11392_ _11394_ VGND VGND VPWR VPWR _11395_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_180_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18509_ net3229 _10304_ _10357_ VGND VGND VPWR VPWR _10358_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_119_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19489_ net3190 _11325_ VGND VGND VPWR VPWR _11326_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21520_ _01521_ net478 VGND VGND VPWR VPWR _01533_ sky130_fd_sc_hd__xor2_1
XFILLER_0_180_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21451_ _01348_ _01355_ _01463_ _01351_ VGND VGND VPWR VPWR _01464_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20402_ net811 _12199_ VGND VGND VPWR VPWR _12200_ sky130_fd_sc_hd__xor2_1
X_24170_ pid_q.prev_error\[8\] pid_q.curr_error\[8\] VGND VGND VPWR VPWR _04032_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21382_ net1182 _01395_ VGND VGND VPWR VPWR _01396_ sky130_fd_sc_hd__xnor2_2
Xwire5408 net5406 VGND VGND VPWR VPWR net5408 sky130_fd_sc_hd__buf_1
XFILLER_0_160_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5419 net5420 VGND VGND VPWR VPWR net5419 sky130_fd_sc_hd__clkbuf_1
X_23121_ net5062 net4683 VGND VGND VPWR VPWR _02991_ sky130_fd_sc_hd__nand2_1
X_20333_ net6515 net2586 net949 VGND VGND VPWR VPWR _12136_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_141_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4707 net4701 VGND VGND VPWR VPWR net4707 sky130_fd_sc_hd__buf_1
XFILLER_0_189_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4718 net4715 VGND VGND VPWR VPWR net4718 sky130_fd_sc_hd__buf_1
Xwire4729 net4730 VGND VGND VPWR VPWR net4729 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23052_ net4865 net4742 VGND VGND VPWR VPWR _02922_ sky130_fd_sc_hd__xor2_1
XFILLER_0_113_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20264_ _12075_ VGND VGND VPWR VPWR _00478_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22003_ pid_d.prev_error\[8\] pid_d.curr_error\[8\] VGND VGND VPWR VPWR _02011_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20195_ _11984_ _11981_ _12018_ _12019_ VGND VGND VPWR VPWR _12020_ sky130_fd_sc_hd__a31o_1
Xinput106 pid_d_data[3] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_1
Xinput117 pid_q_addr[12] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_1
Xinput128 pid_q_addr[8] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_1
Xinput139 pid_q_data[3] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_1
X_23954_ net5020 net4499 VGND VGND VPWR VPWR _03818_ sky130_fd_sc_hd__nand2_1
X_22905_ pid_d.curr_int\[10\] _02797_ VGND VGND VPWR VPWR _02798_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23885_ _03641_ _03650_ _03749_ VGND VGND VPWR VPWR _03750_ sky130_fd_sc_hd__a21o_1
X_25624_ clknet_leaf_117_clk _00497_ net8331 VGND VGND VPWR VPWR cordic0.slte0.opA\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_22836_ _02733_ _02727_ _02728_ _02735_ VGND VGND VPWR VPWR _02736_ sky130_fd_sc_hd__a31o_1
XFILLER_0_149_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22767_ _02689_ VGND VGND VPWR VPWR _00612_ sky130_fd_sc_hd__clkbuf_1
X_25555_ clknet_leaf_72_clk net6632 net8468 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8012 net8013 VGND VGND VPWR VPWR net8012 sky130_fd_sc_hd__clkbuf_2
X_24506_ _04361_ _04362_ VGND VGND VPWR VPWR _04363_ sky130_fd_sc_hd__xor2_1
X_21718_ _01728_ _01638_ pid_d.prev_error\[4\] VGND VGND VPWR VPWR _01729_ sky130_fd_sc_hd__o21ba_1
X_25486_ clknet_leaf_46_clk _00366_ net8780 VGND VGND VPWR VPWR svm0.tA\[8\] sky130_fd_sc_hd__dfrtp_1
Xwire8023 net8024 VGND VGND VPWR VPWR net8023 sky130_fd_sc_hd__buf_1
X_22698_ _02640_ VGND VGND VPWR VPWR _00592_ sky130_fd_sc_hd__clkbuf_1
Xwire8034 net8035 VGND VGND VPWR VPWR net8034 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_117_Right_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout7249 net7262 VGND VGND VPWR VPWR net7249 sky130_fd_sc_hd__clkbuf_1
Xwire8045 net8041 VGND VGND VPWR VPWR net8045 sky130_fd_sc_hd__buf_1
Xwire7300 net7301 VGND VGND VPWR VPWR net7300 sky130_fd_sc_hd__clkbuf_1
Xfanout6515 net6517 VGND VGND VPWR VPWR net6515 sky130_fd_sc_hd__clkbuf_2
Xwire8056 net8057 VGND VGND VPWR VPWR net8056 sky130_fd_sc_hd__buf_1
Xwire7311 net7312 VGND VGND VPWR VPWR net7311 sky130_fd_sc_hd__clkbuf_1
X_24437_ net4493 _04294_ VGND VGND VPWR VPWR _04295_ sky130_fd_sc_hd__nand2_1
X_21649_ _01557_ _01559_ _01659_ VGND VGND VPWR VPWR _01660_ sky130_fd_sc_hd__a21oi_2
Xwire8067 net8068 VGND VGND VPWR VPWR net8067 sky130_fd_sc_hd__clkbuf_1
Xwire7322 net7323 VGND VGND VPWR VPWR net7322 sky130_fd_sc_hd__clkbuf_1
Xwire8078 net8079 VGND VGND VPWR VPWR net8078 sky130_fd_sc_hd__clkbuf_1
Xwire7333 net7334 VGND VGND VPWR VPWR net7333 sky130_fd_sc_hd__clkbuf_1
Xwire7344 net7345 VGND VGND VPWR VPWR net7344 sky130_fd_sc_hd__clkbuf_1
Xwire8089 net8090 VGND VGND VPWR VPWR net8089 sky130_fd_sc_hd__clkbuf_1
Xwire6610 net6612 VGND VGND VPWR VPWR net6610 sky130_fd_sc_hd__buf_1
XFILLER_0_90_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15170_ _07191_ _07243_ VGND VGND VPWR VPWR _07244_ sky130_fd_sc_hd__xnor2_1
X_24368_ _04221_ _04226_ VGND VGND VPWR VPWR _04227_ sky130_fd_sc_hd__xnor2_2
Xwire7366 net7367 VGND VGND VPWR VPWR net7366 sky130_fd_sc_hd__clkbuf_1
Xwire6621 net6618 VGND VGND VPWR VPWR net6621 sky130_fd_sc_hd__buf_1
Xwire6643 net6644 VGND VGND VPWR VPWR net6643 sky130_fd_sc_hd__buf_1
Xwire6654 net6655 VGND VGND VPWR VPWR net6654 sky130_fd_sc_hd__clkbuf_1
X_14121_ net1560 net1124 net7603 VGND VGND VPWR VPWR _06383_ sky130_fd_sc_hd__and3b_1
Xmax_length3086 _02599_ VGND VGND VPWR VPWR net3086 sky130_fd_sc_hd__buf_1
Xwire7399 net7400 VGND VGND VPWR VPWR net7399 sky130_fd_sc_hd__clkbuf_1
X_23319_ _03187_ _03188_ VGND VGND VPWR VPWR _03189_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5920 net5921 VGND VGND VPWR VPWR net5920 sky130_fd_sc_hd__buf_1
Xwire6665 net6666 VGND VGND VPWR VPWR net6665 sky130_fd_sc_hd__clkbuf_1
Xmax_length2363 net2364 VGND VGND VPWR VPWR net2363 sky130_fd_sc_hd__clkbuf_1
X_24299_ _04157_ _04158_ VGND VGND VPWR VPWR _04159_ sky130_fd_sc_hd__xnor2_1
Xwire6687 net6686 VGND VGND VPWR VPWR net6687 sky130_fd_sc_hd__buf_1
Xwire5942 net5945 VGND VGND VPWR VPWR net5942 sky130_fd_sc_hd__clkbuf_1
Xwire6698 net6699 VGND VGND VPWR VPWR net6698 sky130_fd_sc_hd__buf_1
XFILLER_0_104_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14052_ _06315_ VGND VGND VPWR VPWR _06316_ sky130_fd_sc_hd__inv_2
Xwire5964 pid_d.curr_error\[15\] VGND VGND VPWR VPWR net5964 sky130_fd_sc_hd__buf_1
Xwire5975 pid_d.curr_int\[12\] VGND VGND VPWR VPWR net5975 sky130_fd_sc_hd__buf_1
Xwire5986 pid_d.curr_int\[0\] VGND VGND VPWR VPWR net5986 sky130_fd_sc_hd__buf_1
X_13003_ _05274_ _05275_ VGND VGND VPWR VPWR _05276_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5997 net5998 VGND VGND VPWR VPWR net5997 sky130_fd_sc_hd__buf_1
X_18860_ _10686_ _10688_ _10701_ net3221 VGND VGND VPWR VPWR _10702_ sky130_fd_sc_hd__o2bb2a_1
X_17811_ net3988 _09661_ VGND VGND VPWR VPWR _09662_ sky130_fd_sc_hd__or2_1
X_18791_ net6855 _10584_ _10633_ _10634_ VGND VGND VPWR VPWR _10635_ sky130_fd_sc_hd__a31o_1
X_17742_ net4235 net6454 _06646_ _09595_ VGND VGND VPWR VPWR _00436_ sky130_fd_sc_hd__a31o_1
X_14954_ _07027_ VGND VGND VPWR VPWR _07028_ sky130_fd_sc_hd__buf_1
X_13905_ _06169_ _06170_ VGND VGND VPWR VPWR _06171_ sky130_fd_sc_hd__xor2_1
X_17673_ _09550_ _09546_ net4002 svm0.tA\[2\] VGND VGND VPWR VPWR _09553_ sky130_fd_sc_hd__o2bb2a_1
X_14885_ _06960_ VGND VGND VPWR VPWR _00213_ sky130_fd_sc_hd__clkbuf_1
X_19412_ _11248_ _11107_ _11096_ VGND VGND VPWR VPWR _11249_ sky130_fd_sc_hd__mux2_1
X_16624_ matmul0.alpha_pass\[1\] net3383 net6551 VGND VGND VPWR VPWR _08664_ sky130_fd_sc_hd__mux2_1
X_13836_ _06099_ _06102_ VGND VGND VPWR VPWR _06103_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19343_ _11174_ _11176_ _11178_ _11179_ VGND VGND VPWR VPWR _11180_ sky130_fd_sc_hd__a211o_1
X_16555_ net3420 net2622 net2219 net1841 VGND VGND VPWR VPWR _08614_ sky130_fd_sc_hd__or4_1
X_13767_ net7721 net1307 VGND VGND VPWR VPWR _06035_ sky130_fd_sc_hd__nand2_1
X_15506_ net3573 net3569 net4098 net4096 VGND VGND VPWR VPWR _07579_ sky130_fd_sc_hd__o22a_1
X_12718_ _04942_ _04943_ VGND VGND VPWR VPWR _04991_ sky130_fd_sc_hd__xnor2_1
X_19274_ _11109_ _11110_ VGND VGND VPWR VPWR _11111_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16486_ _08546_ VGND VGND VPWR VPWR _00228_ sky130_fd_sc_hd__clkbuf_1
X_13698_ _05965_ _05966_ VGND VGND VPWR VPWR _05967_ sky130_fd_sc_hd__nor2_1
Xfanout8462 net8483 VGND VGND VPWR VPWR net8462 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_127_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18225_ _09696_ _09604_ _10038_ VGND VGND VPWR VPWR _10076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15437_ net4092 net4089 VGND VGND VPWR VPWR _07511_ sky130_fd_sc_hd__or2_1
Xfanout8495 net8504 VGND VGND VPWR VPWR net8495 sky130_fd_sc_hd__buf_1
X_12649_ net7813 net1346 VGND VGND VPWR VPWR _04922_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18156_ _09960_ _09969_ _09968_ VGND VGND VPWR VPWR _10007_ sky130_fd_sc_hd__a21o_1
X_15368_ _07420_ _07421_ VGND VGND VPWR VPWR _07442_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17107_ _09060_ _09062_ VGND VGND VPWR VPWR _09064_ sky130_fd_sc_hd__and2_1
X_14319_ net4235 net6443 net3638 _06536_ _06540_ VGND VGND VPWR VPWR _06541_ sky130_fd_sc_hd__a311o_2
Xwire280 _08432_ VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__clkbuf_1
Xwire291 net292 VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__clkbuf_1
X_18087_ _09935_ _09937_ _08914_ VGND VGND VPWR VPWR _09938_ sky130_fd_sc_hd__mux2_2
XFILLER_0_180_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15299_ net3596 net3590 net4198 net4197 VGND VGND VPWR VPWR _07373_ sky130_fd_sc_hd__o22a_1
XFILLER_0_151_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17038_ net7053 _08997_ net1804 VGND VGND VPWR VPWR _08998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18989_ _10821_ net3899 _10825_ net6339 net6262 VGND VGND VPWR VPWR _10826_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_139_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20951_ _00944_ _00963_ _00966_ VGND VGND VPWR VPWR _00967_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23670_ _03525_ _03536_ VGND VGND VPWR VPWR _03537_ sky130_fd_sc_hd__nor2_1
XFILLER_0_191_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20882_ net5491 net5935 VGND VGND VPWR VPWR _00898_ sky130_fd_sc_hd__and2_1
XFILLER_0_191_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6629 net6630 VGND VGND VPWR VPWR net6629 sky130_fd_sc_hd__buf_1
X_22621_ net3089 _02590_ _02591_ VGND VGND VPWR VPWR _02592_ sky130_fd_sc_hd__and3_1
XFILLER_0_177_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length5939 net5940 VGND VGND VPWR VPWR net5939 sky130_fd_sc_hd__clkbuf_1
X_25340_ clknet_leaf_56_clk _00223_ net8723 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_22552_ net9159 net2049 _02538_ VGND VGND VPWR VPWR _00548_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21503_ net1182 net1181 _01392_ VGND VGND VPWR VPWR _01516_ sky130_fd_sc_hd__o21ba_1
X_25271_ clknet_leaf_88_clk _00154_ net8438 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.c\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_22483_ net5671 net5647 VGND VGND VPWR VPWR _02484_ sky130_fd_sc_hd__and2b_1
XFILLER_0_63_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24222_ _03964_ _03966_ _04082_ VGND VGND VPWR VPWR _04083_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_118_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21434_ _01444_ _01445_ _01446_ VGND VGND VPWR VPWR _01447_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5205 net5207 VGND VGND VPWR VPWR net5205 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24153_ _04005_ _04014_ VGND VGND VPWR VPWR _04015_ sky130_fd_sc_hd__xnor2_1
Xwire5216 net5217 VGND VGND VPWR VPWR net5216 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21365_ _01257_ _01258_ _01378_ VGND VGND VPWR VPWR _01379_ sky130_fd_sc_hd__a21bo_1
Xwire5238 net5239 VGND VGND VPWR VPWR net5238 sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_110_clk clknet_4_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_110_clk
+ sky130_fd_sc_hd__clkbuf_16
Xwire4504 net4503 VGND VGND VPWR VPWR net4504 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire5249 net5243 VGND VGND VPWR VPWR net5249 sky130_fd_sc_hd__clkbuf_1
X_23104_ net4968 net4755 VGND VGND VPWR VPWR _02974_ sky130_fd_sc_hd__nand2_1
X_20316_ net1223 _12119_ VGND VGND VPWR VPWR _12120_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4526 net4527 VGND VGND VPWR VPWR net4526 sky130_fd_sc_hd__clkbuf_1
X_24084_ _03946_ _03854_ pid_q.prev_error\[6\] VGND VGND VPWR VPWR _03947_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_102_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4537 net4539 VGND VGND VPWR VPWR net4537 sky130_fd_sc_hd__buf_1
X_21296_ net5889 _01310_ VGND VGND VPWR VPWR _01311_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3803 net3804 VGND VGND VPWR VPWR net3803 sky130_fd_sc_hd__clkbuf_1
Xwire4559 net4560 VGND VGND VPWR VPWR net4559 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3814 net3815 VGND VGND VPWR VPWR net3814 sky130_fd_sc_hd__clkbuf_1
X_23035_ _02899_ _02904_ VGND VGND VPWR VPWR _02905_ sky130_fd_sc_hd__nand2_1
Xwire3825 net3826 VGND VGND VPWR VPWR net3825 sky130_fd_sc_hd__clkbuf_1
X_20247_ net8121 _12061_ VGND VGND VPWR VPWR _12062_ sky130_fd_sc_hd__nor2_1
Xwire3836 net3837 VGND VGND VPWR VPWR net3836 sky130_fd_sc_hd__clkbuf_2
Xwire3847 _12276_ VGND VGND VPWR VPWR net3847 sky130_fd_sc_hd__buf_1
Xwire3869 _11271_ VGND VGND VPWR VPWR net3869 sky130_fd_sc_hd__buf_1
X_20178_ _12000_ _12003_ _11410_ VGND VGND VPWR VPWR _12004_ sky130_fd_sc_hd__o21a_1
XFILLER_0_157_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24986_ pid_q.kp\[12\] _04726_ net1634 VGND VGND VPWR VPWR _04748_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23937_ _03797_ _03799_ VGND VGND VPWR VPWR _03801_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length8565 net8566 VGND VGND VPWR VPWR net8565 sky130_fd_sc_hd__buf_1
Xmax_length7831 net7832 VGND VGND VPWR VPWR net7831 sky130_fd_sc_hd__buf_1
XFILLER_0_169_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14670_ net7160 _06821_ VGND VGND VPWR VPWR _06822_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_168_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23868_ _03731_ _03732_ VGND VGND VPWR VPWR _03733_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13621_ _05791_ _05796_ _05789_ VGND VGND VPWR VPWR _05891_ sky130_fd_sc_hd__a21o_1
X_25607_ clknet_leaf_109_clk _00480_ net8344 VGND VGND VPWR VPWR cordic0.slte0.opB\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22819_ _02721_ VGND VGND VPWR VPWR _00632_ sky130_fd_sc_hd__clkbuf_1
X_23799_ pid_q.prev_error\[4\] pid_q.curr_error\[4\] VGND VGND VPWR VPWR _03665_ sky130_fd_sc_hd__xnor2_1
Xmax_length7897 net7898 VGND VGND VPWR VPWR net7897 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16340_ _08325_ net1249 _08323_ VGND VGND VPWR VPWR _08403_ sky130_fd_sc_hd__o21ba_1
X_13552_ net1573 net1347 net7617 VGND VGND VPWR VPWR _05823_ sky130_fd_sc_hd__and3b_1
X_25538_ clknet_leaf_33_clk _00418_ net8687 VGND VGND VPWR VPWR pid_q.prev_int\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6301 net6307 VGND VGND VPWR VPWR net6301 sky130_fd_sc_hd__buf_1
X_13483_ _05754_ _05755_ VGND VGND VPWR VPWR _05756_ sky130_fd_sc_hd__nand2_1
X_16271_ _08264_ _08261_ _08334_ VGND VGND VPWR VPWR _08335_ sky130_fd_sc_hd__a21o_1
X_25469_ clknet_leaf_52_clk _00349_ net8806 VGND VGND VPWR VPWR svm0.tB\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_192_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18010_ net7051 net7006 VGND VGND VPWR VPWR _09861_ sky130_fd_sc_hd__or2b_1
Xfanout5600 pid_d.mult0.a\[3\] VGND VGND VPWR VPWR net5600 sky130_fd_sc_hd__clkbuf_1
X_15222_ net1882 net1544 VGND VGND VPWR VPWR _07296_ sky130_fd_sc_hd__xnor2_1
Xwire7141 net7142 VGND VGND VPWR VPWR net7141 sky130_fd_sc_hd__buf_1
XFILLER_0_125_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5611 net5616 VGND VGND VPWR VPWR net5611 sky130_fd_sc_hd__buf_1
Xwire7152 matmul0.sin\[7\] VGND VGND VPWR VPWR net7152 sky130_fd_sc_hd__clkbuf_2
Xwire7163 net7164 VGND VGND VPWR VPWR net7163 sky130_fd_sc_hd__buf_1
Xwire7174 matmul0.cos\[8\] VGND VGND VPWR VPWR net7174 sky130_fd_sc_hd__clkbuf_1
Xwire6440 net6441 VGND VGND VPWR VPWR net6440 sky130_fd_sc_hd__clkbuf_1
Xwire7185 matmul0.b\[7\] VGND VGND VPWR VPWR net7185 sky130_fd_sc_hd__clkbuf_1
Xwire6451 net6450 VGND VGND VPWR VPWR net6451 sky130_fd_sc_hd__clkbuf_2
Xwire7196 net7197 VGND VGND VPWR VPWR net7196 sky130_fd_sc_hd__clkbuf_1
X_15153_ net3583 net3581 net3511 net3506 VGND VGND VPWR VPWR _07227_ sky130_fd_sc_hd__o22a_1
Xwire6473 net6469 VGND VGND VPWR VPWR net6473 sky130_fd_sc_hd__buf_1
Xwire6484 net6485 VGND VGND VPWR VPWR net6484 sky130_fd_sc_hd__buf_1
X_14104_ net217 net403 VGND VGND VPWR VPWR _06366_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5750 net5744 VGND VGND VPWR VPWR net5750 sky130_fd_sc_hd__buf_1
X_19961_ net3153 _11755_ VGND VGND VPWR VPWR _11792_ sky130_fd_sc_hd__or2_1
X_15084_ net3559 _07157_ VGND VGND VPWR VPWR _07158_ sky130_fd_sc_hd__nor2_1
Xfanout4965 net4977 VGND VGND VPWR VPWR net4965 sky130_fd_sc_hd__clkbuf_1
Xwire5761 net5758 VGND VGND VPWR VPWR net5761 sky130_fd_sc_hd__buf_1
Xwire5772 net5773 VGND VGND VPWR VPWR net5772 sky130_fd_sc_hd__clkbuf_1
Xmax_length1470 net1471 VGND VGND VPWR VPWR net1470 sky130_fd_sc_hd__buf_1
X_14035_ net7680 net1323 VGND VGND VPWR VPWR _06299_ sky130_fd_sc_hd__nand2_1
X_18912_ _10278_ _10531_ _10751_ net6828 net6864 VGND VGND VPWR VPWR _10752_ sky130_fd_sc_hd__a221oi_1
Xwire5794 net5792 VGND VGND VPWR VPWR net5794 sky130_fd_sc_hd__buf_1
X_19892_ _11667_ _11720_ _11724_ VGND VGND VPWR VPWR _11725_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_38_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18843_ _10666_ _10685_ VGND VGND VPWR VPWR _10686_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18774_ net764 _10600_ VGND VGND VPWR VPWR _10618_ sky130_fd_sc_hd__or2_1
X_15986_ net2712 net4076 VGND VGND VPWR VPWR _08054_ sky130_fd_sc_hd__nor2_1
X_17725_ net6506 net1831 VGND VGND VPWR VPWR _09585_ sky130_fd_sc_hd__nor2_1
X_14937_ net4161 net4157 VGND VGND VPWR VPWR _07011_ sky130_fd_sc_hd__or2_1
X_17656_ net3279 svm0.tA\[10\] VGND VGND VPWR VPWR _09536_ sky130_fd_sc_hd__or2_1
XFILLER_0_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14868_ matmul0.b\[6\] matmul0.matmul_stage_inst.f\[6\] _06950_ VGND VGND VPWR VPWR
+ _06952_ sky130_fd_sc_hd__mux2_1
X_16607_ _08653_ VGND VGND VPWR VPWR _00242_ sky130_fd_sc_hd__clkbuf_1
X_13819_ net9137 net1126 net256 net1926 VGND VGND VPWR VPWR _00021_ sky130_fd_sc_hd__a22o_1
X_17587_ svm0.tC\[15\] _09422_ _09468_ VGND VGND VPWR VPWR _09469_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_159_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14799_ net8981 net2871 _06916_ VGND VGND VPWR VPWR _00171_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19326_ _10821_ net3210 _11140_ VGND VGND VPWR VPWR _11163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16538_ net1084 _08596_ _08594_ VGND VGND VPWR VPWR _08597_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_85_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19257_ _11070_ _11092_ _11093_ VGND VGND VPWR VPWR _11094_ sky130_fd_sc_hd__o21a_1
XFILLER_0_169_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16469_ _08528_ _08529_ VGND VGND VPWR VPWR _08530_ sky130_fd_sc_hd__nor2b_1
XFILLER_0_183_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18208_ _09798_ _09676_ net6997 VGND VGND VPWR VPWR _10059_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19188_ net6201 net6240 VGND VGND VPWR VPWR _11025_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18139_ _09945_ VGND VGND VPWR VPWR _09990_ sky130_fd_sc_hd__inv_2
Xhold102 pid_q.curr_error\[1\] VGND VGND VPWR VPWR net9055 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 pid_q.curr_int\[13\] VGND VGND VPWR VPWR net9066 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 pid_q.curr_int\[11\] VGND VGND VPWR VPWR net9077 sky130_fd_sc_hd__dlygate4sd3_1
X_21150_ _01148_ _01165_ VGND VGND VPWR VPWR _01166_ sky130_fd_sc_hd__xnor2_1
Xhold135 cordic0.sin\[2\] VGND VGND VPWR VPWR net9088 sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 svm0.tB\[8\] VGND VGND VPWR VPWR net9099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 svm0.in_valid VGND VGND VPWR VPWR net9110 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold168 pid_d.prev_error\[10\] VGND VGND VPWR VPWR net9121 sky130_fd_sc_hd__dlygate4sd3_1
X_20101_ _11928_ _11920_ VGND VGND VPWR VPWR _11929_ sky130_fd_sc_hd__nand2_1
Xhold179 svm0.tB\[5\] VGND VGND VPWR VPWR net9132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21081_ net5556 _01068_ _01094_ _01096_ _01093_ VGND VGND VPWR VPWR _01097_ sky130_fd_sc_hd__a32o_1
Xwire2409 net2410 VGND VGND VPWR VPWR net2409 sky130_fd_sc_hd__buf_1
X_20032_ _11490_ _11861_ VGND VGND VPWR VPWR _11862_ sky130_fd_sc_hd__xor2_1
Xwire1708 net1709 VGND VGND VPWR VPWR net1708 sky130_fd_sc_hd__buf_1
Xwire1719 _01843_ VGND VGND VPWR VPWR net1719 sky130_fd_sc_hd__buf_1
X_24840_ net7482 net629 _04115_ VGND VGND VPWR VPWR _04653_ sky130_fd_sc_hd__a21o_1
X_24771_ _04597_ _04598_ net5220 VGND VGND VPWR VPWR _04599_ sky130_fd_sc_hd__a21oi_1
X_21983_ _01989_ _01990_ VGND VGND VPWR VPWR _01991_ sky130_fd_sc_hd__and2_1
X_23722_ _03518_ _03522_ _03587_ VGND VGND VPWR VPWR _03588_ sky130_fd_sc_hd__a21oi_2
Xmax_length7127 net7128 VGND VGND VPWR VPWR net7127 sky130_fd_sc_hd__clkbuf_1
X_20934_ _00901_ _00902_ VGND VGND VPWR VPWR _00950_ sky130_fd_sc_hd__xor2_1
XFILLER_0_68_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6426 cordic0.sin\[5\] VGND VGND VPWR VPWR net6426 sky130_fd_sc_hd__clkbuf_1
X_23653_ net4495 _03519_ VGND VGND VPWR VPWR _03520_ sky130_fd_sc_hd__nand2_1
X_20865_ net5613 VGND VGND VPWR VPWR _00881_ sky130_fd_sc_hd__inv_2
Xmax_length6448 net6449 VGND VGND VPWR VPWR net6448 sky130_fd_sc_hd__buf_1
Xmax_length6459 net6457 VGND VGND VPWR VPWR net6459 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_76_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22604_ net9013 net2045 net2042 _02578_ VGND VGND VPWR VPWR _00560_ sky130_fd_sc_hd__a22o_1
X_23584_ net1670 net1667 _03363_ VGND VGND VPWR VPWR _03452_ sky130_fd_sc_hd__a21bo_1
X_20796_ net5635 net5730 VGND VGND VPWR VPWR _00812_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25323_ clknet_leaf_74_clk _00206_ net8464 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.f\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_22535_ net5969 net2379 net2047 VGND VGND VPWR VPWR _02530_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22466_ _02464_ _02466_ VGND VGND VPWR VPWR _02467_ sky130_fd_sc_hd__xnor2_1
X_25254_ clknet_leaf_88_clk _00137_ net8430 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.b\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5002 net5003 VGND VGND VPWR VPWR net5002 sky130_fd_sc_hd__clkbuf_1
X_24205_ _04060_ _04065_ VGND VGND VPWR VPWR _04066_ sky130_fd_sc_hd__xnor2_1
X_21417_ pid_d.prev_error\[2\] net5971 VGND VGND VPWR VPWR _01431_ sky130_fd_sc_hd__xor2_1
Xwire5013 net5014 VGND VGND VPWR VPWR net5013 sky130_fd_sc_hd__buf_1
X_25185_ clknet_leaf_69_clk _00074_ net8468 VGND VGND VPWR VPWR matmul0.a_in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire5024 net5025 VGND VGND VPWR VPWR net5024 sky130_fd_sc_hd__buf_1
X_22397_ _02397_ _02398_ VGND VGND VPWR VPWR _02399_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5035 pid_q.mult0.b\[5\] VGND VGND VPWR VPWR net5035 sky130_fd_sc_hd__clkbuf_1
Xwire5046 net5047 VGND VGND VPWR VPWR net5046 sky130_fd_sc_hd__clkbuf_1
X_24136_ _03996_ _03997_ VGND VGND VPWR VPWR _03998_ sky130_fd_sc_hd__nor2_1
Xwire4301 _04872_ VGND VGND VPWR VPWR net4301 sky130_fd_sc_hd__buf_1
Xwire5057 net5058 VGND VGND VPWR VPWR net5057 sky130_fd_sc_hd__buf_1
Xwire4312 _04861_ VGND VGND VPWR VPWR net4312 sky130_fd_sc_hd__clkbuf_1
X_21348_ net5777 net5535 VGND VGND VPWR VPWR _01362_ sky130_fd_sc_hd__nand2_1
Xwire4323 pid_d.state\[5\] VGND VGND VPWR VPWR net4323 sky130_fd_sc_hd__buf_1
Xwire5079 net5080 VGND VGND VPWR VPWR net5079 sky130_fd_sc_hd__buf_1
Xwire3600 net3601 VGND VGND VPWR VPWR net3600 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4345 net4346 VGND VGND VPWR VPWR net4345 sky130_fd_sc_hd__clkbuf_1
X_24067_ net1160 _03929_ VGND VGND VPWR VPWR _03930_ sky130_fd_sc_hd__xnor2_1
Xwire3611 _06928_ VGND VGND VPWR VPWR net3611 sky130_fd_sc_hd__buf_1
Xwire4356 net4357 VGND VGND VPWR VPWR net4356 sky130_fd_sc_hd__buf_1
Xwire4367 net4361 VGND VGND VPWR VPWR net4367 sky130_fd_sc_hd__buf_1
Xwire3622 _06823_ VGND VGND VPWR VPWR net3622 sky130_fd_sc_hd__clkbuf_1
X_21279_ net5731 net5598 VGND VGND VPWR VPWR _01294_ sky130_fd_sc_hd__nand2_1
Xwire4378 pid_d.state\[2\] VGND VGND VPWR VPWR net4378 sky130_fd_sc_hd__clkbuf_1
Xwire3633 net3634 VGND VGND VPWR VPWR net3633 sky130_fd_sc_hd__buf_1
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4389 net4390 VGND VGND VPWR VPWR net4389 sky130_fd_sc_hd__buf_1
XFILLER_0_60_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3644 net3645 VGND VGND VPWR VPWR net3644 sky130_fd_sc_hd__clkbuf_1
X_23018_ _02886_ _02887_ VGND VGND VPWR VPWR _02888_ sky130_fd_sc_hd__nor2_1
Xwire2910 net2911 VGND VGND VPWR VPWR net2910 sky130_fd_sc_hd__clkbuf_1
Xwire3655 net3656 VGND VGND VPWR VPWR net3655 sky130_fd_sc_hd__clkbuf_1
Xwire2921 net2930 VGND VGND VPWR VPWR net2921 sky130_fd_sc_hd__clkbuf_1
Xwire3677 net3678 VGND VGND VPWR VPWR net3677 sky130_fd_sc_hd__buf_1
Xwire2932 net2933 VGND VGND VPWR VPWR net2932 sky130_fd_sc_hd__clkbuf_2
Xwire3688 net3692 VGND VGND VPWR VPWR net3688 sky130_fd_sc_hd__buf_1
Xwire2943 _06501_ VGND VGND VPWR VPWR net2943 sky130_fd_sc_hd__clkbuf_1
Xwire3699 net3700 VGND VGND VPWR VPWR net3699 sky130_fd_sc_hd__buf_1
Xwire2954 net2955 VGND VGND VPWR VPWR net2954 sky130_fd_sc_hd__buf_1
Xwire2965 _05190_ VGND VGND VPWR VPWR net2965 sky130_fd_sc_hd__buf_1
X_15840_ _07802_ _07817_ _07800_ VGND VGND VPWR VPWR _07910_ sky130_fd_sc_hd__a21o_1
Xwire2987 _04909_ VGND VGND VPWR VPWR net2987 sky130_fd_sc_hd__clkbuf_1
Xwire2998 net2999 VGND VGND VPWR VPWR net2998 sky130_fd_sc_hd__clkbuf_1
X_15771_ net2699 net2727 VGND VGND VPWR VPWR _07841_ sky130_fd_sc_hd__nor2_1
X_24969_ _04739_ VGND VGND VPWR VPWR _00764_ sky130_fd_sc_hd__clkbuf_1
X_12983_ net7728 net1616 VGND VGND VPWR VPWR _05256_ sky130_fd_sc_hd__nand2_1
X_17510_ net4067 _09396_ net6659 VGND VGND VPWR VPWR _09397_ sky130_fd_sc_hd__o21a_1
Xmax_length8351 net8352 VGND VGND VPWR VPWR net8351 sky130_fd_sc_hd__buf_1
X_14722_ net8991 _06814_ _06861_ VGND VGND VPWR VPWR _00149_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18490_ _10336_ _10339_ VGND VGND VPWR VPWR _10340_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17441_ net2578 _09336_ VGND VGND VPWR VPWR _09338_ sky130_fd_sc_hd__nor2_1
XFILLER_0_170_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14653_ net7440 net7172 net2874 VGND VGND VPWR VPWR _06811_ sky130_fd_sc_hd__and3_1
XFILLER_0_196_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length7683 net7679 VGND VGND VPWR VPWR net7683 sky130_fd_sc_hd__buf_1
X_13604_ net7770 net1306 VGND VGND VPWR VPWR _05874_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17372_ _09281_ net667 VGND VGND VPWR VPWR _09283_ sky130_fd_sc_hd__and2_1
XFILLER_0_184_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14584_ net3640 _06754_ _06752_ VGND VGND VPWR VPWR _06759_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19111_ _10849_ _10850_ net6182 VGND VGND VPWR VPWR _10948_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16323_ net2629 _08385_ VGND VGND VPWR VPWR _08386_ sky130_fd_sc_hd__nor2_1
X_13535_ _05798_ _05805_ VGND VGND VPWR VPWR _05806_ sky130_fd_sc_hd__xnor2_2
X_19042_ net6252 VGND VGND VPWR VPWR _10879_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16254_ _08311_ _08317_ VGND VGND VPWR VPWR _08318_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_168_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13466_ _05592_ _05593_ _05738_ VGND VGND VPWR VPWR _05739_ sky130_fd_sc_hd__a21o_1
Xfanout6153 net6158 VGND VGND VPWR VPWR net6153 sky130_fd_sc_hd__buf_1
XFILLER_0_3_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6164 cordic0.vec\[0\]\[9\] VGND VGND VPWR VPWR net6164 sky130_fd_sc_hd__buf_1
XFILLER_0_180_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5430 net5439 VGND VGND VPWR VPWR net5430 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout6175 net6192 VGND VGND VPWR VPWR net6175 sky130_fd_sc_hd__buf_1
X_15205_ _07237_ _07239_ VGND VGND VPWR VPWR _07279_ sky130_fd_sc_hd__xor2_1
XFILLER_0_129_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16185_ net2692 net2651 net2214 net2222 net3409 VGND VGND VPWR VPWR _08250_ sky130_fd_sc_hd__o32a_1
X_13397_ net583 _05663_ net581 VGND VGND VPWR VPWR _05670_ sky130_fd_sc_hd__or3b_1
XFILLER_0_50_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15136_ net1894 _07181_ _07176_ VGND VGND VPWR VPWR _07210_ sky130_fd_sc_hd__o21ba_1
Xfanout5496 pid_d.mult0.a\[9\] VGND VGND VPWR VPWR net5496 sky130_fd_sc_hd__clkbuf_1
Xfanout4773 net4780 VGND VGND VPWR VPWR net4773 sky130_fd_sc_hd__buf_1
XFILLER_0_26_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5591 net5592 VGND VGND VPWR VPWR net5591 sky130_fd_sc_hd__clkbuf_1
X_19944_ _11698_ _11703_ _11775_ VGND VGND VPWR VPWR _11776_ sky130_fd_sc_hd__o21a_1
X_15067_ net4111 net4108 VGND VGND VPWR VPWR _07141_ sky130_fd_sc_hd__nor2_1
X_14018_ _06248_ _06256_ _06281_ VGND VGND VPWR VPWR _06282_ sky130_fd_sc_hd__o21a_1
Xwire4890 net4885 VGND VGND VPWR VPWR net4890 sky130_fd_sc_hd__buf_1
X_19875_ _11705_ _11707_ VGND VGND VPWR VPWR _11708_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18826_ net6826 net3920 VGND VGND VPWR VPWR _10669_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18757_ _10558_ _10600_ _10569_ VGND VGND VPWR VPWR _10602_ sky130_fd_sc_hd__or3_1
X_15969_ _08032_ _08036_ VGND VGND VPWR VPWR _08037_ sky130_fd_sc_hd__xnor2_1
X_17708_ net1788 VGND VGND VPWR VPWR _09584_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18688_ net6955 net6867 VGND VGND VPWR VPWR _10534_ sky130_fd_sc_hd__xor2_2
XFILLER_0_172_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17639_ svm0.calc_ready net2568 net876 net8962 net3384 VGND VGND VPWR VPWR _00408_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_72_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20650_ net6484 _12426_ _12427_ VGND VGND VPWR VPWR _12428_ sky130_fd_sc_hd__a21o_1
XFILLER_0_175_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length4309 _04866_ VGND VGND VPWR VPWR net4309 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19309_ net6224 net6290 net6334 VGND VGND VPWR VPWR _11146_ sky130_fd_sc_hd__and3_1
XFILLER_0_162_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20581_ _12295_ _12297_ net2602 VGND VGND VPWR VPWR _12364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length3608 net3609 VGND VGND VPWR VPWR net3608 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_27_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22320_ _02279_ net552 VGND VGND VPWR VPWR _02324_ sky130_fd_sc_hd__or2_1
XFILLER_0_143_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22251_ _02254_ _02176_ _02255_ VGND VGND VPWR VPWR _02256_ sky130_fd_sc_hd__a21o_1
XFILLER_0_103_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21202_ _01029_ _01217_ VGND VGND VPWR VPWR _01218_ sky130_fd_sc_hd__xnor2_1
X_22182_ _02185_ _02186_ VGND VGND VPWR VPWR _02187_ sky130_fd_sc_hd__xnor2_1
X_21133_ net5614 net5908 VGND VGND VPWR VPWR _01149_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2206 net2207 VGND VGND VPWR VPWR net2206 sky130_fd_sc_hd__buf_1
X_21064_ net5552 net5949 VGND VGND VPWR VPWR _01080_ sky130_fd_sc_hd__nand2_1
Xwire2217 net2219 VGND VGND VPWR VPWR net2217 sky130_fd_sc_hd__buf_1
X_25941_ clknet_leaf_120_clk net2379 net8419 VGND VGND VPWR VPWR pid_d.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire2228 _07570_ VGND VGND VPWR VPWR net2228 sky130_fd_sc_hd__buf_1
Xwire2239 net2240 VGND VGND VPWR VPWR net2239 sky130_fd_sc_hd__clkbuf_2
Xwire1505 net1506 VGND VGND VPWR VPWR net1505 sky130_fd_sc_hd__buf_1
X_20015_ _11814_ _11815_ VGND VGND VPWR VPWR _11845_ sky130_fd_sc_hd__nor2_1
Xwire1516 _08101_ VGND VGND VPWR VPWR net1516 sky130_fd_sc_hd__buf_1
X_25872_ clknet_leaf_17_clk _00745_ net8626 VGND VGND VPWR VPWR pid_q.ki\[0\] sky130_fd_sc_hd__dfrtp_1
Xwire1527 net1528 VGND VGND VPWR VPWR net1527 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1538 _07531_ VGND VGND VPWR VPWR net1538 sky130_fd_sc_hd__buf_1
X_24823_ net5156 _04642_ net2000 _04644_ VGND VGND VPWR VPWR _00713_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24754_ _04582_ _04584_ VGND VGND VPWR VPWR _04585_ sky130_fd_sc_hd__xnor2_1
X_21966_ net1047 net1171 VGND VGND VPWR VPWR _01974_ sky130_fd_sc_hd__and2_1
X_23705_ pid_q.prev_error\[3\] pid_q.curr_error\[3\] VGND VGND VPWR VPWR _03572_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_178_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20917_ _00921_ _00924_ _00932_ VGND VGND VPWR VPWR _00933_ sky130_fd_sc_hd__a21o_1
X_24685_ pid_q.curr_error\[14\] net3021 _04509_ VGND VGND VPWR VPWR _04525_ sky130_fd_sc_hd__and3_1
X_21897_ net599 _01905_ VGND VGND VPWR VPWR _01906_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6256 net6257 VGND VGND VPWR VPWR net6256 sky130_fd_sc_hd__clkbuf_1
X_23636_ _03493_ _03502_ VGND VGND VPWR VPWR _03503_ sky130_fd_sc_hd__xnor2_2
X_20848_ _12514_ _12515_ _00863_ VGND VGND VPWR VPWR _00864_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_154_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23567_ net4702 net4876 VGND VGND VPWR VPWR _03435_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20779_ net5597 net5761 VGND VGND VPWR VPWR _12550_ sky130_fd_sc_hd__nand2_1
XFILLER_0_193_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length4843 net4844 VGND VGND VPWR VPWR net4843 sky130_fd_sc_hd__buf_1
Xwire802 _02074_ VGND VGND VPWR VPWR net802 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_119_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire813 _11238_ VGND VGND VPWR VPWR net813 sky130_fd_sc_hd__clkbuf_1
X_13320_ net7747 net2330 net2325 VGND VGND VPWR VPWR _05593_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25306_ clknet_leaf_71_clk _00189_ net8461 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.e\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire824 net825 VGND VGND VPWR VPWR net824 sky130_fd_sc_hd__clkbuf_1
X_22518_ net4390 net4380 net4316 net4346 VGND VGND VPWR VPWR _02518_ sky130_fd_sc_hd__or4_1
XFILLER_0_52_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23498_ net1670 net1667 VGND VGND VPWR VPWR _03367_ sky130_fd_sc_hd__xnor2_1
Xwire835 _06240_ VGND VGND VPWR VPWR net835 sky130_fd_sc_hd__buf_1
Xmax_length411 _02180_ VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__clkbuf_1
Xwire846 _05549_ VGND VGND VPWR VPWR net846 sky130_fd_sc_hd__buf_1
Xmax_length422 _10407_ VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire868 _11978_ VGND VGND VPWR VPWR net868 sky130_fd_sc_hd__buf_1
XFILLER_0_161_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13251_ _05518_ _05523_ VGND VGND VPWR VPWR _05524_ sky130_fd_sc_hd__xnor2_1
X_22449_ _02341_ _02377_ _02378_ VGND VGND VPWR VPWR _02451_ sky130_fd_sc_hd__o21ai_2
X_25237_ clknet_leaf_23_clk _00010_ net8582 VGND VGND VPWR VPWR pid_q.state\[4\] sky130_fd_sc_hd__dfrtp_1
Xwire879 _08568_ VGND VGND VPWR VPWR net879 sky130_fd_sc_hd__buf_1
X_13182_ _05366_ _05367_ _05368_ VGND VGND VPWR VPWR _05455_ sky130_fd_sc_hd__a21o_1
X_25168_ clknet_leaf_55_clk _00057_ net8728 VGND VGND VPWR VPWR svm0.periodTop\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire4120 net4122 VGND VGND VPWR VPWR net4120 sky130_fd_sc_hd__buf_1
Xwire4131 net4132 VGND VGND VPWR VPWR net4131 sky130_fd_sc_hd__buf_1
X_24119_ _03979_ _03980_ VGND VGND VPWR VPWR _03981_ sky130_fd_sc_hd__xor2_2
XFILLER_0_20_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4142 _07023_ VGND VGND VPWR VPWR net4142 sky130_fd_sc_hd__buf_1
X_25099_ net1994 _04840_ _04841_ VGND VGND VPWR VPWR _04843_ sky130_fd_sc_hd__o21ai_1
X_17990_ _09777_ _09778_ _09779_ _09839_ _09840_ VGND VGND VPWR VPWR _09841_ sky130_fd_sc_hd__a311o_1
Xwire4153 net4154 VGND VGND VPWR VPWR net4153 sky130_fd_sc_hd__buf_1
XFILLER_0_20_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4164 net4165 VGND VGND VPWR VPWR net4164 sky130_fd_sc_hd__buf_1
Xwire3430 _07485_ VGND VGND VPWR VPWR net3430 sky130_fd_sc_hd__buf_1
Xwire4175 net4176 VGND VGND VPWR VPWR net4175 sky130_fd_sc_hd__buf_1
X_16941_ net1827 VGND VGND VPWR VPWR _08905_ sky130_fd_sc_hd__clkbuf_1
Xwire3441 _07353_ VGND VGND VPWR VPWR net3441 sky130_fd_sc_hd__buf_1
Xwire4186 net4187 VGND VGND VPWR VPWR net4186 sky130_fd_sc_hd__buf_1
Xwire4197 _06977_ VGND VGND VPWR VPWR net4197 sky130_fd_sc_hd__buf_1
Xwire2740 net2741 VGND VGND VPWR VPWR net2740 sky130_fd_sc_hd__buf_1
X_19660_ net3142 net3291 net2504 VGND VGND VPWR VPWR _11496_ sky130_fd_sc_hd__and3_1
Xwire3485 _07150_ VGND VGND VPWR VPWR net3485 sky130_fd_sc_hd__clkbuf_1
X_16872_ net5992 net4057 _08836_ VGND VGND VPWR VPWR _08837_ sky130_fd_sc_hd__mux2_1
Xwire2751 net2752 VGND VGND VPWR VPWR net2751 sky130_fd_sc_hd__buf_1
Xwire2762 net2763 VGND VGND VPWR VPWR net2762 sky130_fd_sc_hd__buf_1
Xwire2773 net2774 VGND VGND VPWR VPWR net2773 sky130_fd_sc_hd__clkbuf_1
X_18611_ net6377 net422 _10458_ VGND VGND VPWR VPWR _10459_ sky130_fd_sc_hd__a21o_1
Xwire2784 net2785 VGND VGND VPWR VPWR net2784 sky130_fd_sc_hd__buf_1
X_15823_ _07794_ _07796_ _07792_ VGND VGND VPWR VPWR _07893_ sky130_fd_sc_hd__o21ba_1
X_19591_ _11375_ _11417_ VGND VGND VPWR VPWR _11428_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18542_ net3930 VGND VGND VPWR VPWR _10391_ sky130_fd_sc_hd__clkbuf_1
X_15754_ _07645_ _07734_ net778 VGND VGND VPWR VPWR _07825_ sky130_fd_sc_hd__a21boi_1
X_12966_ _05237_ _05238_ net1155 VGND VGND VPWR VPWR _05239_ sky130_fd_sc_hd__mux2_1
X_14705_ net7149 _06848_ VGND VGND VPWR VPWR _06849_ sky130_fd_sc_hd__xnor2_1
X_18473_ net1773 _10243_ VGND VGND VPWR VPWR _10323_ sky130_fd_sc_hd__or2b_1
X_15685_ _07752_ _07755_ VGND VGND VPWR VPWR _07756_ sky130_fd_sc_hd__xnor2_2
X_12897_ net7737 net1617 VGND VGND VPWR VPWR _05170_ sky130_fd_sc_hd__nand2_1
X_17424_ net2615 _09324_ VGND VGND VPWR VPWR _00388_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14636_ net3629 VGND VGND VPWR VPWR _06801_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_184_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17355_ net6658 net4253 VGND VGND VPWR VPWR _09268_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14567_ net7260 net3640 _06730_ VGND VGND VPWR VPWR _06744_ sky130_fd_sc_hd__o21a_1
X_16306_ _08359_ _08369_ VGND VGND VPWR VPWR _08370_ sky130_fd_sc_hd__xnor2_1
X_13518_ _05785_ _05788_ VGND VGND VPWR VPWR _05789_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_181_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17286_ net6727 net6719 _09197_ _09200_ VGND VGND VPWR VPWR _09201_ sky130_fd_sc_hd__or4_1
X_14498_ net7313 net5270 VGND VGND VPWR VPWR _06681_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_36_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19025_ _10809_ _10835_ _10861_ VGND VGND VPWR VPWR _10862_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_28_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16237_ net491 _08301_ VGND VGND VPWR VPWR _08302_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13449_ _05719_ _05720_ _05621_ _05622_ VGND VGND VPWR VPWR _05722_ sky130_fd_sc_hd__and4_1
XFILLER_0_140_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16168_ _08231_ _08233_ VGND VGND VPWR VPWR _08234_ sky130_fd_sc_hd__xor2_1
XFILLER_0_23_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout4570 net4577 VGND VGND VPWR VPWR net4570 sky130_fd_sc_hd__buf_1
X_15119_ net3603 _07192_ VGND VGND VPWR VPWR _07193_ sky130_fd_sc_hd__nor2_1
X_16099_ net2234 _08163_ _08164_ VGND VGND VPWR VPWR _08165_ sky130_fd_sc_hd__a21oi_2
X_19927_ _11757_ _11758_ VGND VGND VPWR VPWR _11759_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_177_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19858_ _11689_ _11690_ VGND VGND VPWR VPWR _11691_ sky130_fd_sc_hd__xor2_1
XFILLER_0_183_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18809_ _10596_ _10598_ _10595_ VGND VGND VPWR VPWR _10653_ sky130_fd_sc_hd__a21o_1
X_19789_ _11584_ _11592_ _11622_ VGND VGND VPWR VPWR _11623_ sky130_fd_sc_hd__a21oi_1
X_21820_ _01748_ _01775_ _01828_ VGND VGND VPWR VPWR _01829_ sky130_fd_sc_hd__o21ai_1
X_21751_ _01755_ _01760_ VGND VGND VPWR VPWR _01761_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_90_clk clknet_4_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_90_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_175_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20702_ _12472_ _12475_ VGND VGND VPWR VPWR _12476_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_176_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24470_ net7522 _04263_ net236 net7465 net290 VGND VGND VPWR VPWR _04328_ sky130_fd_sc_hd__a221o_1
X_21682_ _01691_ _01692_ VGND VGND VPWR VPWR _01693_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8419 net8414 VGND VGND VPWR VPWR net8419 sky130_fd_sc_hd__buf_1
X_23421_ _03208_ _03209_ _03290_ VGND VGND VPWR VPWR _03291_ sky130_fd_sc_hd__a21oi_2
Xclkbuf_4_9__f_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_4_9__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20633_ _12411_ _12412_ VGND VGND VPWR VPWR _12413_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7707 net7709 VGND VGND VPWR VPWR net7707 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire7718 net7721 VGND VGND VPWR VPWR net7718 sky130_fd_sc_hd__buf_1
Xmax_length3405 net3406 VGND VGND VPWR VPWR net3405 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_190_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23352_ _02940_ _02942_ _02941_ VGND VGND VPWR VPWR _03222_ sky130_fd_sc_hd__o21a_1
Xwire7729 net7730 VGND VGND VPWR VPWR net7729 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20564_ _12333_ _12336_ _12344_ VGND VGND VPWR VPWR _12348_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length3449 net3450 VGND VGND VPWR VPWR net3449 sky130_fd_sc_hd__buf_1
XFILLER_0_150_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22303_ net2473 _02305_ _02306_ _02300_ VGND VGND VPWR VPWR _02307_ sky130_fd_sc_hd__a31o_1
XFILLER_0_33_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23283_ _03107_ _03110_ net3060 VGND VGND VPWR VPWR _03153_ sky130_fd_sc_hd__o21a_1
XFILLER_0_131_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20495_ _12280_ _12281_ _12282_ VGND VGND VPWR VPWR _12283_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_132_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22234_ _02152_ _02155_ _02238_ VGND VGND VPWR VPWR _02239_ sky130_fd_sc_hd__a21o_1
X_25022_ _04774_ _04775_ VGND VGND VPWR VPWR _04776_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22165_ _02169_ _02170_ VGND VGND VPWR VPWR _02171_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21116_ _01084_ _01131_ VGND VGND VPWR VPWR _01132_ sky130_fd_sc_hd__xnor2_1
Xwire2003 net2004 VGND VGND VPWR VPWR net2003 sky130_fd_sc_hd__clkbuf_2
Xwire2014 net2015 VGND VGND VPWR VPWR net2014 sky130_fd_sc_hd__clkbuf_1
X_22096_ pid_d.prev_error\[9\] net5967 VGND VGND VPWR VPWR _02103_ sky130_fd_sc_hd__xnor2_1
Xwire2025 _03963_ VGND VGND VPWR VPWR net2025 sky130_fd_sc_hd__buf_1
Xwire2036 _02694_ VGND VGND VPWR VPWR net2036 sky130_fd_sc_hd__dlymetal6s2s_1
X_25924_ clknet_leaf_1_clk _00797_ net8404 VGND VGND VPWR VPWR pid_d.prev_int\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1302 _06522_ VGND VGND VPWR VPWR net1302 sky130_fd_sc_hd__buf_1
X_21047_ net1731 _01061_ _01062_ VGND VGND VPWR VPWR _01063_ sky130_fd_sc_hd__a21o_1
Xwire2047 net2048 VGND VGND VPWR VPWR net2047 sky130_fd_sc_hd__buf_1
Xwire2058 net2059 VGND VGND VPWR VPWR net2058 sky130_fd_sc_hd__clkbuf_2
Xwire1324 net1325 VGND VGND VPWR VPWR net1324 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2069 _01711_ VGND VGND VPWR VPWR net2069 sky130_fd_sc_hd__buf_1
Xwire1335 _05133_ VGND VGND VPWR VPWR net1335 sky130_fd_sc_hd__clkbuf_1
Xwire1346 _04921_ VGND VGND VPWR VPWR net1346 sky130_fd_sc_hd__buf_1
Xwire1357 net1358 VGND VGND VPWR VPWR net1357 sky130_fd_sc_hd__buf_1
X_25855_ clknet_leaf_23_clk _00728_ net8586 VGND VGND VPWR VPWR pid_q.mult0.b\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1368 net1369 VGND VGND VPWR VPWR net1368 sky130_fd_sc_hd__buf_1
Xwire1379 _04072_ VGND VGND VPWR VPWR net1379 sky130_fd_sc_hd__buf_1
X_24806_ net7955 _04629_ VGND VGND VPWR VPWR _04630_ sky130_fd_sc_hd__xor2_1
X_12820_ _05089_ _05092_ VGND VGND VPWR VPWR _05093_ sky130_fd_sc_hd__xnor2_2
X_25786_ clknet_leaf_58_clk _00659_ net8712 VGND VGND VPWR VPWR matmul0.beta_pass\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_22998_ net3758 VGND VGND VPWR VPWR _02868_ sky130_fd_sc_hd__inv_2
X_24737_ pid_q.curr_error\[5\] net1371 net1365 net1009 VGND VGND VPWR VPWR _00702_
+ sky130_fd_sc_hd__a22o_1
X_12751_ _05004_ net851 VGND VGND VPWR VPWR _05024_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21949_ net5839 net5420 net5395 net3776 _01956_ VGND VGND VPWR VPWR _01957_ sky130_fd_sc_hd__a41o_1
XFILLER_0_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8803 net8808 VGND VGND VPWR VPWR net8803 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_167_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_81_clk clknet_4_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_81_clk sky130_fd_sc_hd__clkbuf_16
Xfanout8814 net8856 VGND VGND VPWR VPWR net8814 sky130_fd_sc_hd__buf_1
XFILLER_0_38_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15470_ _07343_ _07344_ net1542 VGND VGND VPWR VPWR _07544_ sky130_fd_sc_hd__and3_1
X_24668_ net9144 net1375 _04516_ VGND VGND VPWR VPWR _00686_ sky130_fd_sc_hd__a21o_1
X_12682_ _04945_ net1008 _04954_ VGND VGND VPWR VPWR _04955_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_166_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14421_ matmul0.beta_pass\[7\] net1293 net2889 net4436 _06619_ VGND VGND VPWR VPWR
+ _06620_ sky130_fd_sc_hd__a221o_1
Xfanout8869 net8873 VGND VGND VPWR VPWR net8869 sky130_fd_sc_hd__buf_1
Xwire8920 net8921 VGND VGND VPWR VPWR net8920 sky130_fd_sc_hd__clkbuf_1
X_23619_ net696 _03473_ VGND VGND VPWR VPWR _03486_ sky130_fd_sc_hd__nand2_1
Xwire8931 net111 VGND VGND VPWR VPWR net8931 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length5363 pid_d.out\[6\] VGND VGND VPWR VPWR net5363 sky130_fd_sc_hd__buf_1
Xwire8942 net8943 VGND VGND VPWR VPWR net8942 sky130_fd_sc_hd__clkbuf_1
X_24599_ net5170 _02866_ net2433 _04454_ VGND VGND VPWR VPWR _00679_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8953 net1 VGND VGND VPWR VPWR net8953 sky130_fd_sc_hd__dlymetal6s2s_1
X_17140_ net5988 net2597 net3343 net3305 VGND VGND VPWR VPWR _09094_ sky130_fd_sc_hd__a22o_1
Xwire610 _10260_ VGND VGND VPWR VPWR net610 sky130_fd_sc_hd__clkbuf_1
X_14352_ net8210 net3646 VGND VGND VPWR VPWR _06566_ sky130_fd_sc_hd__and2_1
Xwire621 _05937_ VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__buf_1
Xwire632 _04443_ VGND VGND VPWR VPWR net632 sky130_fd_sc_hd__clkbuf_1
Xwire643 net644 VGND VGND VPWR VPWR net643 sky130_fd_sc_hd__clkbuf_1
X_13303_ _05491_ _05574_ _05575_ VGND VGND VPWR VPWR _05576_ sky130_fd_sc_hd__a21o_1
XFILLER_0_122_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17071_ net3332 net6474 VGND VGND VPWR VPWR _09029_ sky130_fd_sc_hd__nor2_1
Xwire654 net655 VGND VGND VPWR VPWR net654 sky130_fd_sc_hd__clkbuf_1
X_14283_ net8118 net2902 net2265 net7855 VGND VGND VPWR VPWR _00054_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire665 net666 VGND VGND VPWR VPWR net665 sky130_fd_sc_hd__clkbuf_1
Xwire676 _06707_ VGND VGND VPWR VPWR net676 sky130_fd_sc_hd__clkbuf_1
Xwire687 _04651_ VGND VGND VPWR VPWR net687 sky130_fd_sc_hd__clkbuf_1
Xwire698 _01921_ VGND VGND VPWR VPWR net698 sky130_fd_sc_hd__clkbuf_1
X_16022_ _08007_ _08082_ VGND VGND VPWR VPWR _08089_ sky130_fd_sc_hd__nand2_1
X_13234_ net7745 net2321 net2317 VGND VGND VPWR VPWR _05507_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13165_ _05434_ _05435_ _05436_ _05437_ VGND VGND VPWR VPWR _05438_ sky130_fd_sc_hd__a211o_1
XFILLER_0_23_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13096_ _05367_ _05368_ VGND VGND VPWR VPWR _05369_ sky130_fd_sc_hd__xnor2_1
X_17973_ _09790_ net1213 VGND VGND VPWR VPWR _09824_ sky130_fd_sc_hd__xnor2_1
Xwire3260 _09633_ VGND VGND VPWR VPWR net3260 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_97_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3271 net3272 VGND VGND VPWR VPWR net3271 sky130_fd_sc_hd__buf_1
X_16924_ net6420 _08886_ _08887_ VGND VGND VPWR VPWR _08888_ sky130_fd_sc_hd__a21bo_1
X_19712_ net653 _11424_ _11481_ _11547_ VGND VGND VPWR VPWR _11548_ sky130_fd_sc_hd__a31o_1
Xwire3293 net3294 VGND VGND VPWR VPWR net3293 sky130_fd_sc_hd__clkbuf_1
X_16855_ net6082 net6055 net6501 VGND VGND VPWR VPWR _08820_ sky130_fd_sc_hd__mux2_1
X_19643_ _11472_ _11479_ VGND VGND VPWR VPWR _11480_ sky130_fd_sc_hd__xnor2_1
Xwire2581 net2582 VGND VGND VPWR VPWR net2581 sky130_fd_sc_hd__buf_1
X_15806_ _07872_ _07875_ VGND VGND VPWR VPWR _07876_ sky130_fd_sc_hd__xnor2_2
X_19574_ net3146 net3142 VGND VGND VPWR VPWR _11411_ sky130_fd_sc_hd__nor2_1
Xwire1880 _07286_ VGND VGND VPWR VPWR net1880 sky130_fd_sc_hd__clkbuf_2
Xwire1891 _07209_ VGND VGND VPWR VPWR net1891 sky130_fd_sc_hd__clkbuf_1
X_16786_ net7589 matmul0.a\[12\] net3372 VGND VGND VPWR VPWR _08783_ sky130_fd_sc_hd__mux2_1
X_13998_ _06167_ _06261_ _06262_ VGND VGND VPWR VPWR _06263_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_99_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18525_ _10371_ _10372_ net6833 VGND VGND VPWR VPWR _10374_ sky130_fd_sc_hd__a21oi_1
X_15737_ _07647_ _07649_ _07648_ VGND VGND VPWR VPWR _07808_ sky130_fd_sc_hd__a21bo_1
X_12949_ _05214_ net1593 VGND VGND VPWR VPWR _05222_ sky130_fd_sc_hd__nand2_1
XFILLER_0_158_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_72_clk clknet_4_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18456_ net3229 _10305_ VGND VGND VPWR VPWR _10306_ sky130_fd_sc_hd__xnor2_1
X_15668_ _07737_ _07739_ VGND VGND VPWR VPWR _07740_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17407_ svm0.delta\[10\] VGND VGND VPWR VPWR _09311_ sky130_fd_sc_hd__inv_2
Xclkbuf_2_1_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1_0_clk sky130_fd_sc_hd__clkbuf_8
X_14619_ net1622 _06786_ clarke_done VGND VGND VPWR VPWR _06790_ sky130_fd_sc_hd__a21o_1
X_18387_ _10231_ _10232_ _10236_ _10237_ VGND VGND VPWR VPWR _10238_ sky130_fd_sc_hd__o211ai_1
X_15599_ net3531 net2725 VGND VGND VPWR VPWR _07671_ sky130_fd_sc_hd__nor2_1
X_17338_ net6698 net7661 VGND VGND VPWR VPWR _09252_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17269_ net2159 net191 net1797 net9136 VGND VGND VPWR VPWR _00363_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_183_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19008_ net6268 _10828_ net3202 VGND VGND VPWR VPWR _10845_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_178_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20280_ net1835 net2091 net8055 VGND VGND VPWR VPWR _12087_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold17 matmul0.matmul_stage_inst.a\[8\] VGND VGND VPWR VPWR net8970 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 matmul0.matmul_stage_inst.a\[3\] VGND VGND VPWR VPWR net8981 sky130_fd_sc_hd__dlygate4sd3_1
X_23970_ _03742_ _03833_ VGND VGND VPWR VPWR _03834_ sky130_fd_sc_hd__xnor2_1
Xhold39 pid_d.iterate_enable VGND VGND VPWR VPWR net8992 sky130_fd_sc_hd__dlygate4sd3_1
X_22921_ _02811_ VGND VGND VPWR VPWR _02812_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25640_ clknet_leaf_102_clk _00513_ net8366 VGND VGND VPWR VPWR cordic0.vec\[0\]\[12\]
+ sky130_fd_sc_hd__dfstp_1
X_22852_ pid_d.out\[4\] net3065 _02750_ net8897 VGND VGND VPWR VPWR _00636_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21803_ pid_d.prev_error\[6\] net5968 VGND VGND VPWR VPWR _01813_ sky130_fd_sc_hd__xnor2_1
X_25571_ clknet_leaf_98_clk _00444_ net8381 VGND VGND VPWR VPWR cordic0.sin\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22783_ _02699_ VGND VGND VPWR VPWR _00618_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_63_clk clknet_4_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_63_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24522_ net792 _04315_ _04376_ _04268_ VGND VGND VPWR VPWR _04379_ sky130_fd_sc_hd__o22a_1
X_21734_ net1173 _01706_ _01743_ VGND VGND VPWR VPWR _01744_ sky130_fd_sc_hd__o21a_2
Xwire8205 net8206 VGND VGND VPWR VPWR net8205 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8216 net31 VGND VGND VPWR VPWR net8216 sky130_fd_sc_hd__clkbuf_1
X_24453_ _04229_ _04233_ _04310_ VGND VGND VPWR VPWR _04311_ sky130_fd_sc_hd__a21o_1
Xwire8227 net8228 VGND VGND VPWR VPWR net8227 sky130_fd_sc_hd__clkbuf_1
X_21665_ _01674_ _01675_ VGND VGND VPWR VPWR _01676_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8238 net8239 VGND VGND VPWR VPWR net8238 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7504 net7505 VGND VGND VPWR VPWR net7504 sky130_fd_sc_hd__buf_1
XFILLER_0_4_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8249 net8250 VGND VGND VPWR VPWR net8249 sky130_fd_sc_hd__clkbuf_1
X_23404_ net4575 net5080 VGND VGND VPWR VPWR _03274_ sky130_fd_sc_hd__nand2_1
Xwire7515 net7507 VGND VGND VPWR VPWR net7515 sky130_fd_sc_hd__buf_1
XFILLER_0_152_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7526 net7527 VGND VGND VPWR VPWR net7526 sky130_fd_sc_hd__buf_1
X_20616_ net1740 _12367_ net1396 VGND VGND VPWR VPWR _12397_ sky130_fd_sc_hd__or3b_1
X_24384_ _04240_ net929 VGND VGND VPWR VPWR _04243_ sky130_fd_sc_hd__nor2_1
X_21596_ net5928 net5909 net5951 VGND VGND VPWR VPWR _01608_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7537 net7538 VGND VGND VPWR VPWR net7537 sky130_fd_sc_hd__clkbuf_1
Xwire7548 net7549 VGND VGND VPWR VPWR net7548 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire6814 net6812 VGND VGND VPWR VPWR net6814 sky130_fd_sc_hd__buf_1
XFILLER_0_85_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7559 net7560 VGND VGND VPWR VPWR net7559 sky130_fd_sc_hd__clkbuf_1
X_23335_ _03201_ _03204_ VGND VGND VPWR VPWR _03205_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_149_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20547_ _12330_ _12331_ net2082 VGND VGND VPWR VPWR _12332_ sky130_fd_sc_hd__a21bo_1
Xwire6836 net6838 VGND VGND VPWR VPWR net6836 sky130_fd_sc_hd__buf_1
XFILLER_0_104_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6847 net6848 VGND VGND VPWR VPWR net6847 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire6869 net6866 VGND VGND VPWR VPWR net6869 sky130_fd_sc_hd__buf_1
X_23266_ _03134_ _03135_ VGND VGND VPWR VPWR _03136_ sky130_fd_sc_hd__nand2_1
X_20478_ net7147 net7129 net7113 net7088 net6512 net6489 VGND VGND VPWR VPWR _12267_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25005_ net4474 net5183 pid_q.out\[1\] net5181 VGND VGND VPWR VPWR _04761_ sky130_fd_sc_hd__a22o_1
X_22217_ _02128_ _02133_ _02126_ VGND VGND VPWR VPWR _02222_ sky130_fd_sc_hd__a21bo_1
X_23197_ _03064_ _03066_ VGND VGND VPWR VPWR _03067_ sky130_fd_sc_hd__nor2_1
X_22148_ _02045_ _02047_ _02153_ VGND VGND VPWR VPWR _02154_ sky130_fd_sc_hd__o21a_1
X_22079_ net1717 _01980_ VGND VGND VPWR VPWR _02086_ sky130_fd_sc_hd__nand2_1
X_14970_ net4139 _07027_ VGND VGND VPWR VPWR _07044_ sky130_fd_sc_hd__nor2_1
Xwire1110 net1111 VGND VGND VPWR VPWR net1110 sky130_fd_sc_hd__clkbuf_1
Xwire1121 net1123 VGND VGND VPWR VPWR net1121 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_22_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13921_ net7668 net1944 net2293 VGND VGND VPWR VPWR _06187_ sky130_fd_sc_hd__and3_1
Xwire1132 _05557_ VGND VGND VPWR VPWR net1132 sky130_fd_sc_hd__buf_1
X_25907_ clknet_leaf_60_clk _00780_ net8691 VGND VGND VPWR VPWR pid_q.out\[3\] sky130_fd_sc_hd__dfrtp_1
Xwire1143 _05174_ VGND VGND VPWR VPWR net1143 sky130_fd_sc_hd__buf_1
Xwire1165 _03545_ VGND VGND VPWR VPWR net1165 sky130_fd_sc_hd__buf_1
X_16640_ matmul0.alpha_pass\[3\] net2202 net6552 VGND VGND VPWR VPWR _08678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13852_ _06116_ _06118_ VGND VGND VPWR VPWR _06119_ sky130_fd_sc_hd__xnor2_1
X_25838_ clknet_leaf_31_clk _00711_ net8684 VGND VGND VPWR VPWR pid_q.curr_error\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1187 _00913_ VGND VGND VPWR VPWR net1187 sky130_fd_sc_hd__buf_1
Xwire1198 _10362_ VGND VGND VPWR VPWR net1198 sky130_fd_sc_hd__clkbuf_1
X_12803_ _04955_ _05075_ _05074_ VGND VGND VPWR VPWR _05076_ sky130_fd_sc_hd__a21o_1
X_16571_ _08550_ _08554_ _08623_ _08629_ VGND VGND VPWR VPWR _08630_ sky130_fd_sc_hd__a31o_1
X_13783_ net909 net781 VGND VGND VPWR VPWR _06051_ sky130_fd_sc_hd__or2_1
X_25769_ clknet_leaf_26_clk _00642_ net8576 VGND VGND VPWR VPWR pid_d.out\[10\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_54_clk clknet_4_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_16
X_18310_ net7072 _09675_ VGND VGND VPWR VPWR _10161_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15522_ net2717 net3537 VGND VGND VPWR VPWR _07595_ sky130_fd_sc_hd__nor2_1
X_12734_ net7917 net1350 _05005_ _05006_ VGND VGND VPWR VPWR _05007_ sky130_fd_sc_hd__a22o_1
X_19290_ net3205 VGND VGND VPWR VPWR _11127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout8622 net8643 VGND VGND VPWR VPWR net8622 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_84_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8633 net8826 VGND VGND VPWR VPWR net8633 sky130_fd_sc_hd__clkbuf_1
X_18241_ net7063 _10037_ net2564 _10091_ VGND VGND VPWR VPWR _10092_ sky130_fd_sc_hd__o31a_1
X_15453_ net2807 net3555 VGND VGND VPWR VPWR _07527_ sky130_fd_sc_hd__nor2_1
X_12665_ _04936_ _04937_ net7836 net1346 VGND VGND VPWR VPWR _04938_ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout8677 net8699 VGND VGND VPWR VPWR net8677 sky130_fd_sc_hd__buf_1
XFILLER_0_26_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14404_ _06605_ matmul0.b_in\[3\] net898 VGND VGND VPWR VPWR _06607_ sky130_fd_sc_hd__mux2_1
Xwire8750 net8747 VGND VGND VPWR VPWR net8750 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_155_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length5182 pid_q.curr_int\[1\] VGND VGND VPWR VPWR net5182 sky130_fd_sc_hd__buf_1
X_18172_ _09842_ net768 net817 _10022_ VGND VGND VPWR VPWR _10023_ sky130_fd_sc_hd__a31o_1
X_15384_ net990 _07457_ VGND VGND VPWR VPWR _07458_ sky130_fd_sc_hd__xnor2_1
Xwire8772 net8769 VGND VGND VPWR VPWR net8772 sky130_fd_sc_hd__buf_1
X_12596_ net4292 VGND VGND VPWR VPWR _04877_ sky130_fd_sc_hd__buf_1
Xmax_length4470 pid_q.out\[1\] VGND VGND VPWR VPWR net4470 sky130_fd_sc_hd__clkbuf_1
Xwire8783 net8781 VGND VGND VPWR VPWR net8783 sky130_fd_sc_hd__buf_1
X_17123_ _09068_ _09078_ net3350 VGND VGND VPWR VPWR _09079_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8794 net8795 VGND VGND VPWR VPWR net8794 sky130_fd_sc_hd__clkbuf_1
Xwire440 net441 VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__buf_1
X_14335_ _06553_ VGND VGND VPWR VPWR _00070_ sky130_fd_sc_hd__clkbuf_1
Xwire451 _05933_ VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__clkbuf_2
Xwire462 net463 VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__clkbuf_1
Xwire473 net474 VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__buf_1
XFILLER_0_150_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17054_ net1804 net1483 _08952_ VGND VGND VPWR VPWR _09013_ sky130_fd_sc_hd__o21ai_1
Xwire484 net485 VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__clkbuf_1
X_14266_ net59 net2931 net2278 net9004 VGND VGND VPWR VPWR _00039_ sky130_fd_sc_hd__a22o_1
Xwire495 net496 VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__clkbuf_1
X_16005_ _08068_ _08072_ VGND VGND VPWR VPWR _08073_ sky130_fd_sc_hd__xnor2_2
X_13217_ _05488_ _05489_ VGND VGND VPWR VPWR _05490_ sky130_fd_sc_hd__xor2_1
X_14197_ _06401_ _06419_ _06402_ VGND VGND VPWR VPWR _06457_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13148_ net4261 net2302 net2298 VGND VGND VPWR VPWR _05421_ sky130_fd_sc_hd__or3_1
XFILLER_0_148_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13079_ _05290_ _05296_ _05351_ net4259 _05287_ VGND VGND VPWR VPWR _05352_ sky130_fd_sc_hd__o221a_1
X_17956_ _09805_ _09806_ VGND VGND VPWR VPWR _09807_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3090 net3091 VGND VGND VPWR VPWR net3090 sky130_fd_sc_hd__buf_1
XFILLER_0_174_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16907_ cordic0.slte0.opA\[6\] net6413 VGND VGND VPWR VPWR _08871_ sky130_fd_sc_hd__or2b_1
X_17887_ net6966 net7005 VGND VGND VPWR VPWR _09738_ sky130_fd_sc_hd__nand2_1
XFILLER_0_174_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19626_ net6225 _11401_ _11462_ VGND VGND VPWR VPWR _11463_ sky130_fd_sc_hd__nand3_1
X_16838_ net6424 matmul0.sin\[7\] net3366 VGND VGND VPWR VPWR _08810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19557_ _10938_ _11393_ net2513 net6252 VGND VGND VPWR VPWR _11394_ sky130_fd_sc_hd__a211o_1
X_16769_ matmul0.a_in\[4\] matmul0.a\[4\] net3378 VGND VGND VPWR VPWR _08774_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_45_clk clknet_4_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18508_ net3229 _10304_ net3941 VGND VGND VPWR VPWR _10357_ sky130_fd_sc_hd__a21o_1
X_19488_ _11323_ _11324_ VGND VGND VPWR VPWR _11325_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18439_ _10284_ _10287_ VGND VGND VPWR VPWR _10289_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21450_ _01348_ _01462_ net5638 VGND VGND VPWR VPWR _01463_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20401_ _12187_ _12197_ _12198_ VGND VGND VPWR VPWR _12199_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_43_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21381_ _01392_ net1181 VGND VGND VPWR VPWR _01395_ sky130_fd_sc_hd__xor2_1
XFILLER_0_189_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23120_ _02981_ _02989_ VGND VGND VPWR VPWR _02990_ sky130_fd_sc_hd__xnor2_2
X_20332_ _12134_ VGND VGND VPWR VPWR _12135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4708 net4709 VGND VGND VPWR VPWR net4708 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4719 net4720 VGND VGND VPWR VPWR net4719 sky130_fd_sc_hd__buf_1
XFILLER_0_113_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23051_ _02889_ _02908_ _02920_ VGND VGND VPWR VPWR _02921_ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20263_ _12074_ cordic0.slte0.opB\[13\] net2531 VGND VGND VPWR VPWR _12075_ sky130_fd_sc_hd__mux2_1
X_22002_ _02008_ _01910_ _02009_ VGND VGND VPWR VPWR _02010_ sky130_fd_sc_hd__a21o_1
XFILLER_0_179_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20194_ net952 _11995_ net867 VGND VGND VPWR VPWR _12019_ sky130_fd_sc_hd__a21oi_1
Xinput107 pid_d_data[4] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_1
Xinput118 pid_q_addr[13] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_1
Xinput129 pid_q_addr[9] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_1
X_23953_ _03811_ _03816_ VGND VGND VPWR VPWR _03817_ sky130_fd_sc_hd__xnor2_2
X_22904_ _02109_ _02787_ _02796_ VGND VGND VPWR VPWR _02797_ sky130_fd_sc_hd__a21o_1
X_23884_ _03641_ _03650_ net855 VGND VGND VPWR VPWR _03749_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25623_ clknet_leaf_116_clk _00496_ net8329 VGND VGND VPWR VPWR cordic0.slte0.opA\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_22835_ net5365 VGND VGND VPWR VPWR _02735_ sky130_fd_sc_hd__inv_2
XFILLER_0_196_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_36_clk clknet_4_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_6_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25554_ clknet_leaf_78_clk net3003 net8439 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_22766_ pid_d.ki\[13\] _02688_ net2038 VGND VGND VPWR VPWR _02689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24505_ net4582 net3045 _04273_ VGND VGND VPWR VPWR _04362_ sky130_fd_sc_hd__or3b_1
XFILLER_0_93_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8002 net8003 VGND VGND VPWR VPWR net8002 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21717_ pid_d.curr_error\[4\] VGND VGND VPWR VPWR _01728_ sky130_fd_sc_hd__inv_2
X_25485_ clknet_leaf_45_clk _00365_ net8788 VGND VGND VPWR VPWR svm0.tA\[7\] sky130_fd_sc_hd__dfrtp_1
Xwire8013 net8014 VGND VGND VPWR VPWR net8013 sky130_fd_sc_hd__clkbuf_1
Xwire8024 net8025 VGND VGND VPWR VPWR net8024 sky130_fd_sc_hd__clkbuf_1
X_22697_ _02639_ net5496 net2451 VGND VGND VPWR VPWR _02640_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8035 net8036 VGND VGND VPWR VPWR net8035 sky130_fd_sc_hd__clkbuf_1
Xwire7301 matmul0.alpha_pass\[6\] VGND VGND VPWR VPWR net7301 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24436_ net4918 _04290_ _04291_ _04293_ net4896 VGND VGND VPWR VPWR _04294_ sky130_fd_sc_hd__a32o_1
Xwire7312 net7316 VGND VGND VPWR VPWR net7312 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21648_ _01557_ _01559_ _01558_ VGND VGND VPWR VPWR _01659_ sky130_fd_sc_hd__o21a_1
Xwire8057 net8054 VGND VGND VPWR VPWR net8057 sky130_fd_sc_hd__clkbuf_2
Xwire8068 net8064 VGND VGND VPWR VPWR net8068 sky130_fd_sc_hd__clkbuf_1
Xwire7323 net7328 VGND VGND VPWR VPWR net7323 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8079 net8080 VGND VGND VPWR VPWR net8079 sky130_fd_sc_hd__clkbuf_1
Xwire7334 net7335 VGND VGND VPWR VPWR net7334 sky130_fd_sc_hd__clkbuf_1
Xwire6600 net6601 VGND VGND VPWR VPWR net6600 sky130_fd_sc_hd__buf_1
XFILLER_0_105_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7345 net7346 VGND VGND VPWR VPWR net7345 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7356 net7357 VGND VGND VPWR VPWR net7356 sky130_fd_sc_hd__buf_1
X_24367_ _04222_ _04225_ VGND VGND VPWR VPWR _04226_ sky130_fd_sc_hd__xnor2_1
Xwire7367 net7374 VGND VGND VPWR VPWR net7367 sky130_fd_sc_hd__clkbuf_1
X_21579_ _01484_ _01485_ _01590_ VGND VGND VPWR VPWR _01591_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_50_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6633 net6636 VGND VGND VPWR VPWR net6633 sky130_fd_sc_hd__clkbuf_1
Xmax_length2331 net2332 VGND VGND VPWR VPWR net2331 sky130_fd_sc_hd__buf_1
Xwire7378 net7379 VGND VGND VPWR VPWR net7378 sky130_fd_sc_hd__buf_1
X_14120_ _06378_ _06381_ VGND VGND VPWR VPWR _06382_ sky130_fd_sc_hd__xor2_1
Xwire6644 net6641 VGND VGND VPWR VPWR net6644 sky130_fd_sc_hd__clkbuf_2
Xwire7389 net7390 VGND VGND VPWR VPWR net7389 sky130_fd_sc_hd__clkbuf_1
X_23318_ net4723 net4913 VGND VGND VPWR VPWR _03188_ sky130_fd_sc_hd__nand2_1
Xwire6655 svm0.ready VGND VGND VPWR VPWR net6655 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6666 net6667 VGND VGND VPWR VPWR net6666 sky130_fd_sc_hd__clkbuf_1
Xwire5921 net5922 VGND VGND VPWR VPWR net5921 sky130_fd_sc_hd__buf_1
X_24298_ net4624 net3044 _04090_ VGND VGND VPWR VPWR _04158_ sky130_fd_sc_hd__or3b_1
Xwire5943 net5944 VGND VGND VPWR VPWR net5943 sky130_fd_sc_hd__buf_1
Xwire6688 net6686 VGND VGND VPWR VPWR net6688 sky130_fd_sc_hd__buf_1
Xwire6699 net6700 VGND VGND VPWR VPWR net6699 sky130_fd_sc_hd__buf_1
X_14051_ _06311_ _06314_ VGND VGND VPWR VPWR _06315_ sky130_fd_sc_hd__nand2_1
Xwire5954 net5953 VGND VGND VPWR VPWR net5954 sky130_fd_sc_hd__buf_1
X_23249_ _03117_ _03118_ VGND VGND VPWR VPWR _03119_ sky130_fd_sc_hd__xnor2_2
Xwire5965 pid_d.curr_error\[13\] VGND VGND VPWR VPWR net5965 sky130_fd_sc_hd__buf_1
XFILLER_0_24_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5976 pid_d.curr_int\[9\] VGND VGND VPWR VPWR net5976 sky130_fd_sc_hd__clkbuf_2
X_13002_ _05272_ _05273_ _05270_ _05271_ VGND VGND VPWR VPWR _05275_ sky130_fd_sc_hd__o211a_1
Xwire5998 net5994 VGND VGND VPWR VPWR net5998 sky130_fd_sc_hd__buf_1
X_17810_ net6954 net6885 VGND VGND VPWR VPWR _09661_ sky130_fd_sc_hd__nand2_1
X_18790_ net6855 _10579_ _10584_ VGND VGND VPWR VPWR _10634_ sky130_fd_sc_hd__nor3_1
X_17741_ _06536_ _09594_ net6449 VGND VGND VPWR VPWR _09595_ sky130_fd_sc_hd__o21a_1
X_14953_ net6610 net7429 matmul0.matmul_stage_inst.a\[4\] net6582 VGND VGND VPWR VPWR
+ _07027_ sky130_fd_sc_hd__a22o_1
X_13904_ net7766 net1931 VGND VGND VPWR VPWR _06170_ sky130_fd_sc_hd__nand2_1
X_17672_ net4011 svm0.tA\[4\] VGND VGND VPWR VPWR _09552_ sky130_fd_sc_hd__nor2_1
X_14884_ matmul0.b\[14\] matmul0.matmul_stage_inst.f\[14\] net3605 VGND VGND VPWR
+ VPWR _06960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19411_ _11099_ _11102_ VGND VGND VPWR VPWR _11248_ sky130_fd_sc_hd__or2_1
X_16623_ _08661_ _08662_ VGND VGND VPWR VPWR _08663_ sky130_fd_sc_hd__xnor2_1
X_13835_ _06100_ _06101_ VGND VGND VPWR VPWR _06102_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_27_clk clknet_4_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_16
X_19342_ net6335 _11076_ _10812_ _11177_ VGND VGND VPWR VPWR _11179_ sky130_fd_sc_hd__and4b_1
X_16554_ net2624 net3401 net1847 net2664 VGND VGND VPWR VPWR _08613_ sky130_fd_sc_hd__a31o_1
X_13766_ _06031_ _06032_ _06025_ _06026_ VGND VGND VPWR VPWR _06034_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_57_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15505_ _07133_ _07146_ net3566 _07360_ _07577_ VGND VGND VPWR VPWR _07578_ sky130_fd_sc_hd__a32o_1
X_12717_ net7853 net1615 VGND VGND VPWR VPWR _04990_ sky130_fd_sc_hd__nand2_1
X_19273_ _10966_ _10968_ VGND VGND VPWR VPWR _11110_ sky130_fd_sc_hd__nor2_1
XFILLER_0_183_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8441 net8519 VGND VGND VPWR VPWR net8441 sky130_fd_sc_hd__clkbuf_1
X_16485_ matmul0.matmul_stage_inst.mult1\[13\] net181 net3475 VGND VGND VPWR VPWR
+ _08546_ sky130_fd_sc_hd__mux2_1
X_13697_ _05896_ _05898_ VGND VGND VPWR VPWR _05966_ sky130_fd_sc_hd__nor2_1
X_18224_ _10029_ _10073_ VGND VGND VPWR VPWR _10075_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15436_ _07506_ _07509_ VGND VGND VPWR VPWR _07510_ sky130_fd_sc_hd__xnor2_1
X_12648_ net1616 VGND VGND VPWR VPWR _04921_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18155_ _10003_ _10005_ VGND VGND VPWR VPWR _10006_ sky130_fd_sc_hd__or2_1
Xwire8591 net8592 VGND VGND VPWR VPWR net8591 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15367_ net2726 net2782 _07439_ _07440_ VGND VGND VPWR VPWR _07441_ sky130_fd_sc_hd__a31o_1
XFILLER_0_81_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12579_ net8906 VGND VGND VPWR VPWR _04865_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17106_ _09060_ _09062_ VGND VGND VPWR VPWR _09063_ sky130_fd_sc_hd__nor2_1
Xwire270 _04108_ VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__clkbuf_1
X_14318_ _06539_ VGND VGND VPWR VPWR _06540_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7890 net7891 VGND VGND VPWR VPWR net7890 sky130_fd_sc_hd__buf_1
XFILLER_0_151_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire281 _06760_ VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__buf_1
X_18086_ net7054 _09936_ VGND VGND VPWR VPWR _09937_ sky130_fd_sc_hd__nand2_1
X_15298_ _07368_ net3438 VGND VGND VPWR VPWR _07372_ sky130_fd_sc_hd__nor2_1
Xwire292 net293 VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__buf_1
XFILLER_0_68_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17037_ net7053 net967 VGND VGND VPWR VPWR _08997_ sky130_fd_sc_hd__nand2_1
X_14249_ net6477 net6467 VGND VGND VPWR VPWR _06504_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18988_ _10823_ _10824_ net6296 VGND VGND VPWR VPWR _10825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_183_Right_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17939_ _09686_ _09783_ _09789_ VGND VGND VPWR VPWR _09790_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_175_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20950_ _12526_ _00918_ _00939_ _00965_ net3830 VGND VGND VPWR VPWR _00966_ sky130_fd_sc_hd__o32a_1
XFILLER_0_191_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19609_ _11445_ VGND VGND VPWR VPWR _11446_ sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20881_ net5507 net5905 VGND VGND VPWR VPWR _00897_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_18_clk clknet_4_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_177_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22620_ net7218 _02586_ VGND VGND VPWR VPWR _02591_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22551_ net5965 net3018 net2460 VGND VGND VPWR VPWR _02538_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21502_ net1179 _01514_ VGND VGND VPWR VPWR _01515_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25270_ clknet_leaf_92_clk _00153_ net8433 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.c\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_172_Left_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22482_ net5433 net5692 VGND VGND VPWR VPWR _02483_ sky130_fd_sc_hd__and2b_1
XFILLER_0_90_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24221_ _03964_ _03966_ _03965_ VGND VGND VPWR VPWR _04082_ sky130_fd_sc_hd__o21a_1
X_21433_ _01444_ _01445_ _01400_ VGND VGND VPWR VPWR _01446_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24152_ net1015 _04013_ VGND VGND VPWR VPWR _04014_ sky130_fd_sc_hd__xnor2_2
Xwire5217 net5218 VGND VGND VPWR VPWR net5217 sky130_fd_sc_hd__clkbuf_1
X_21364_ _01257_ _01258_ _01259_ VGND VGND VPWR VPWR _01378_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5228 net5229 VGND VGND VPWR VPWR net5228 sky130_fd_sc_hd__clkbuf_1
Xwire5239 net5240 VGND VGND VPWR VPWR net5239 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_31_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23103_ net5062 net4683 _02971_ _02972_ VGND VGND VPWR VPWR _02973_ sky130_fd_sc_hd__a31o_1
X_20315_ net6467 _12118_ net6509 VGND VGND VPWR VPWR _12119_ sky130_fd_sc_hd__a21o_1
Xwire4516 net4514 VGND VGND VPWR VPWR net4516 sky130_fd_sc_hd__buf_1
XFILLER_0_13_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4527 net4530 VGND VGND VPWR VPWR net4527 sky130_fd_sc_hd__buf_1
X_24083_ pid_q.curr_error\[6\] VGND VGND VPWR VPWR _03946_ sky130_fd_sc_hd__inv_2
X_21295_ net5455 _01309_ VGND VGND VPWR VPWR _01310_ sky130_fd_sc_hd__xnor2_1
Xwire4538 net4539 VGND VGND VPWR VPWR net4538 sky130_fd_sc_hd__clkbuf_1
Xwire3804 _01174_ VGND VGND VPWR VPWR net3804 sky130_fd_sc_hd__clkbuf_1
Xwire4549 net4540 VGND VGND VPWR VPWR net4549 sky130_fd_sc_hd__buf_1
X_23034_ net4981 net4715 _02902_ _02903_ VGND VGND VPWR VPWR _02904_ sky130_fd_sc_hd__a31o_1
X_20246_ net13 net14 _12054_ VGND VGND VPWR VPWR _12061_ sky130_fd_sc_hd__and3_1
Xwire3815 _00978_ VGND VGND VPWR VPWR net3815 sky130_fd_sc_hd__clkbuf_1
Xwire3826 net3827 VGND VGND VPWR VPWR net3826 sky130_fd_sc_hd__clkbuf_1
Xwire3837 net3838 VGND VGND VPWR VPWR net3837 sky130_fd_sc_hd__clkbuf_1
Xwire3848 _12274_ VGND VGND VPWR VPWR net3848 sky130_fd_sc_hd__buf_1
Xwire3859 net3860 VGND VGND VPWR VPWR net3859 sky130_fd_sc_hd__buf_1
X_20177_ net3200 net3137 net6013 _11489_ VGND VGND VPWR VPWR _12003_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_181_Left_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24985_ _04747_ VGND VGND VPWR VPWR _00772_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_150_Right_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23936_ _03797_ _03799_ VGND VGND VPWR VPWR _03800_ sky130_fd_sc_hd__and2_1
XFILLER_0_168_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length8566 net8568 VGND VGND VPWR VPWR net8566 sky130_fd_sc_hd__buf_1
X_23867_ _03588_ _03612_ _03611_ VGND VGND VPWR VPWR _03732_ sky130_fd_sc_hd__a21oi_2
Xmax_length8577 net8578 VGND VGND VPWR VPWR net8577 sky130_fd_sc_hd__buf_1
Xmax_length7843 net7835 VGND VGND VPWR VPWR net7843 sky130_fd_sc_hd__clkbuf_1
Xmax_length7865 net7866 VGND VGND VPWR VPWR net7865 sky130_fd_sc_hd__buf_1
X_13620_ _05813_ _05818_ _05819_ VGND VGND VPWR VPWR _05890_ sky130_fd_sc_hd__o21ba_1
X_25606_ clknet_leaf_109_clk _00479_ net8345 VGND VGND VPWR VPWR cordic0.slte0.opB\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_22818_ net8896 _02720_ VGND VGND VPWR VPWR _02721_ sky130_fd_sc_hd__and2_1
XFILLER_0_184_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23798_ _03661_ _03571_ _03663_ VGND VGND VPWR VPWR _03664_ sky130_fd_sc_hd__o21a_1
XFILLER_0_104_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13551_ _05748_ _05755_ _05754_ VGND VGND VPWR VPWR _05822_ sky130_fd_sc_hd__a21bo_1
X_25537_ clknet_leaf_33_clk _00417_ net8691 VGND VGND VPWR VPWR pid_q.prev_int\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22749_ _02677_ VGND VGND VPWR VPWR _00606_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_190_Left_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16270_ _08264_ _08261_ net1250 VGND VGND VPWR VPWR _08334_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25468_ clknet_leaf_52_clk _00348_ net8806 VGND VGND VPWR VPWR svm0.tB\[6\] sky130_fd_sc_hd__dfrtp_1
X_13482_ _05749_ _05750_ net1310 VGND VGND VPWR VPWR _05755_ sky130_fd_sc_hd__nand3_1
Xfanout6313 net6316 VGND VGND VPWR VPWR net6313 sky130_fd_sc_hd__clkbuf_2
Xfanout7058 net7062 VGND VGND VPWR VPWR net7058 sky130_fd_sc_hd__clkbuf_1
Xfanout6324 cordic0.vec\[0\]\[2\] VGND VGND VPWR VPWR net6324 sky130_fd_sc_hd__clkbuf_2
X_15221_ _07292_ net1276 VGND VGND VPWR VPWR _07295_ sky130_fd_sc_hd__nand2_1
X_24419_ net4589 net4791 _04230_ VGND VGND VPWR VPWR _04277_ sky130_fd_sc_hd__and3b_1
Xwire7142 net7139 VGND VGND VPWR VPWR net7142 sky130_fd_sc_hd__clkbuf_2
Xwire7153 net7154 VGND VGND VPWR VPWR net7153 sky130_fd_sc_hd__dlymetal6s2s_1
X_25399_ clknet_leaf_70_clk _00282_ net8451 VGND VGND VPWR VPWR matmul0.a\[2\] sky130_fd_sc_hd__dfrtp_1
Xwire7164 net7165 VGND VGND VPWR VPWR net7164 sky130_fd_sc_hd__buf_1
Xfanout5634 net5636 VGND VGND VPWR VPWR net5634 sky130_fd_sc_hd__buf_1
Xwire6430 cordic0.sin\[1\] VGND VGND VPWR VPWR net6430 sky130_fd_sc_hd__clkbuf_1
Xwire7175 net7176 VGND VGND VPWR VPWR net7175 sky130_fd_sc_hd__clkbuf_1
Xmax_cap1659 _03706_ VGND VGND VPWR VPWR net1659 sky130_fd_sc_hd__buf_1
X_15152_ net3512 net3507 net4170 net4165 VGND VGND VPWR VPWR _07226_ sky130_fd_sc_hd__o22a_1
Xwire6441 net6442 VGND VGND VPWR VPWR net6441 sky130_fd_sc_hd__clkbuf_1
Xwire7186 matmul0.b\[4\] VGND VGND VPWR VPWR net7186 sky130_fd_sc_hd__clkbuf_1
Xfanout5645 net5663 VGND VGND VPWR VPWR net5645 sky130_fd_sc_hd__buf_1
XFILLER_0_62_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout4911 net4927 VGND VGND VPWR VPWR net4911 sky130_fd_sc_hd__buf_1
Xwire7197 matmul0.alpha_pass\[15\] VGND VGND VPWR VPWR net7197 sky130_fd_sc_hd__clkbuf_1
X_14103_ _06356_ _06357_ VGND VGND VPWR VPWR _06365_ sky130_fd_sc_hd__or2_1
Xfanout4933 net4945 VGND VGND VPWR VPWR net4933 sky130_fd_sc_hd__buf_1
Xwire6474 cordic0.gm0.iter\[3\] VGND VGND VPWR VPWR net6474 sky130_fd_sc_hd__clkbuf_1
Xfanout5689 net5695 VGND VGND VPWR VPWR net5689 sky130_fd_sc_hd__buf_1
Xwire6485 net6481 VGND VGND VPWR VPWR net6485 sky130_fd_sc_hd__buf_1
XFILLER_0_1_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5740 net5741 VGND VGND VPWR VPWR net5740 sky130_fd_sc_hd__buf_1
X_19960_ net6111 _11789_ _11790_ VGND VGND VPWR VPWR _11791_ sky130_fd_sc_hd__o21ai_1
Xwire6496 net6497 VGND VGND VPWR VPWR net6496 sky130_fd_sc_hd__clkbuf_1
X_15083_ net4105 net4101 VGND VGND VPWR VPWR _07157_ sky130_fd_sc_hd__nor2_1
Xwire5773 pid_d.mult0.b\[9\] VGND VGND VPWR VPWR net5773 sky130_fd_sc_hd__clkbuf_1
X_14034_ _06220_ _06296_ _06297_ VGND VGND VPWR VPWR _06298_ sky130_fd_sc_hd__o21a_1
Xfanout4988 net4999 VGND VGND VPWR VPWR net4988 sky130_fd_sc_hd__clkbuf_1
Xwire5784 net5785 VGND VGND VPWR VPWR net5784 sky130_fd_sc_hd__buf_1
X_18911_ net6876 net6814 VGND VGND VPWR VPWR _10751_ sky130_fd_sc_hd__nor2_1
Xfanout4999 pid_q.mult0.b\[6\] VGND VGND VPWR VPWR net4999 sky130_fd_sc_hd__buf_1
Xmax_length1493 net1494 VGND VGND VPWR VPWR net1493 sky130_fd_sc_hd__clkbuf_1
X_19891_ _11667_ _11720_ net708 VGND VGND VPWR VPWR _11724_ sky130_fd_sc_hd__o21ai_1
X_18842_ _10682_ _10684_ VGND VGND VPWR VPWR _10685_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15985_ net2239 net3499 VGND VGND VPWR VPWR _08053_ sky130_fd_sc_hd__xnor2_2
X_18773_ net9064 net2287 net1450 _10617_ VGND VGND VPWR VPWR _00445_ sky130_fd_sc_hd__a31o_1
X_17724_ net9122 net1457 net1790 net5169 VGND VGND VPWR VPWR _00429_ sky130_fd_sc_hd__a22o_1
X_14936_ net6611 net7427 matmul0.matmul_stage_inst.a\[5\] net6585 VGND VGND VPWR VPWR
+ _07010_ sky130_fd_sc_hd__a22o_1
X_17655_ net3279 svm0.tA\[10\] VGND VGND VPWR VPWR _09535_ sky130_fd_sc_hd__nand2_1
X_14867_ _06951_ VGND VGND VPWR VPWR _00204_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13818_ net283 _06085_ VGND VGND VPWR VPWR _06086_ sky130_fd_sc_hd__xnor2_1
X_16606_ matmul0.matmul_stage_inst.mult2\[10\] net247 net3471 VGND VGND VPWR VPWR
+ _08653_ sky130_fd_sc_hd__mux2_1
X_17586_ svm0.tC\[15\] _09422_ net4031 VGND VGND VPWR VPWR _09468_ sky130_fd_sc_hd__a21o_1
X_14798_ net7445 matmul0.cos\[3\] net3697 VGND VGND VPWR VPWR _06916_ sky130_fd_sc_hd__and3_1
X_19325_ net6263 _11161_ VGND VGND VPWR VPWR _11162_ sky130_fd_sc_hd__nand2_1
X_16537_ net976 net879 net880 VGND VGND VPWR VPWR _08596_ sky130_fd_sc_hd__o21ba_1
X_13749_ net404 _06003_ VGND VGND VPWR VPWR _06017_ sky130_fd_sc_hd__or2_1
XFILLER_0_156_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19256_ net1422 _11069_ VGND VGND VPWR VPWR _11093_ sky130_fd_sc_hd__nand2_1
X_16468_ _08527_ _08526_ VGND VGND VPWR VPWR _08529_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15419_ _07492_ VGND VGND VPWR VPWR _07493_ sky130_fd_sc_hd__inv_2
X_18207_ net3956 _09676_ _09796_ VGND VGND VPWR VPWR _10058_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_72_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19187_ net6259 net6315 VGND VGND VPWR VPWR _11024_ sky130_fd_sc_hd__or2b_1
X_16399_ net2772 net2204 _08387_ _08460_ VGND VGND VPWR VPWR _08461_ sky130_fd_sc_hd__o31a_1
XFILLER_0_53_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18138_ _09930_ _09987_ VGND VGND VPWR VPWR _09989_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold103 svm0.vC\[10\] VGND VGND VPWR VPWR net9056 sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 pid_q.prev_error\[14\] VGND VGND VPWR VPWR net9067 sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 pid_q.target\[10\] VGND VGND VPWR VPWR net9078 sky130_fd_sc_hd__dlygate4sd3_1
X_18069_ _09902_ _09919_ VGND VGND VPWR VPWR _09920_ sky130_fd_sc_hd__xor2_1
Xhold136 svm0.tA\[0\] VGND VGND VPWR VPWR net9089 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 svm0.tA\[8\] VGND VGND VPWR VPWR net9100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 svm0.tA\[14\] VGND VGND VPWR VPWR net9111 sky130_fd_sc_hd__dlygate4sd3_1
X_20100_ _11909_ VGND VGND VPWR VPWR _11928_ sky130_fd_sc_hd__inv_2
XFILLER_0_186_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold169 pid_q.prev_int\[15\] VGND VGND VPWR VPWR net9122 sky130_fd_sc_hd__dlygate4sd3_1
X_21080_ net5556 _01068_ _01095_ VGND VGND VPWR VPWR _01096_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_112_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20031_ net6112 net6057 VGND VGND VPWR VPWR _11861_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_186_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1709 _02154_ VGND VGND VPWR VPWR net1709 sky130_fd_sc_hd__clkbuf_1
X_24770_ _04596_ _04593_ VGND VGND VPWR VPWR _04598_ sky130_fd_sc_hd__nand2_1
X_21982_ net2477 net1046 VGND VGND VPWR VPWR _01990_ sky130_fd_sc_hd__nor2_1
X_23721_ _03518_ _03522_ _03516_ VGND VGND VPWR VPWR _03587_ sky130_fd_sc_hd__o21ba_1
X_20933_ net5621 net5821 _00947_ _00948_ VGND VGND VPWR VPWR _00949_ sky130_fd_sc_hd__a31o_1
XFILLER_0_178_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23652_ net5154 net5120 VGND VGND VPWR VPWR _03519_ sky130_fd_sc_hd__xor2_1
XFILLER_0_166_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20864_ _12539_ _00879_ VGND VGND VPWR VPWR _00880_ sky130_fd_sc_hd__xnor2_1
X_22603_ _02576_ _02577_ VGND VGND VPWR VPWR _02578_ sky130_fd_sc_hd__and2_1
XFILLER_0_152_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23583_ _03349_ _03368_ _03450_ VGND VGND VPWR VPWR _03451_ sky130_fd_sc_hd__a21o_1
XFILLER_0_165_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20795_ net5627 net5740 VGND VGND VPWR VPWR _00811_ sky130_fd_sc_hd__nand2_1
Xmax_length5759 net5760 VGND VGND VPWR VPWR net5759 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_187_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25322_ clknet_leaf_75_clk _00205_ net8467 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.f\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22534_ net9138 net1700 _02529_ VGND VGND VPWR VPWR _00539_ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25253_ clknet_leaf_88_clk _00136_ net8431 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.a\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_22465_ pid_d.prev_int\[14\] _02397_ _02465_ VGND VGND VPWR VPWR _02466_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24204_ _04061_ _04064_ VGND VGND VPWR VPWR _04065_ sky130_fd_sc_hd__xnor2_1
X_21416_ _01428_ _01429_ VGND VGND VPWR VPWR _01430_ sky130_fd_sc_hd__and2_1
Xwire5003 net5004 VGND VGND VPWR VPWR net5003 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25184_ clknet_leaf_72_clk _00073_ net8470 VGND VGND VPWR VPWR matmul0.a_in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire5014 net5019 VGND VGND VPWR VPWR net5014 sky130_fd_sc_hd__clkbuf_1
X_22396_ pid_d.curr_int\[14\] pid_d.prev_int\[14\] VGND VGND VPWR VPWR _02398_ sky130_fd_sc_hd__xor2_1
Xwire5025 net5026 VGND VGND VPWR VPWR net5025 sky130_fd_sc_hd__buf_1
X_24135_ _03897_ _03906_ _03907_ VGND VGND VPWR VPWR _03997_ sky130_fd_sc_hd__a21bo_1
Xwire4302 net4303 VGND VGND VPWR VPWR net4302 sky130_fd_sc_hd__buf_1
Xwire5047 net5048 VGND VGND VPWR VPWR net5047 sky130_fd_sc_hd__clkbuf_1
X_21347_ net5758 net5543 VGND VGND VPWR VPWR _01361_ sky130_fd_sc_hd__nand2_1
Xwire5058 net5059 VGND VGND VPWR VPWR net5058 sky130_fd_sc_hd__clkbuf_1
Xwire4313 _04861_ VGND VGND VPWR VPWR net4313 sky130_fd_sc_hd__clkbuf_1
Xwire5069 net5070 VGND VGND VPWR VPWR net5069 sky130_fd_sc_hd__buf_1
Xwire4346 net4351 VGND VGND VPWR VPWR net4346 sky130_fd_sc_hd__buf_1
Xwire3601 _06967_ VGND VGND VPWR VPWR net3601 sky130_fd_sc_hd__buf_1
XFILLER_0_102_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24066_ _03927_ _03928_ VGND VGND VPWR VPWR _03929_ sky130_fd_sc_hd__xor2_1
Xwire4357 net4358 VGND VGND VPWR VPWR net4357 sky130_fd_sc_hd__buf_1
X_21278_ net5741 net5590 VGND VGND VPWR VPWR _01293_ sky130_fd_sc_hd__nand2_1
Xwire3634 _06609_ VGND VGND VPWR VPWR net3634 sky130_fd_sc_hd__buf_1
X_23017_ _02880_ _02885_ VGND VGND VPWR VPWR _02887_ sky130_fd_sc_hd__nor2_1
Xwire2900 _06525_ VGND VGND VPWR VPWR net2900 sky130_fd_sc_hd__buf_1
Xwire3645 net3646 VGND VGND VPWR VPWR net3645 sky130_fd_sc_hd__buf_1
Xwire2911 net2912 VGND VGND VPWR VPWR net2911 sky130_fd_sc_hd__clkbuf_1
Xwire3656 net3666 VGND VGND VPWR VPWR net3656 sky130_fd_sc_hd__clkbuf_1
X_20229_ net11 _12047_ VGND VGND VPWR VPWR _12048_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2933 net2934 VGND VGND VPWR VPWR net2933 sky130_fd_sc_hd__clkbuf_1
Xwire3678 net3679 VGND VGND VPWR VPWR net3678 sky130_fd_sc_hd__buf_1
Xwire2944 net2945 VGND VGND VPWR VPWR net2944 sky130_fd_sc_hd__buf_1
Xwire3689 net3690 VGND VGND VPWR VPWR net3689 sky130_fd_sc_hd__buf_1
Xwire2955 _05346_ VGND VGND VPWR VPWR net2955 sky130_fd_sc_hd__buf_1
Xwire2966 _05128_ VGND VGND VPWR VPWR net2966 sky130_fd_sc_hd__buf_1
Xwire2977 net2978 VGND VGND VPWR VPWR net2977 sky130_fd_sc_hd__clkbuf_1
Xwire2988 _04909_ VGND VGND VPWR VPWR net2988 sky130_fd_sc_hd__clkbuf_1
Xwire2999 _00003_ VGND VGND VPWR VPWR net2999 sky130_fd_sc_hd__clkbuf_1
X_15770_ net2234 _07838_ _07839_ VGND VGND VPWR VPWR _07840_ sky130_fd_sc_hd__a21oi_1
X_24968_ pid_q.kp\[3\] _04708_ net1359 VGND VGND VPWR VPWR _04739_ sky130_fd_sc_hd__mux2_1
X_12982_ _05171_ _05172_ _05254_ VGND VGND VPWR VPWR _05255_ sky130_fd_sc_hd__a21o_1
XFILLER_0_188_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length8341 net8342 VGND VGND VPWR VPWR net8341 sky130_fd_sc_hd__buf_1
X_14721_ _06859_ _06860_ net7441 net2876 VGND VGND VPWR VPWR _06861_ sky130_fd_sc_hd__o211a_1
X_23919_ net4572 net4915 VGND VGND VPWR VPWR _03783_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24899_ _04690_ net4507 net2399 VGND VGND VPWR VPWR _04691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17440_ net4251 _09336_ net3386 VGND VGND VPWR VPWR _09337_ sky130_fd_sc_hd__a21o_1
X_14652_ net8958 _06801_ _06810_ VGND VGND VPWR VPWR _00130_ sky130_fd_sc_hd__a21o_1
Xmax_length7662 net7663 VGND VGND VPWR VPWR net7662 sky130_fd_sc_hd__buf_1
Xmax_length7673 net7674 VGND VGND VPWR VPWR net7673 sky130_fd_sc_hd__clkbuf_1
X_13603_ net1589 VGND VGND VPWR VPWR _05873_ sky130_fd_sc_hd__buf_1
XFILLER_0_129_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length6950 net6951 VGND VGND VPWR VPWR net6950 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17371_ net667 VGND VGND VPWR VPWR _09282_ sky130_fd_sc_hd__buf_1
Xmax_length7695 net7696 VGND VGND VPWR VPWR net7695 sky130_fd_sc_hd__clkbuf_1
X_14583_ net2390 _06754_ _06752_ VGND VGND VPWR VPWR _06758_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19110_ _10946_ _10849_ net6181 net6205 VGND VGND VPWR VPWR _10947_ sky130_fd_sc_hd__o2bb2a_1
Xmax_length6994 net6995 VGND VGND VPWR VPWR net6994 sky130_fd_sc_hd__clkbuf_1
X_16322_ net2841 _08382_ _08384_ VGND VGND VPWR VPWR _08385_ sky130_fd_sc_hd__a21oi_1
X_13534_ _05803_ _05804_ VGND VGND VPWR VPWR _05805_ sky130_fd_sc_hd__nand2_1
XFILLER_0_193_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19041_ net6298 net6266 VGND VGND VPWR VPWR _10878_ sky130_fd_sc_hd__nor2b_1
XFILLER_0_40_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16253_ net1509 net1083 VGND VGND VPWR VPWR _08317_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_164_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13465_ _05592_ _05593_ net7769 net1313 VGND VGND VPWR VPWR _05738_ sky130_fd_sc_hd__o211a_1
Xfanout6132 net6146 VGND VGND VPWR VPWR net6132 sky130_fd_sc_hd__buf_1
XFILLER_0_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15204_ net1882 net1544 VGND VGND VPWR VPWR _07278_ sky130_fd_sc_hd__or2b_1
XFILLER_0_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16184_ net1089 net983 _08248_ VGND VGND VPWR VPWR _08249_ sky130_fd_sc_hd__o21a_1
X_13396_ net583 _05668_ net581 VGND VGND VPWR VPWR _05669_ sky130_fd_sc_hd__or3_1
Xfanout5453 net5467 VGND VGND VPWR VPWR net5453 sky130_fd_sc_hd__clkbuf_1
Xwire6260 net6258 VGND VGND VPWR VPWR net6260 sky130_fd_sc_hd__buf_1
XFILLER_0_140_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6271 net6274 VGND VGND VPWR VPWR net6271 sky130_fd_sc_hd__buf_2
XFILLER_0_26_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15135_ _07206_ _07208_ VGND VGND VPWR VPWR _07209_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout4741 net4747 VGND VGND VPWR VPWR net4741 sky130_fd_sc_hd__buf_1
Xwire6282 net6283 VGND VGND VPWR VPWR net6282 sky130_fd_sc_hd__buf_1
Xwire6293 net6291 VGND VGND VPWR VPWR net6293 sky130_fd_sc_hd__buf_1
XFILLER_0_26_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5570 net5571 VGND VGND VPWR VPWR net5570 sky130_fd_sc_hd__buf_1
XFILLER_0_65_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5581 net5584 VGND VGND VPWR VPWR net5581 sky130_fd_sc_hd__buf_1
X_15066_ _07139_ VGND VGND VPWR VPWR _07140_ sky130_fd_sc_hd__buf_1
X_19943_ _11698_ _11703_ _11677_ VGND VGND VPWR VPWR _11775_ sky130_fd_sc_hd__a21bo_1
Xwire5592 net5593 VGND VGND VPWR VPWR net5592 sky130_fd_sc_hd__buf_1
X_14017_ _06246_ _06247_ _06256_ _06249_ VGND VGND VPWR VPWR _06281_ sky130_fd_sc_hd__a31o_1
Xwire4880 net4881 VGND VGND VPWR VPWR net4880 sky130_fd_sc_hd__buf_1
Xwire4891 net4892 VGND VGND VPWR VPWR net4891 sky130_fd_sc_hd__clkbuf_1
X_19874_ net6016 net6033 _11706_ VGND VGND VPWR VPWR _11707_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18825_ _10638_ _10667_ VGND VGND VPWR VPWR _10668_ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18756_ _10558_ _10569_ _10600_ VGND VGND VPWR VPWR _10601_ sky130_fd_sc_hd__o21ai_1
X_15968_ _08034_ net1261 VGND VGND VPWR VPWR _08036_ sky130_fd_sc_hd__xor2_1
XFILLER_0_65_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17707_ _09582_ VGND VGND VPWR VPWR _09583_ sky130_fd_sc_hd__clkbuf_1
X_14919_ net6556 net6587 matmul0.matmul_stage_inst.e\[5\] VGND VGND VPWR VPWR _06993_
+ sky130_fd_sc_hd__o21a_1
X_15899_ net2647 net2748 _07872_ VGND VGND VPWR VPWR _07968_ sky130_fd_sc_hd__o21ai_1
X_18687_ net6796 _10532_ VGND VGND VPWR VPWR _10533_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_81_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17638_ net2153 net1792 _09493_ net2151 _09518_ VGND VGND VPWR VPWR _09519_ sky130_fd_sc_hd__a41o_1
XFILLER_0_187_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17569_ net6734 VGND VGND VPWR VPWR _09451_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19308_ _11140_ _11144_ VGND VGND VPWR VPWR _11145_ sky130_fd_sc_hd__xor2_1
XFILLER_0_144_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20580_ net3325 net3846 _12351_ VGND VGND VPWR VPWR _12363_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length3609 _06939_ VGND VGND VPWR VPWR net3609 sky130_fd_sc_hd__buf_1
XFILLER_0_74_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19239_ net6222 net6323 VGND VGND VPWR VPWR _11076_ sky130_fd_sc_hd__or2b_1
XFILLER_0_33_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22250_ _02254_ _02176_ pid_d.prev_error\[10\] VGND VGND VPWR VPWR _02255_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_121_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21201_ _01065_ _01074_ VGND VGND VPWR VPWR _01217_ sky130_fd_sc_hd__xnor2_1
X_22181_ pid_d.curr_int\[11\] pid_d.prev_int\[11\] VGND VGND VPWR VPWR _02186_ sky130_fd_sc_hd__xor2_1
XFILLER_0_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21132_ _01130_ _01132_ VGND VGND VPWR VPWR _01148_ sky130_fd_sc_hd__xor2_1
X_25940_ clknet_leaf_25_clk _00005_ net8581 VGND VGND VPWR VPWR pid_d.state\[4\] sky130_fd_sc_hd__dfrtp_1
X_21063_ net5581 net5911 VGND VGND VPWR VPWR _01079_ sky130_fd_sc_hd__nand2_1
Xwire2207 _08051_ VGND VGND VPWR VPWR net2207 sky130_fd_sc_hd__clkbuf_1
Xwire2229 net2230 VGND VGND VPWR VPWR net2229 sky130_fd_sc_hd__clkbuf_2
X_20014_ _11841_ _11843_ VGND VGND VPWR VPWR _11844_ sky130_fd_sc_hd__nand2_1
Xwire1506 _08905_ VGND VGND VPWR VPWR net1506 sky130_fd_sc_hd__buf_1
X_25871_ clknet_leaf_18_clk _00744_ net8630 VGND VGND VPWR VPWR pid_q.mult0.a\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1517 _08070_ VGND VGND VPWR VPWR net1517 sky130_fd_sc_hd__buf_1
Xwire1539 net1540 VGND VGND VPWR VPWR net1539 sky130_fd_sc_hd__clkbuf_2
X_24822_ _03313_ _04533_ VGND VGND VPWR VPWR _04644_ sky130_fd_sc_hd__or2_1
X_24753_ net7996 net2009 VGND VGND VPWR VPWR _04584_ sky130_fd_sc_hd__xor2_1
X_21965_ net1045 _01972_ VGND VGND VPWR VPWR _01973_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_90_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23704_ _03568_ _03570_ VGND VGND VPWR VPWR _03571_ sky130_fd_sc_hd__and2_1
X_20916_ _00921_ _00924_ _00916_ VGND VGND VPWR VPWR _00932_ sky130_fd_sc_hd__o21ba_1
X_24684_ net9179 _04507_ _04524_ VGND VGND VPWR VPWR _00694_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21896_ _01742_ _01802_ _01904_ VGND VGND VPWR VPWR _01905_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_65_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23635_ _03496_ net2413 VGND VGND VPWR VPWR _03502_ sky130_fd_sc_hd__xor2_1
X_20847_ _12514_ _12515_ _12516_ VGND VGND VPWR VPWR _00863_ sky130_fd_sc_hd__o21a_1
XFILLER_0_182_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23566_ net4727 net4845 VGND VGND VPWR VPWR _03434_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20778_ net5577 net5774 VGND VGND VPWR VPWR _12549_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25305_ clknet_leaf_69_clk _00188_ net8451 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.e\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire803 _01823_ VGND VGND VPWR VPWR net803 sky130_fd_sc_hd__clkbuf_1
X_22517_ net9195 _12499_ net2489 _02468_ _02517_ VGND VGND VPWR VPWR _00534_ sky130_fd_sc_hd__a221o_1
Xwire814 _10415_ VGND VGND VPWR VPWR net814 sky130_fd_sc_hd__buf_1
Xwire825 _08702_ VGND VGND VPWR VPWR net825 sky130_fd_sc_hd__clkbuf_1
X_23497_ _03289_ _03291_ _03365_ VGND VGND VPWR VPWR _03366_ sky130_fd_sc_hd__o21a_1
Xwire836 _06184_ VGND VGND VPWR VPWR net836 sky130_fd_sc_hd__buf_1
XFILLER_0_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire847 _05503_ VGND VGND VPWR VPWR net847 sky130_fd_sc_hd__buf_1
XFILLER_0_51_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13250_ _05520_ _05522_ VGND VGND VPWR VPWR _05523_ sky130_fd_sc_hd__xor2_1
X_25236_ clknet_leaf_23_clk _00009_ net8582 VGND VGND VPWR VPWR pid_q.state\[3\] sky130_fd_sc_hd__dfrtp_1
Xwire858 _02592_ VGND VGND VPWR VPWR net858 sky130_fd_sc_hd__buf_1
X_22448_ _02417_ _02449_ VGND VGND VPWR VPWR _02450_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire869 net870 VGND VGND VPWR VPWR net869 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13181_ _05450_ _05453_ VGND VGND VPWR VPWR _05454_ sky130_fd_sc_hd__xnor2_1
X_25167_ clknet_leaf_55_clk _00056_ net8728 VGND VGND VPWR VPWR svm0.periodTop\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_22379_ _02313_ _02316_ _02381_ VGND VGND VPWR VPWR _02382_ sky130_fd_sc_hd__a21o_1
Xwire4110 _07127_ VGND VGND VPWR VPWR net4110 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4121 net4122 VGND VGND VPWR VPWR net4121 sky130_fd_sc_hd__buf_1
X_24118_ net4604 net4835 VGND VGND VPWR VPWR _03980_ sky130_fd_sc_hd__nand2_1
Xwire4132 net4133 VGND VGND VPWR VPWR net4132 sky130_fd_sc_hd__buf_1
XFILLER_0_130_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25098_ net1627 _04840_ _04841_ net2148 VGND VGND VPWR VPWR _04842_ sky130_fd_sc_hd__a211o_1
Xwire4143 net4144 VGND VGND VPWR VPWR net4143 sky130_fd_sc_hd__clkbuf_2
Xwire4154 net4155 VGND VGND VPWR VPWR net4154 sky130_fd_sc_hd__buf_1
Xwire4165 net4166 VGND VGND VPWR VPWR net4165 sky130_fd_sc_hd__buf_1
Xwire3420 net3421 VGND VGND VPWR VPWR net3420 sky130_fd_sc_hd__buf_1
XFILLER_0_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3431 net3432 VGND VGND VPWR VPWR net3431 sky130_fd_sc_hd__buf_1
Xwire4176 net4177 VGND VGND VPWR VPWR net4176 sky130_fd_sc_hd__buf_1
X_24049_ _03788_ _03793_ net2411 VGND VGND VPWR VPWR _03912_ sky130_fd_sc_hd__o21a_1
X_16940_ _08856_ _08860_ net2176 net2174 _08903_ VGND VGND VPWR VPWR _08904_ sky130_fd_sc_hd__o221a_1
Xwire3442 _07353_ VGND VGND VPWR VPWR net3442 sky130_fd_sc_hd__buf_1
XFILLER_0_159_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4187 net4188 VGND VGND VPWR VPWR net4187 sky130_fd_sc_hd__buf_1
XFILLER_0_25_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4198 net4199 VGND VGND VPWR VPWR net4198 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3453 _07194_ VGND VGND VPWR VPWR net3453 sky130_fd_sc_hd__buf_1
Xwire3464 _07179_ VGND VGND VPWR VPWR net3464 sky130_fd_sc_hd__buf_1
Xwire2730 _07240_ VGND VGND VPWR VPWR net2730 sky130_fd_sc_hd__buf_1
Xwire3475 net3476 VGND VGND VPWR VPWR net3475 sky130_fd_sc_hd__buf_1
Xwire2741 net2742 VGND VGND VPWR VPWR net2741 sky130_fd_sc_hd__clkbuf_1
Xwire3486 net3487 VGND VGND VPWR VPWR net3486 sky130_fd_sc_hd__buf_1
X_16871_ net6468 _08835_ VGND VGND VPWR VPWR _08836_ sky130_fd_sc_hd__nor2_2
Xwire3497 net3498 VGND VGND VPWR VPWR net3497 sky130_fd_sc_hd__buf_1
Xwire2752 net2753 VGND VGND VPWR VPWR net2752 sky130_fd_sc_hd__buf_1
Xwire2774 net2775 VGND VGND VPWR VPWR net2774 sky130_fd_sc_hd__clkbuf_1
X_18610_ net714 _10457_ VGND VGND VPWR VPWR _10458_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_189_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15822_ _07775_ _07798_ _07891_ VGND VGND VPWR VPWR _07892_ sky130_fd_sc_hd__a21o_1
Xwire2785 net2786 VGND VGND VPWR VPWR net2785 sky130_fd_sc_hd__clkbuf_1
X_19590_ _11375_ _11417_ VGND VGND VPWR VPWR _11427_ sky130_fd_sc_hd__nor2_1
Xwire2796 net2797 VGND VGND VPWR VPWR net2796 sky130_fd_sc_hd__buf_1
XFILLER_0_95_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15753_ _07645_ _07734_ VGND VGND VPWR VPWR _07824_ sky130_fd_sc_hd__nor2_1
X_18541_ _10387_ _10309_ net2587 VGND VGND VPWR VPWR _10390_ sky130_fd_sc_hd__a21oi_1
X_12965_ _05024_ _05020_ _05030_ VGND VGND VPWR VPWR _05238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14704_ net7459 _06847_ VGND VGND VPWR VPWR _06848_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15684_ _07753_ _07754_ VGND VGND VPWR VPWR _07755_ sky130_fd_sc_hd__xnor2_1
X_18472_ net3930 _10317_ _10320_ _10321_ VGND VGND VPWR VPWR _10322_ sky130_fd_sc_hd__o211a_1
X_12896_ _05153_ _05154_ _05166_ _05167_ VGND VGND VPWR VPWR _05169_ sky130_fd_sc_hd__or4_2
XFILLER_0_185_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17423_ net9162 _09323_ VGND VGND VPWR VPWR _09324_ sky130_fd_sc_hd__xnor2_1
X_14635_ net4282 VGND VGND VPWR VPWR _06800_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17354_ net1465 _09267_ VGND VGND VPWR VPWR _00375_ sky130_fd_sc_hd__nand2_1
X_14566_ net1625 _06742_ _06730_ VGND VGND VPWR VPWR _06743_ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13517_ _05786_ _05787_ VGND VGND VPWR VPWR _05788_ sky130_fd_sc_hd__xor2_1
X_16305_ _08363_ _08368_ VGND VGND VPWR VPWR _08369_ sky130_fd_sc_hd__or2_1
X_17285_ _09198_ _09199_ VGND VGND VPWR VPWR _09200_ sky130_fd_sc_hd__or2_1
X_14497_ net7324 net5278 VGND VGND VPWR VPWR _06680_ sky130_fd_sc_hd__nor2_1
X_19024_ _10809_ _10835_ _10860_ VGND VGND VPWR VPWR _10861_ sky130_fd_sc_hd__a21o_1
X_16236_ _08245_ _08300_ VGND VGND VPWR VPWR _08301_ sky130_fd_sc_hd__xnor2_1
X_13448_ _05719_ _05720_ _05621_ _05622_ VGND VGND VPWR VPWR _05721_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16167_ _08150_ _08155_ _08232_ VGND VGND VPWR VPWR _08233_ sky130_fd_sc_hd__o21ai_2
X_13379_ net628 _05651_ VGND VGND VPWR VPWR _05652_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6090 cordic0.vec\[0\]\[13\] VGND VGND VPWR VPWR net6090 sky130_fd_sc_hd__buf_1
X_15118_ net4175 net4173 VGND VGND VPWR VPWR _07192_ sky130_fd_sc_hd__nor2_1
X_16098_ _07841_ net1260 VGND VGND VPWR VPWR _08164_ sky130_fd_sc_hd__and2b_1
XFILLER_0_76_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19926_ net6168 net6081 VGND VGND VPWR VPWR _11758_ sky130_fd_sc_hd__xnor2_2
X_15049_ _07075_ net1285 net1283 VGND VGND VPWR VPWR _07123_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_167_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19857_ net6169 net6098 VGND VGND VPWR VPWR _11690_ sky130_fd_sc_hd__xnor2_2
X_18808_ _10627_ _10651_ VGND VGND VPWR VPWR _10652_ sky130_fd_sc_hd__xnor2_1
X_19788_ _11584_ _11592_ _11580_ VGND VGND VPWR VPWR _11622_ sky130_fd_sc_hd__o21a_1
X_18739_ _10582_ _10583_ VGND VGND VPWR VPWR _10584_ sky130_fd_sc_hd__nor2_1
XFILLER_0_183_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_188_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21750_ _01756_ _01759_ VGND VGND VPWR VPWR _01760_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_25_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20701_ _12473_ _12474_ VGND VGND VPWR VPWR _12475_ sky130_fd_sc_hd__xor2_2
X_21681_ net5813 net5440 VGND VGND VPWR VPWR _01692_ sky130_fd_sc_hd__nand2_1
XFILLER_0_164_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_191_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23420_ _03208_ _03209_ _03210_ VGND VGND VPWR VPWR _03290_ sky130_fd_sc_hd__o21a_1
X_20632_ _12410_ _12406_ VGND VGND VPWR VPWR _12412_ sky130_fd_sc_hd__or2b_1
XFILLER_0_50_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7708 net7709 VGND VGND VPWR VPWR net7708 sky130_fd_sc_hd__buf_1
XFILLER_0_135_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7719 net7720 VGND VGND VPWR VPWR net7719 sky130_fd_sc_hd__buf_1
XFILLER_0_18_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23351_ _03217_ _03220_ VGND VGND VPWR VPWR _03221_ sky130_fd_sc_hd__xnor2_2
X_20563_ net8057 net2516 _12346_ _12347_ VGND VGND VPWR VPWR _00505_ sky130_fd_sc_hd__a31o_1
XFILLER_0_61_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3439 net3440 VGND VGND VPWR VPWR net3439 sky130_fd_sc_hd__buf_1
X_22302_ net5762 net3786 _02228_ VGND VGND VPWR VPWR _02306_ sky130_fd_sc_hd__nand3_1
XFILLER_0_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23282_ net4912 net4775 VGND VGND VPWR VPWR _03152_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20494_ net2088 VGND VGND VPWR VPWR _12282_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25021_ net4457 pid_q.curr_int\[4\] VGND VGND VPWR VPWR _04775_ sky130_fd_sc_hd__xnor2_1
X_22233_ _02152_ _02155_ net1712 VGND VGND VPWR VPWR _02238_ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22164_ _02116_ _02168_ VGND VGND VPWR VPWR _02170_ sky130_fd_sc_hd__or2_1
X_21115_ _01086_ _01083_ VGND VGND VPWR VPWR _01131_ sky130_fd_sc_hd__xnor2_1
Xwire2004 net2005 VGND VGND VPWR VPWR net2004 sky130_fd_sc_hd__clkbuf_1
X_22095_ _02100_ _02010_ _02101_ VGND VGND VPWR VPWR _02102_ sky130_fd_sc_hd__a21o_1
Xwire2015 _04535_ VGND VGND VPWR VPWR net2015 sky130_fd_sc_hd__buf_1
Xwire2026 _02930_ VGND VGND VPWR VPWR net2026 sky130_fd_sc_hd__buf_1
Xwire2037 net2039 VGND VGND VPWR VPWR net2037 sky130_fd_sc_hd__buf_1
X_25923_ clknet_leaf_96_clk _00796_ net8402 VGND VGND VPWR VPWR pid_d.prev_int\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_100_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21046_ net2075 net2074 net2480 VGND VGND VPWR VPWR _01062_ sky130_fd_sc_hd__and3_1
Xwire2048 _02524_ VGND VGND VPWR VPWR net2048 sky130_fd_sc_hd__buf_1
Xwire1314 net1315 VGND VGND VPWR VPWR net1314 sky130_fd_sc_hd__buf_1
Xwire2059 _01894_ VGND VGND VPWR VPWR net2059 sky130_fd_sc_hd__buf_1
Xwire1325 net1326 VGND VGND VPWR VPWR net1325 sky130_fd_sc_hd__clkbuf_1
Xwire1336 _05098_ VGND VGND VPWR VPWR net1336 sky130_fd_sc_hd__clkbuf_2
Xwire1347 net1348 VGND VGND VPWR VPWR net1347 sky130_fd_sc_hd__clkbuf_1
X_25854_ clknet_leaf_23_clk _00727_ net8586 VGND VGND VPWR VPWR pid_q.mult0.b\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1358 net1359 VGND VGND VPWR VPWR net1358 sky130_fd_sc_hd__clkbuf_2
X_24805_ net5194 net2385 VGND VGND VPWR VPWR _04629_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25785_ clknet_leaf_57_clk _00658_ net8716 VGND VGND VPWR VPWR matmul0.beta_pass\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_22997_ _02866_ VGND VGND VPWR VPWR _02867_ sky130_fd_sc_hd__buf_1
XFILLER_0_9_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24736_ _04567_ _04568_ VGND VGND VPWR VPWR _04569_ sky130_fd_sc_hd__xnor2_1
X_12750_ net1608 net1342 net3689 VGND VGND VPWR VPWR _05023_ sky130_fd_sc_hd__and3_1
X_21948_ _01783_ _01955_ _01781_ VGND VGND VPWR VPWR _01956_ sky130_fd_sc_hd__a21oi_1
X_24667_ pid_q.curr_error\[5\] net2383 net1373 VGND VGND VPWR VPWR _04516_ sky130_fd_sc_hd__and3_1
X_12681_ _04945_ net1008 _04953_ VGND VGND VPWR VPWR _04954_ sky130_fd_sc_hd__o21a_1
XFILLER_0_167_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21879_ _01887_ _01788_ VGND VGND VPWR VPWR _01888_ sky130_fd_sc_hd__nand2_1
Xmax_length6054 net6057 VGND VGND VPWR VPWR net6054 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14420_ net8132 net3631 VGND VGND VPWR VPWR _06619_ sky130_fd_sc_hd__and2_1
X_23618_ _03483_ _03484_ VGND VGND VPWR VPWR _03485_ sky130_fd_sc_hd__xnor2_1
Xwire8910 net8911 VGND VGND VPWR VPWR net8910 sky130_fd_sc_hd__clkbuf_1
Xwire8921 net8922 VGND VGND VPWR VPWR net8921 sky130_fd_sc_hd__buf_1
XFILLER_0_166_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24598_ net7522 _04392_ net234 net7465 net230 VGND VGND VPWR VPWR _04454_ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8932 net8933 VGND VGND VPWR VPWR net8932 sky130_fd_sc_hd__clkbuf_1
Xwire8943 net8944 VGND VGND VPWR VPWR net8943 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire600 net601 VGND VGND VPWR VPWR net600 sky130_fd_sc_hd__buf_1
X_14351_ _06565_ VGND VGND VPWR VPWR _00074_ sky130_fd_sc_hd__clkbuf_1
X_23549_ _03337_ _03338_ _03416_ VGND VGND VPWR VPWR _03417_ sky130_fd_sc_hd__a21oi_2
Xwire611 net613 VGND VGND VPWR VPWR net611 sky130_fd_sc_hd__buf_1
XFILLER_0_135_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire622 net623 VGND VGND VPWR VPWR net622 sky130_fd_sc_hd__buf_1
XFILLER_0_37_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13302_ _05499_ net1135 VGND VGND VPWR VPWR _05575_ sky130_fd_sc_hd__and2b_1
Xwire633 _04167_ VGND VGND VPWR VPWR net633 sky130_fd_sc_hd__clkbuf_2
Xwire644 net645 VGND VGND VPWR VPWR net644 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17070_ _08946_ _08947_ net2601 VGND VGND VPWR VPWR _09028_ sky130_fd_sc_hd__mux2_1
X_14282_ net73 net2902 net2265 net7880 VGND VGND VPWR VPWR _00053_ sky130_fd_sc_hd__a22o_1
Xwire655 net656 VGND VGND VPWR VPWR net655 sky130_fd_sc_hd__clkbuf_1
Xmax_length3951 _09876_ VGND VGND VPWR VPWR net3951 sky130_fd_sc_hd__clkbuf_1
Xwire666 _10266_ VGND VGND VPWR VPWR net666 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire677 _06204_ VGND VGND VPWR VPWR net677 sky130_fd_sc_hd__buf_1
XFILLER_0_126_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16021_ _08008_ _08082_ VGND VGND VPWR VPWR _08088_ sky130_fd_sc_hd__or2b_1
Xwire688 net689 VGND VGND VPWR VPWR net688 sky130_fd_sc_hd__clkbuf_1
X_13233_ net7780 net3685 net2967 VGND VGND VPWR VPWR _05506_ sky130_fd_sc_hd__and3_1
X_25219_ clknet_leaf_59_clk _00108_ net8688 VGND VGND VPWR VPWR svm0.vC\[7\] sky130_fd_sc_hd__dfrtp_1
Xwire699 _01914_ VGND VGND VPWR VPWR net699 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13164_ _05374_ _05375_ net7757 net1620 VGND VGND VPWR VPWR _05437_ sky130_fd_sc_hd__o211a_1
X_13095_ net7716 net2351 net2347 VGND VGND VPWR VPWR _05368_ sky130_fd_sc_hd__and3_1
X_17972_ _09817_ _09822_ VGND VGND VPWR VPWR _09823_ sky130_fd_sc_hd__xor2_1
Xwire3250 net3251 VGND VGND VPWR VPWR net3250 sky130_fd_sc_hd__clkbuf_1
X_19711_ _11425_ _11481_ _11482_ VGND VGND VPWR VPWR _11547_ sky130_fd_sc_hd__a21o_1
X_16923_ cordic0.slte0.opA\[2\] cordic0.slte0.opA\[1\] cordic0.slte0.opA\[0\] VGND
+ VGND VPWR VPWR _08887_ sky130_fd_sc_hd__or3_1
Xwire3272 _09393_ VGND VGND VPWR VPWR net3272 sky130_fd_sc_hd__buf_1
XFILLER_0_137_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3283 _09177_ VGND VGND VPWR VPWR net3283 sky130_fd_sc_hd__buf_1
Xwire3294 net3295 VGND VGND VPWR VPWR net3294 sky130_fd_sc_hd__buf_1
Xwire2560 _09683_ VGND VGND VPWR VPWR net2560 sky130_fd_sc_hd__clkbuf_1
Xwire2571 _09286_ VGND VGND VPWR VPWR net2571 sky130_fd_sc_hd__buf_1
X_19642_ net1191 _11478_ VGND VGND VPWR VPWR _11479_ sky130_fd_sc_hd__xor2_1
X_16854_ net2196 VGND VGND VPWR VPWR _08819_ sky130_fd_sc_hd__buf_1
Xwire2582 _09170_ VGND VGND VPWR VPWR net2582 sky130_fd_sc_hd__buf_1
X_15805_ _07873_ _07874_ VGND VGND VPWR VPWR _07875_ sky130_fd_sc_hd__xor2_1
Xwire1870 net1871 VGND VGND VPWR VPWR net1870 sky130_fd_sc_hd__clkbuf_1
X_19573_ _10996_ VGND VGND VPWR VPWR _11410_ sky130_fd_sc_hd__buf_1
Xwire1881 _07283_ VGND VGND VPWR VPWR net1881 sky130_fd_sc_hd__buf_1
X_13997_ net7766 net1569 _06169_ VGND VGND VPWR VPWR _06262_ sky130_fd_sc_hd__and3_1
Xwire1892 _07197_ VGND VGND VPWR VPWR net1892 sky130_fd_sc_hd__buf_1
X_16785_ _08782_ VGND VGND VPWR VPWR _00291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18524_ _10371_ _10372_ net3981 VGND VGND VPWR VPWR _10373_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12948_ _05214_ net1593 net1003 VGND VGND VPWR VPWR _05221_ sky130_fd_sc_hd__o21ai_1
X_15736_ net2250 net2672 _07805_ _07806_ _07724_ VGND VGND VPWR VPWR _07807_ sky130_fd_sc_hd__o32a_1
XFILLER_0_87_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18455_ _10301_ _10304_ VGND VGND VPWR VPWR _10305_ sky130_fd_sc_hd__xnor2_1
X_12879_ _05151_ _05144_ VGND VGND VPWR VPWR _05152_ sky130_fd_sc_hd__nor2_1
X_15667_ _07736_ _07738_ VGND VGND VPWR VPWR _07739_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17406_ _09307_ net616 _09308_ _09310_ VGND VGND VPWR VPWR _00384_ sky130_fd_sc_hd__a31o_1
XFILLER_0_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14618_ _06789_ VGND VGND VPWR VPWR _00117_ sky130_fd_sc_hd__clkbuf_1
X_18386_ net3241 _09909_ _09701_ VGND VGND VPWR VPWR _10237_ sky130_fd_sc_hd__or3b_1
X_15598_ net3447 net3537 VGND VGND VPWR VPWR _07670_ sky130_fd_sc_hd__nor2_1
X_17337_ net6698 net7661 VGND VGND VPWR VPWR _09251_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14549_ _06710_ _06725_ _06726_ net5250 VGND VGND VPWR VPWR _06727_ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17268_ net2160 net256 net1797 net9186 VGND VGND VPWR VPWR _00362_ sky130_fd_sc_hd__a22o_1
X_19007_ net3202 net3898 _10800_ VGND VGND VPWR VPWR _10844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16219_ _08193_ _08198_ _08191_ VGND VGND VPWR VPWR _08284_ sky130_fd_sc_hd__a21o_1
XFILLER_0_140_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17199_ net6850 net618 VGND VGND VPWR VPWR _09149_ sky130_fd_sc_hd__nor2_1
XFILLER_0_178_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5091 net5103 VGND VGND VPWR VPWR net5091 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19909_ _11716_ _11737_ _11740_ VGND VGND VPWR VPWR _11741_ sky130_fd_sc_hd__o21ba_1
Xhold18 svm0.tA\[9\] VGND VGND VPWR VPWR net8971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 matmul0.matmul_stage_inst.a\[12\] VGND VGND VPWR VPWR net8982 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_3_Left_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22920_ _02270_ _02802_ _02810_ VGND VGND VPWR VPWR _02811_ sky130_fd_sc_hd__a21o_1
XFILLER_0_194_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22851_ net4360 net475 _02749_ net4336 net2465 VGND VGND VPWR VPWR _02750_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21802_ _01810_ _01730_ _01811_ VGND VGND VPWR VPWR _01812_ sky130_fd_sc_hd__a21o_1
X_25570_ clknet_leaf_97_clk _00443_ net8398 VGND VGND VPWR VPWR cordic0.sin\[4\] sky130_fd_sc_hd__dfrtp_1
X_22782_ pid_d.kp\[3\] _02668_ net1679 VGND VGND VPWR VPWR _02699_ sky130_fd_sc_hd__mux2_1
X_24521_ _04268_ _04376_ _04314_ _04377_ VGND VGND VPWR VPWR _04378_ sky130_fd_sc_hd__o2bb2a_1
X_21733_ net1173 _01706_ net1174 VGND VGND VPWR VPWR _01743_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24452_ _04229_ _04233_ _04234_ VGND VGND VPWR VPWR _04310_ sky130_fd_sc_hd__o21a_1
Xwire8206 net8207 VGND VGND VPWR VPWR net8206 sky130_fd_sc_hd__clkbuf_1
X_21664_ net5798 net5460 VGND VGND VPWR VPWR _01675_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8217 net8218 VGND VGND VPWR VPWR net8217 sky130_fd_sc_hd__clkbuf_1
Xwire8228 net8229 VGND VGND VPWR VPWR net8228 sky130_fd_sc_hd__clkbuf_1
Xwire8239 net8240 VGND VGND VPWR VPWR net8239 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23403_ net5054 net4597 VGND VGND VPWR VPWR _03273_ sky130_fd_sc_hd__nand2_1
Xwire7505 net7506 VGND VGND VPWR VPWR net7505 sky130_fd_sc_hd__buf_1
Xwire7516 net7517 VGND VGND VPWR VPWR net7516 sky130_fd_sc_hd__clkbuf_1
Xmax_length3203 _10843_ VGND VGND VPWR VPWR net3203 sky130_fd_sc_hd__buf_1
X_20615_ net2601 _12394_ _12395_ net3325 _12353_ VGND VGND VPWR VPWR _12396_ sky130_fd_sc_hd__o221a_1
X_24383_ _04153_ _04157_ _04241_ VGND VGND VPWR VPWR _04242_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_49_Left_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire7527 net7525 VGND VGND VPWR VPWR net7527 sky130_fd_sc_hd__buf_1
X_21595_ net5961 net5943 net5921 net3115 VGND VGND VPWR VPWR _01607_ sky130_fd_sc_hd__o211a_1
Xmax_length3225 _10223_ VGND VGND VPWR VPWR net3225 sky130_fd_sc_hd__clkbuf_2
Xwire7538 net7539 VGND VGND VPWR VPWR net7538 sky130_fd_sc_hd__clkbuf_1
Xwire7549 svm0.vC\[9\] VGND VGND VPWR VPWR net7549 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6804 net6806 VGND VGND VPWR VPWR net6804 sky130_fd_sc_hd__buf_1
X_23334_ _03202_ _03203_ VGND VGND VPWR VPWR _03204_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20546_ net1822 net2084 _12329_ VGND VGND VPWR VPWR _12331_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire6837 net6838 VGND VGND VPWR VPWR net6837 sky130_fd_sc_hd__buf_1
XFILLER_0_144_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6848 net6849 VGND VGND VPWR VPWR net6848 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6859 net6858 VGND VGND VPWR VPWR net6859 sky130_fd_sc_hd__buf_1
X_23265_ _03026_ _03033_ _03038_ _03043_ VGND VGND VPWR VPWR _03135_ sky130_fd_sc_hd__a22oi_2
X_20477_ net6962 net6917 net6937 net6904 net6491 net6521 VGND VGND VPWR VPWR _12266_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_120_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25004_ pid_q.out\[1\] net5181 VGND VGND VPWR VPWR _04760_ sky130_fd_sc_hd__or2_1
X_22216_ net2052 _02220_ VGND VGND VPWR VPWR _02221_ sky130_fd_sc_hd__xnor2_2
X_23196_ net5065 net5040 _03065_ VGND VGND VPWR VPWR _03066_ sky130_fd_sc_hd__and3_1
X_22147_ _02045_ _02047_ _02043_ VGND VGND VPWR VPWR _02153_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_30_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22078_ net1717 _01980_ VGND VGND VPWR VPWR _02085_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_58_Left_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1100 net1101 VGND VGND VPWR VPWR net1100 sky130_fd_sc_hd__clkbuf_1
Xwire1111 net1112 VGND VGND VPWR VPWR net1111 sky130_fd_sc_hd__clkbuf_1
Xwire1122 net1123 VGND VGND VPWR VPWR net1122 sky130_fd_sc_hd__buf_1
XFILLER_0_156_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13920_ net7645 net1331 VGND VGND VPWR VPWR _06186_ sky130_fd_sc_hd__nand2_1
X_25906_ clknet_leaf_65_clk _00779_ net8703 VGND VGND VPWR VPWR pid_q.out\[2\] sky130_fd_sc_hd__dfrtp_1
X_21029_ _01043_ _01044_ VGND VGND VPWR VPWR _01045_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_96_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1133 net1134 VGND VGND VPWR VPWR net1133 sky130_fd_sc_hd__buf_1
Xwire1144 net1145 VGND VGND VPWR VPWR net1144 sky130_fd_sc_hd__clkbuf_1
Xwire1155 net1156 VGND VGND VPWR VPWR net1155 sky130_fd_sc_hd__buf_1
XFILLER_0_107_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1166 _03301_ VGND VGND VPWR VPWR net1166 sky130_fd_sc_hd__buf_1
X_13851_ _06117_ net1950 VGND VGND VPWR VPWR _06118_ sky130_fd_sc_hd__nor2_1
X_25837_ clknet_leaf_31_clk _00710_ net8684 VGND VGND VPWR VPWR pid_q.curr_error\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1177 _01584_ VGND VGND VPWR VPWR net1177 sky130_fd_sc_hd__buf_1
XFILLER_0_18_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1188 net1189 VGND VGND VPWR VPWR net1188 sky130_fd_sc_hd__clkbuf_2
X_12802_ net1343 _04969_ VGND VGND VPWR VPWR _05075_ sky130_fd_sc_hd__or2_1
X_13782_ _06042_ _06049_ VGND VGND VPWR VPWR _06050_ sky130_fd_sc_hd__xnor2_2
X_16570_ _08550_ _08554_ _08628_ VGND VGND VPWR VPWR _08629_ sky130_fd_sc_hd__o21a_1
XFILLER_0_186_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25768_ clknet_leaf_27_clk _00641_ net8646 VGND VGND VPWR VPWR pid_d.out\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12733_ net7853 net2338 net1968 VGND VGND VPWR VPWR _05006_ sky130_fd_sc_hd__and3_1
X_15521_ net3447 net3518 VGND VGND VPWR VPWR _07594_ sky130_fd_sc_hd__nor2_1
X_24719_ _04552_ _04553_ VGND VGND VPWR VPWR _04554_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25699_ clknet_leaf_0_clk _00572_ net8409 VGND VGND VPWR VPWR pid_d.mult0.b\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout8623 net8629 VGND VGND VPWR VPWR net8623 sky130_fd_sc_hd__clkbuf_1
X_15452_ net4161 net4157 net4143 net4140 VGND VGND VPWR VPWR _07526_ sky130_fd_sc_hd__o22a_1
X_18240_ _10037_ net2564 _10030_ net3254 VGND VGND VPWR VPWR _10091_ sky130_fd_sc_hd__a211o_1
X_12664_ net7777 net2340 _04932_ VGND VGND VPWR VPWR _04937_ sky130_fd_sc_hd__and3_1
Xfanout8645 net8660 VGND VGND VPWR VPWR net8645 sky130_fd_sc_hd__buf_1
XFILLER_0_127_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_67_Left_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14403_ net994 VGND VGND VPWR VPWR _06606_ sky130_fd_sc_hd__buf_1
Xwire8740 net8741 VGND VGND VPWR VPWR net8740 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15383_ _07455_ _07456_ VGND VGND VPWR VPWR _07457_ sky130_fd_sc_hd__nand2_1
X_18171_ _10020_ _09776_ _10021_ _09841_ VGND VGND VPWR VPWR _10022_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12595_ matmul0.state\[0\] matmul0.start VGND VGND VPWR VPWR _04876_ sky130_fd_sc_hd__nand2_1
Xwire8762 net8760 VGND VGND VPWR VPWR net8762 sky130_fd_sc_hd__clkbuf_2
X_17122_ _09075_ _09077_ VGND VGND VPWR VPWR _09078_ sky130_fd_sc_hd__xnor2_1
Xwire430 net431 VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__clkbuf_1
X_14334_ _06552_ matmul0.a_in\[3\] net902 VGND VGND VPWR VPWR _06553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8795 net8796 VGND VGND VPWR VPWR net8795 sky130_fd_sc_hd__clkbuf_1
Xwire441 net442 VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__clkbuf_1
Xwire452 net453 VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__clkbuf_1
Xwire463 net464 VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__buf_1
XFILLER_0_40_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17053_ net1802 _09011_ VGND VGND VPWR VPWR _09012_ sky130_fd_sc_hd__xor2_2
Xwire474 _01809_ VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__clkbuf_1
X_14265_ net58 _06511_ _06515_ net8985 VGND VGND VPWR VPWR _00038_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire485 net486 VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire496 net497 VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__clkbuf_1
X_16004_ net1521 net1257 VGND VGND VPWR VPWR _08072_ sky130_fd_sc_hd__xnor2_1
X_13216_ net7713 net1606 VGND VGND VPWR VPWR _05489_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_164_Right_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14196_ _06450_ _06455_ VGND VGND VPWR VPWR _06456_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13147_ net5199 net3028 net3693 net2992 svm0.vC\[13\] VGND VGND VPWR VPWR _05420_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_148_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_76_Left_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13078_ _05345_ net4255 VGND VGND VPWR VPWR _05351_ sky130_fd_sc_hd__nand2_1
X_17955_ _09803_ _09804_ net2552 VGND VGND VPWR VPWR _09806_ sky130_fd_sc_hd__o21ai_1
Xwire3080 net3081 VGND VGND VPWR VPWR net3080 sky130_fd_sc_hd__buf_1
X_16906_ net6402 _08865_ _08867_ _08868_ _08869_ VGND VGND VPWR VPWR _08870_ sky130_fd_sc_hd__a221o_1
X_17886_ net3964 _09736_ VGND VGND VPWR VPWR _09737_ sky130_fd_sc_hd__xnor2_1
Xwire2390 _04858_ VGND VGND VPWR VPWR net2390 sky130_fd_sc_hd__buf_1
XFILLER_0_189_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19625_ net3176 _10917_ net3186 VGND VGND VPWR VPWR _11462_ sky130_fd_sc_hd__mux2_1
X_16837_ _08809_ VGND VGND VPWR VPWR _00316_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_178_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19556_ _11076_ _11075_ VGND VGND VPWR VPWR _11393_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16768_ _08773_ VGND VGND VPWR VPWR _00283_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18507_ _10352_ _10353_ _10355_ VGND VGND VPWR VPWR _10356_ sky130_fd_sc_hd__and3_1
X_15719_ net2225 _07789_ VGND VGND VPWR VPWR _07790_ sky130_fd_sc_hd__xnor2_2
X_19487_ _11076_ _11075_ VGND VGND VPWR VPWR _11324_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_85_Left_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16699_ matmul0.matmul_stage_inst.mult1\[11\] VGND VGND VPWR VPWR _08728_ sky130_fd_sc_hd__inv_2
X_18438_ _10284_ _10287_ VGND VGND VPWR VPWR _10288_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18369_ net6858 net6879 VGND VGND VPWR VPWR _10220_ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20400_ cordic0.slte0.opA\[8\] net865 VGND VGND VPWR VPWR _12198_ sky130_fd_sc_hd__or2_1
X_21380_ _01288_ _01289_ _01393_ VGND VGND VPWR VPWR _01394_ sky130_fd_sc_hd__o21a_1
XFILLER_0_154_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20331_ net3667 _12133_ VGND VGND VPWR VPWR _12134_ sky130_fd_sc_hd__or2_1
Xmax_length1119 net1120 VGND VGND VPWR VPWR net1119 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_109_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4709 net4710 VGND VGND VPWR VPWR net4709 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23050_ _02889_ _02908_ _02919_ VGND VGND VPWR VPWR _02920_ sky130_fd_sc_hd__a21bo_1
X_20262_ net3 _12073_ VGND VGND VPWR VPWR _12074_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_131_Right_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_94_Left_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22001_ _02008_ _01910_ pid_d.prev_error\[7\] VGND VGND VPWR VPWR _02009_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_179_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20193_ net952 _11954_ _11934_ VGND VGND VPWR VPWR _12018_ sky130_fd_sc_hd__and3b_1
XFILLER_0_11_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput108 pid_d_data[5] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_1
Xinput119 pid_q_addr[14] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_1
X_23952_ _03813_ _03815_ VGND VGND VPWR VPWR _03816_ sky130_fd_sc_hd__xor2_1
X_22903_ _02109_ _02787_ net5354 VGND VGND VPWR VPWR _02796_ sky130_fd_sc_hd__o21ba_1
X_23883_ _03734_ _03747_ VGND VGND VPWR VPWR _03748_ sky130_fd_sc_hd__xnor2_1
X_25622_ clknet_leaf_115_clk _00495_ net8330 VGND VGND VPWR VPWR cordic0.slte0.opA\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_22834_ _02727_ _02728_ _02733_ VGND VGND VPWR VPWR _02734_ sky130_fd_sc_hd__a21o_1
XFILLER_0_195_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25553_ clknet_leaf_64_clk net6572 net8662 VGND VGND VPWR VPWR matmul0.done_pass
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_177_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22765_ net4302 net8940 VGND VGND VPWR VPWR _02688_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24504_ _04302_ _04359_ net2017 VGND VGND VPWR VPWR _04361_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_176_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21716_ _01649_ _01726_ VGND VGND VPWR VPWR _01727_ sky130_fd_sc_hd__xor2_1
X_25484_ clknet_leaf_45_clk _00364_ net8788 VGND VGND VPWR VPWR svm0.tA\[6\] sky130_fd_sc_hd__dfrtp_1
Xwire8003 net8004 VGND VGND VPWR VPWR net8003 sky130_fd_sc_hd__clkbuf_1
Xwire8014 net8015 VGND VGND VPWR VPWR net8014 sky130_fd_sc_hd__clkbuf_1
X_22696_ pid_d.ki\[9\] net2446 net3696 pid_d.kp\[9\] VGND VGND VPWR VPWR _02639_ sky130_fd_sc_hd__a22o_1
Xwire8025 net8026 VGND VGND VPWR VPWR net8025 sky130_fd_sc_hd__clkbuf_1
Xwire8036 net8037 VGND VGND VPWR VPWR net8036 sky130_fd_sc_hd__clkbuf_1
X_24435_ net3753 _04287_ _04292_ net4515 VGND VGND VPWR VPWR _04293_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7302 net7303 VGND VGND VPWR VPWR net7302 sky130_fd_sc_hd__dlymetal6s2s_1
X_21647_ _01556_ _01566_ _01657_ VGND VGND VPWR VPWR _01658_ sky130_fd_sc_hd__o21ai_2
Xfanout6506 cordic0.gm0.iter\[0\] VGND VGND VPWR VPWR net6506 sky130_fd_sc_hd__buf_1
XFILLER_0_35_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3000 _00003_ VGND VGND VPWR VPWR net3000 sky130_fd_sc_hd__clkbuf_1
Xwire7313 net7314 VGND VGND VPWR VPWR net7313 sky130_fd_sc_hd__clkbuf_2
Xfanout6517 net6524 VGND VGND VPWR VPWR net6517 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7324 net7325 VGND VGND VPWR VPWR net7324 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire8069 net8070 VGND VGND VPWR VPWR net8069 sky130_fd_sc_hd__buf_1
XFILLER_0_35_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7335 matmul0.alpha_pass\[3\] VGND VGND VPWR VPWR net7335 sky130_fd_sc_hd__clkbuf_1
Xwire6601 net6602 VGND VGND VPWR VPWR net6601 sky130_fd_sc_hd__clkbuf_1
Xfanout6539 net6544 VGND VGND VPWR VPWR net6539 sky130_fd_sc_hd__buf_1
X_24366_ net2024 net2404 VGND VGND VPWR VPWR _04225_ sky130_fd_sc_hd__xor2_2
Xwire7346 net7347 VGND VGND VPWR VPWR net7346 sky130_fd_sc_hd__buf_1
Xfanout5816 net5819 VGND VGND VPWR VPWR net5816 sky130_fd_sc_hd__buf_1
X_21578_ _01484_ _01485_ _01483_ VGND VGND VPWR VPWR _01590_ sky130_fd_sc_hd__o21ai_1
Xwire6612 net6609 VGND VGND VPWR VPWR net6612 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire7357 net7358 VGND VGND VPWR VPWR net7357 sky130_fd_sc_hd__clkbuf_1
Xmax_length3055 _03373_ VGND VGND VPWR VPWR net3055 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6623 net6624 VGND VGND VPWR VPWR net6623 sky130_fd_sc_hd__clkbuf_1
Xwire7368 net7369 VGND VGND VPWR VPWR net7368 sky130_fd_sc_hd__buf_1
XFILLER_0_35_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6634 net6636 VGND VGND VPWR VPWR net6634 sky130_fd_sc_hd__buf_1
X_23317_ net4887 net4743 VGND VGND VPWR VPWR _03187_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6645 net6646 VGND VGND VPWR VPWR net6645 sky130_fd_sc_hd__clkbuf_1
Xwire5900 net5901 VGND VGND VPWR VPWR net5900 sky130_fd_sc_hd__clkbuf_1
Xwire5911 net5909 VGND VGND VPWR VPWR net5911 sky130_fd_sc_hd__clkbuf_2
X_20529_ net6901 net6853 net6890 net6840 net6490 net6513 VGND VGND VPWR VPWR _12315_
+ sky130_fd_sc_hd__mux4_2
X_24297_ _04155_ _04156_ net4603 VGND VGND VPWR VPWR _04157_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6667 net6668 VGND VGND VPWR VPWR net6667 sky130_fd_sc_hd__clkbuf_1
Xwire5922 net5923 VGND VGND VPWR VPWR net5922 sky130_fd_sc_hd__buf_1
XFILLER_0_132_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length1620 _04901_ VGND VGND VPWR VPWR net1620 sky130_fd_sc_hd__buf_1
Xwire5933 net5934 VGND VGND VPWR VPWR net5933 sky130_fd_sc_hd__buf_1
X_14050_ _06251_ _06312_ _06313_ VGND VGND VPWR VPWR _06314_ sky130_fd_sc_hd__o21ba_1
Xwire6689 svm0.counter\[14\] VGND VGND VPWR VPWR net6689 sky130_fd_sc_hd__buf_1
X_23248_ net4983 net4754 VGND VGND VPWR VPWR _03118_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5955 net5956 VGND VGND VPWR VPWR net5955 sky130_fd_sc_hd__buf_1
XFILLER_0_123_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5966 pid_d.curr_error\[11\] VGND VGND VPWR VPWR net5966 sky130_fd_sc_hd__buf_1
X_13001_ _05270_ _05271_ _05272_ _05273_ VGND VGND VPWR VPWR _05274_ sky130_fd_sc_hd__a211oi_1
Xwire5977 pid_d.curr_int\[8\] VGND VGND VPWR VPWR net5977 sky130_fd_sc_hd__clkbuf_2
X_23179_ net5089 net4757 VGND VGND VPWR VPWR _03049_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_0_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17740_ net6443 net6650 net6454 VGND VGND VPWR VPWR _09594_ sky130_fd_sc_hd__a21oi_1
X_14952_ net4139 VGND VGND VPWR VPWR _07026_ sky130_fd_sc_hd__buf_1
X_13903_ _06099_ _06101_ _06168_ VGND VGND VPWR VPWR _06169_ sky130_fd_sc_hd__o21a_1
X_17671_ net4011 svm0.tA\[4\] _09545_ net6740 _09550_ VGND VGND VPWR VPWR _09551_
+ sky130_fd_sc_hd__o221a_1
X_14883_ _06959_ VGND VGND VPWR VPWR _00212_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19410_ _11245_ _11246_ _11096_ VGND VGND VPWR VPWR _11247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16622_ matmul0.matmul_stage_inst.mult2\[1\] matmul0.matmul_stage_inst.mult1\[1\]
+ VGND VGND VPWR VPWR _08662_ sky130_fd_sc_hd__xor2_1
X_13834_ net7720 net2952 net3671 VGND VGND VPWR VPWR _06101_ sky130_fd_sc_hd__and3_1
XFILLER_0_159_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19341_ _10812_ _11177_ _11120_ VGND VGND VPWR VPWR _11178_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13765_ _06025_ _06026_ _06031_ _06032_ VGND VGND VPWR VPWR _06033_ sky130_fd_sc_hd__a211o_1
X_16553_ _08608_ _08611_ VGND VGND VPWR VPWR _08612_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_186_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15504_ _07479_ _07480_ VGND VGND VPWR VPWR _07577_ sky130_fd_sc_hd__or2_1
Xfanout8420 net8424 VGND VGND VPWR VPWR net8420 sky130_fd_sc_hd__clkbuf_2
X_12716_ _04985_ _04988_ VGND VGND VPWR VPWR _04989_ sky130_fd_sc_hd__xnor2_4
X_19272_ _10966_ _10968_ VGND VGND VPWR VPWR _11109_ sky130_fd_sc_hd__and2_1
X_13696_ _05896_ _05898_ _05897_ VGND VGND VPWR VPWR _05965_ sky130_fd_sc_hd__a21oi_1
X_16484_ net208 _08544_ VGND VGND VPWR VPWR _08545_ sky130_fd_sc_hd__xnor2_1
Xfanout8453 net8479 VGND VGND VPWR VPWR net8453 sky130_fd_sc_hd__buf_1
X_18223_ _10029_ _10073_ VGND VGND VPWR VPWR _10074_ sky130_fd_sc_hd__or2_1
X_12647_ _04919_ VGND VGND VPWR VPWR _04920_ sky130_fd_sc_hd__buf_1
X_15435_ net3423 net2689 VGND VGND VPWR VPWR _07509_ sky130_fd_sc_hd__xnor2_1
Xfanout8475 net8486 VGND VGND VPWR VPWR net8475 sky130_fd_sc_hd__clkbuf_1
Xfanout7741 net7750 VGND VGND VPWR VPWR net7741 sky130_fd_sc_hd__buf_1
XFILLER_0_109_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout7763 net7772 VGND VGND VPWR VPWR net7763 sky130_fd_sc_hd__clkbuf_1
Xwire8570 net8572 VGND VGND VPWR VPWR net8570 sky130_fd_sc_hd__buf_1
XFILLER_0_5_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18154_ _09758_ _10004_ VGND VGND VPWR VPWR _10005_ sky130_fd_sc_hd__xor2_1
X_15366_ net2233 net2249 net2704 VGND VGND VPWR VPWR _07440_ sky130_fd_sc_hd__and3_1
X_12578_ matmul0.state\[1\] _04864_ net8976 VGND VGND VPWR VPWR _00014_ sky130_fd_sc_hd__a21o_1
Xwire8592 net8593 VGND VGND VPWR VPWR net8592 sky130_fd_sc_hd__buf_1
Xmax_length4290 net4291 VGND VGND VPWR VPWR net4290 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17105_ _09039_ net772 _09061_ VGND VGND VPWR VPWR _09062_ sky130_fd_sc_hd__o21a_1
Xwire260 net261 VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__clkbuf_1
X_14317_ net6448 _06530_ net6443 _06538_ VGND VGND VPWR VPWR _06539_ sky130_fd_sc_hd__or4_1
XFILLER_0_29_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire271 net272 VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__clkbuf_1
X_18085_ net3969 net3995 _09849_ VGND VGND VPWR VPWR _09936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15297_ net4092 net4089 VGND VGND VPWR VPWR _07371_ sky130_fd_sc_hd__nor2_1
Xwire282 _06275_ VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__buf_1
Xwire7891 net7892 VGND VGND VPWR VPWR net7891 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire293 _04250_ VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14248_ net6508 net6496 VGND VGND VPWR VPWR _06503_ sky130_fd_sc_hd__or2_1
X_17036_ net3336 net1804 _08995_ VGND VGND VPWR VPWR _08996_ sky130_fd_sc_hd__or3_1
XFILLER_0_68_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14179_ _06409_ net833 VGND VGND VPWR VPWR _06439_ sky130_fd_sc_hd__nor2_2
XFILLER_0_110_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18987_ net6312 net6352 VGND VGND VPWR VPWR _10824_ sky130_fd_sc_hd__xor2_1
XFILLER_0_84_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17938_ _09781_ _09784_ _09786_ _09686_ _09788_ VGND VGND VPWR VPWR _09789_ sky130_fd_sc_hd__o221a_1
X_17869_ _09050_ net3268 VGND VGND VPWR VPWR _09720_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_178_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19608_ net6065 _11444_ VGND VGND VPWR VPWR _11445_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20880_ net5954 net5472 VGND VGND VPWR VPWR _00896_ sky130_fd_sc_hd__and2_1
XFILLER_0_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19539_ _11035_ VGND VGND VPWR VPWR _11376_ sky130_fd_sc_hd__buf_1
Xmax_length5908 net5903 VGND VGND VPWR VPWR net5908 sky130_fd_sc_hd__buf_1
XFILLER_0_191_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22550_ net9012 net2049 _02537_ VGND VGND VPWR VPWR _00547_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21501_ _01511_ _01513_ VGND VGND VPWR VPWR _01514_ sky130_fd_sc_hd__xor2_1
XFILLER_0_146_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22481_ net5407 net5434 net5647 VGND VGND VPWR VPWR _02482_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_63_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24220_ _04079_ _04080_ VGND VGND VPWR VPWR _04081_ sky130_fd_sc_hd__xor2_2
XFILLER_0_16_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21432_ net5456 net5890 net2479 VGND VGND VPWR VPWR _01445_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24151_ net1658 _04012_ VGND VGND VPWR VPWR _04013_ sky130_fd_sc_hd__xor2_1
Xwire5207 net5208 VGND VGND VPWR VPWR net5207 sky130_fd_sc_hd__clkbuf_2
X_21363_ _01373_ _01376_ VGND VGND VPWR VPWR _01377_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5229 net5230 VGND VGND VPWR VPWR net5229 sky130_fd_sc_hd__clkbuf_1
X_23102_ _02969_ _02970_ VGND VGND VPWR VPWR _02972_ sky130_fd_sc_hd__nor2_1
X_20314_ net4041 net6477 VGND VGND VPWR VPWR _12118_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput90 pid_d_addr[3] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_1
X_24082_ net376 _03944_ VGND VGND VPWR VPWR _03945_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21294_ net5473 _01308_ VGND VGND VPWR VPWR _01309_ sky130_fd_sc_hd__nand2_1
Xwire4528 net4529 VGND VGND VPWR VPWR net4528 sky130_fd_sc_hd__clkbuf_1
Xwire4539 net4533 VGND VGND VPWR VPWR net4539 sky130_fd_sc_hd__buf_1
XFILLER_0_3_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23033_ _02900_ _02901_ VGND VGND VPWR VPWR _02903_ sky130_fd_sc_hd__nor2_1
Xwire3805 _01066_ VGND VGND VPWR VPWR net3805 sky130_fd_sc_hd__buf_1
XFILLER_0_12_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3816 net3817 VGND VGND VPWR VPWR net3816 sky130_fd_sc_hd__buf_1
X_20245_ _12060_ VGND VGND VPWR VPWR _00474_ sky130_fd_sc_hd__clkbuf_1
Xwire3827 net3828 VGND VGND VPWR VPWR net3827 sky130_fd_sc_hd__clkbuf_1
Xwire3838 _00882_ VGND VGND VPWR VPWR net3838 sky130_fd_sc_hd__clkbuf_1
Xwire3849 net3850 VGND VGND VPWR VPWR net3849 sky130_fd_sc_hd__buf_1
X_20176_ _12000_ _12001_ net6042 VGND VGND VPWR VPWR _12002_ sky130_fd_sc_hd__and3b_1
X_24984_ pid_q.kp\[11\] _04724_ net1634 VGND VGND VPWR VPWR _04747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23935_ _03715_ _03720_ _03798_ VGND VGND VPWR VPWR _03799_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23866_ _03722_ _03730_ VGND VGND VPWR VPWR _03731_ sky130_fd_sc_hd__xnor2_2
Xmax_length8567 net8568 VGND VGND VPWR VPWR net8567 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_54_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25605_ clknet_leaf_109_clk _00478_ net8344 VGND VGND VPWR VPWR cordic0.slte0.opB\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_22817_ pid_d.out\[0\] net2463 net2034 net479 _02719_ VGND VGND VPWR VPWR _02720_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_168_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23797_ _03661_ _03568_ _03570_ _03662_ VGND VGND VPWR VPWR _03663_ sky130_fd_sc_hd__a31o_1
XFILLER_0_183_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13550_ _05813_ _05820_ VGND VGND VPWR VPWR _05821_ sky130_fd_sc_hd__xor2_2
Xmax_length7899 net7888 VGND VGND VPWR VPWR net7899 sky130_fd_sc_hd__buf_1
X_25536_ clknet_leaf_33_clk _00416_ net8687 VGND VGND VPWR VPWR pid_q.prev_int\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_22748_ net9234 _02676_ net1690 VGND VGND VPWR VPWR _02677_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout7004 cordic0.vec\[1\]\[6\] VGND VGND VPWR VPWR net7004 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_95_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout7015 net7023 VGND VGND VPWR VPWR net7015 sky130_fd_sc_hd__clkbuf_1
X_25467_ clknet_leaf_53_clk _00347_ net8807 VGND VGND VPWR VPWR svm0.tB\[5\] sky130_fd_sc_hd__dfrtp_1
X_13481_ _05749_ _05750_ net1310 VGND VGND VPWR VPWR _05754_ sky130_fd_sc_hd__a21o_1
XFILLER_0_137_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22679_ _02627_ net5606 net2448 VGND VGND VPWR VPWR _02628_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15220_ net1545 _07293_ VGND VGND VPWR VPWR _07294_ sky130_fd_sc_hd__xnor2_1
X_24418_ _04274_ _04275_ net4581 VGND VGND VPWR VPWR _04276_ sky130_fd_sc_hd__mux2_1
Xwire7132 net7133 VGND VGND VPWR VPWR net7132 sky130_fd_sc_hd__buf_1
XFILLER_0_152_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25398_ clknet_leaf_70_clk _00281_ net8448 VGND VGND VPWR VPWR matmul0.a\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6420 cordic0.slte0.opB\[2\] VGND VGND VPWR VPWR net6420 sky130_fd_sc_hd__clkbuf_1
Xfanout6358 net6365 VGND VGND VPWR VPWR net6358 sky130_fd_sc_hd__buf_1
XFILLER_0_35_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15151_ net3562 _07224_ VGND VGND VPWR VPWR _07225_ sky130_fd_sc_hd__nand2_1
Xwire7165 matmul0.sin\[0\] VGND VGND VPWR VPWR net7165 sky130_fd_sc_hd__clkbuf_1
X_24349_ net4555 net4837 VGND VGND VPWR VPWR _04208_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6431 cordic0.sin\[0\] VGND VGND VPWR VPWR net6431 sky130_fd_sc_hd__clkbuf_1
Xwire7176 net7177 VGND VGND VPWR VPWR net7176 sky130_fd_sc_hd__clkbuf_1
Xwire6442 cordic0.out_valid VGND VGND VPWR VPWR net6442 sky130_fd_sc_hd__clkbuf_1
Xwire7187 matmul0.b\[3\] VGND VGND VPWR VPWR net7187 sky130_fd_sc_hd__clkbuf_1
Xwire7198 net7201 VGND VGND VPWR VPWR net7198 sky130_fd_sc_hd__clkbuf_1
X_14102_ _06356_ _06357_ net255 net254 VGND VGND VPWR VPWR _06364_ sky130_fd_sc_hd__a22o_1
Xfanout4923 pid_q.mult0.b\[9\] VGND VGND VPWR VPWR net4923 sky130_fd_sc_hd__buf_1
XFILLER_0_133_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6464 net6465 VGND VGND VPWR VPWR net6464 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5730 net5731 VGND VGND VPWR VPWR net5730 sky130_fd_sc_hd__buf_1
X_15082_ net2765 VGND VGND VPWR VPWR _07156_ sky130_fd_sc_hd__buf_1
Xfanout4945 pid_q.mult0.b\[8\] VGND VGND VPWR VPWR net4945 sky130_fd_sc_hd__buf_1
Xwire5741 net5739 VGND VGND VPWR VPWR net5741 sky130_fd_sc_hd__buf_1
Xwire6486 net6487 VGND VGND VPWR VPWR net6486 sky130_fd_sc_hd__clkbuf_1
Xfanout4956 pid_q.mult0.b\[7\] VGND VGND VPWR VPWR net4956 sky130_fd_sc_hd__clkbuf_1
Xwire5752 net5753 VGND VGND VPWR VPWR net5752 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6497 net6492 VGND VGND VPWR VPWR net6497 sky130_fd_sc_hd__buf_1
Xwire5763 net5764 VGND VGND VPWR VPWR net5763 sky130_fd_sc_hd__buf_1
X_14033_ _06220_ _06296_ _06219_ VGND VGND VPWR VPWR _06297_ sky130_fd_sc_hd__a21bo_1
X_18910_ net9062 net2288 net1449 _10750_ VGND VGND VPWR VPWR _00449_ sky130_fd_sc_hd__a31o_1
Xwire5785 net5783 VGND VGND VPWR VPWR net5785 sky130_fd_sc_hd__buf_1
Xmax_length1483 _08975_ VGND VGND VPWR VPWR net1483 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19890_ _11661_ _11721_ _11722_ net3858 VGND VGND VPWR VPWR _11723_ sky130_fd_sc_hd__o211a_1
Xwire5796 net5797 VGND VGND VPWR VPWR net5796 sky130_fd_sc_hd__clkbuf_1
X_18841_ net3222 _10683_ VGND VGND VPWR VPWR _10684_ sky130_fd_sc_hd__or2_1
X_18772_ net1437 net180 VGND VGND VPWR VPWR _10617_ sky130_fd_sc_hd__nor2_1
X_15984_ _08050_ net2205 VGND VGND VPWR VPWR _08052_ sky130_fd_sc_hd__or2b_1
X_17723_ net9189 net1457 net1790 net5170 VGND VGND VPWR VPWR _00428_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14935_ net6635 matmul0.matmul_stage_inst.d\[5\] net7413 net6535 VGND VGND VPWR VPWR
+ _07009_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17654_ _09522_ _09523_ _09524_ _09533_ VGND VGND VPWR VPWR _09534_ sky130_fd_sc_hd__or4_1
XFILLER_0_159_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14866_ matmul0.b\[5\] matmul0.matmul_stage_inst.f\[5\] net3606 VGND VGND VPWR VPWR
+ _06951_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16605_ _08652_ VGND VGND VPWR VPWR _00241_ sky130_fd_sc_hd__clkbuf_1
X_13817_ net449 _06084_ VGND VGND VPWR VPWR _06085_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_188_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17585_ net965 _09466_ net2155 VGND VGND VPWR VPWR _09467_ sky130_fd_sc_hd__o21ai_1
X_14797_ net9069 net3005 net2853 _06915_ VGND VGND VPWR VPWR _00170_ sky130_fd_sc_hd__o22a_1
X_19324_ _10837_ net3203 _11140_ VGND VGND VPWR VPWR _11161_ sky130_fd_sc_hd__mux2_1
XFILLER_0_187_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16536_ net1086 _08594_ VGND VGND VPWR VPWR _08595_ sky130_fd_sc_hd__nor2_1
X_13748_ _05869_ _06014_ _06015_ _05934_ VGND VGND VPWR VPWR _06016_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19255_ net1193 _11090_ _11091_ VGND VGND VPWR VPWR _11092_ sky130_fd_sc_hd__a21oi_1
X_16467_ net2625 net2218 _08525_ _08526_ _08527_ VGND VGND VPWR VPWR _08528_ sky130_fd_sc_hd__o311a_1
X_13679_ net3677 _05947_ net2947 net7810 net1939 VGND VGND VPWR VPWR _05948_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_155_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18206_ net2139 _09807_ _10056_ VGND VGND VPWR VPWR _10057_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_143_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15418_ net1865 net1864 VGND VGND VPWR VPWR _07492_ sky130_fd_sc_hd__nand2_1
X_19186_ _10909_ _10966_ _10968_ _10970_ net872 VGND VGND VPWR VPWR _11023_ sky130_fd_sc_hd__a221o_1
XFILLER_0_26_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16398_ net2245 net2642 net2639 VGND VGND VPWR VPWR _08460_ sky130_fd_sc_hd__or3_1
XFILLER_0_79_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18137_ _09930_ _09987_ _09901_ VGND VGND VPWR VPWR _09988_ sky130_fd_sc_hd__mux2_1
X_15349_ _07419_ _07420_ _07421_ _07422_ VGND VGND VPWR VPWR _07423_ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6892 net6899 VGND VGND VPWR VPWR net6892 sky130_fd_sc_hd__buf_2
Xhold104 matmul0.matmul_stage_inst.c\[15\] VGND VGND VPWR VPWR net9057 sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 svm0.vC\[7\] VGND VGND VPWR VPWR net9068 sky130_fd_sc_hd__dlygate4sd3_1
X_18068_ net3256 net7146 net3994 VGND VGND VPWR VPWR _09919_ sky130_fd_sc_hd__a21oi_1
Xhold126 pid_d.curr_int\[2\] VGND VGND VPWR VPWR net9079 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 svm0.tB\[6\] VGND VGND VPWR VPWR net9090 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold148 cordic0.sin\[12\] VGND VGND VPWR VPWR net9101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 svm0.tC\[9\] VGND VGND VPWR VPWR net9112 sky130_fd_sc_hd__dlygate4sd3_1
X_17019_ _08978_ _08979_ VGND VGND VPWR VPWR _08980_ sky130_fd_sc_hd__nand2_2
XFILLER_0_42_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20030_ net2497 _11859_ VGND VGND VPWR VPWR _11860_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21981_ _01879_ _01987_ _01988_ _01883_ VGND VGND VPWR VPWR _01989_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23720_ _03584_ _03585_ VGND VGND VPWR VPWR _03586_ sky130_fd_sc_hd__nand2_1
X_20932_ _00945_ _00946_ VGND VGND VPWR VPWR _00948_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23651_ net3748 _03395_ _03517_ VGND VGND VPWR VPWR _03518_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_135_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6417 cordic0.slte0.opB\[5\] VGND VGND VPWR VPWR net6417 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20863_ _12537_ _12538_ VGND VGND VPWR VPWR _00879_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length5705 net5701 VGND VGND VPWR VPWR net5705 sky130_fd_sc_hd__buf_1
X_22602_ net7265 _02574_ VGND VGND VPWR VPWR _02577_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23582_ _03349_ _03368_ net1028 VGND VGND VPWR VPWR _03450_ sky130_fd_sc_hd__o21a_1
XFILLER_0_187_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20794_ _12559_ net2484 VGND VGND VPWR VPWR _00810_ sky130_fd_sc_hd__xnor2_2
X_25321_ clknet_leaf_74_clk _00204_ net8464 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.f\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22533_ pid_d.curr_error\[4\] net2380 net2047 VGND VGND VPWR VPWR _02529_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25252_ clknet_leaf_88_clk _00135_ net8430 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.a\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_22464_ pid_d.prev_int\[14\] _02397_ pid_d.curr_int\[14\] VGND VGND VPWR VPWR _02465_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length616 _09276_ VGND VGND VPWR VPWR net616 sky130_fd_sc_hd__buf_1
X_24203_ _04062_ _04063_ VGND VGND VPWR VPWR _04064_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length638 _04035_ VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__clkbuf_1
X_21415_ pid_d.prev_error\[0\] net5973 pid_d.prev_error\[1\] net5972 VGND VGND VPWR
+ VPWR _01429_ sky130_fd_sc_hd__a22o_1
X_25183_ clknet_leaf_67_clk _00072_ net8450 VGND VGND VPWR VPWR matmul0.a_in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire5004 net5005 VGND VGND VPWR VPWR net5004 sky130_fd_sc_hd__clkbuf_1
X_22395_ _02330_ _02333_ _02334_ _02331_ VGND VGND VPWR VPWR _02397_ sky130_fd_sc_hd__o31a_1
Xwire5015 net5016 VGND VGND VPWR VPWR net5015 sky130_fd_sc_hd__buf_1
Xwire5026 net5030 VGND VGND VPWR VPWR net5026 sky130_fd_sc_hd__clkbuf_1
X_24134_ _03878_ _03883_ _03995_ VGND VGND VPWR VPWR _03996_ sky130_fd_sc_hd__a21o_1
Xwire5037 net5038 VGND VGND VPWR VPWR net5037 sky130_fd_sc_hd__buf_1
X_21346_ net5807 net5511 VGND VGND VPWR VPWR _01360_ sky130_fd_sc_hd__nand2_2
Xwire5048 net5049 VGND VGND VPWR VPWR net5048 sky130_fd_sc_hd__buf_1
Xwire4303 net4304 VGND VGND VPWR VPWR net4303 sky130_fd_sc_hd__buf_1
XFILLER_0_20_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5059 net5060 VGND VGND VPWR VPWR net5059 sky130_fd_sc_hd__buf_1
XFILLER_0_103_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4325 net4326 VGND VGND VPWR VPWR net4325 sky130_fd_sc_hd__buf_1
XFILLER_0_103_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24065_ net4704 net3747 _03830_ VGND VGND VPWR VPWR _03928_ sky130_fd_sc_hd__or3b_1
Xwire4336 net4337 VGND VGND VPWR VPWR net4336 sky130_fd_sc_hd__buf_1
Xwire4347 net4348 VGND VGND VPWR VPWR net4347 sky130_fd_sc_hd__clkbuf_1
Xwire3602 net3603 VGND VGND VPWR VPWR net3602 sky130_fd_sc_hd__buf_1
X_21277_ _01290_ _01291_ VGND VGND VPWR VPWR _01292_ sky130_fd_sc_hd__xor2_1
Xwire4358 net4352 VGND VGND VPWR VPWR net4358 sky130_fd_sc_hd__buf_1
Xwire4369 net4375 VGND VGND VPWR VPWR net4369 sky130_fd_sc_hd__clkbuf_1
Xwire3624 net3625 VGND VGND VPWR VPWR net3624 sky130_fd_sc_hd__buf_1
X_23016_ _02880_ _02885_ VGND VGND VPWR VPWR _02886_ sky130_fd_sc_hd__and2_1
Xwire3635 net3636 VGND VGND VPWR VPWR net3635 sky130_fd_sc_hd__buf_1
Xwire2901 _06518_ VGND VGND VPWR VPWR net2901 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3646 _06527_ VGND VGND VPWR VPWR net3646 sky130_fd_sc_hd__buf_1
XFILLER_0_21_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20228_ net10 _12043_ net8122 VGND VGND VPWR VPWR _12047_ sky130_fd_sc_hd__a21oi_1
Xwire3657 net3658 VGND VGND VPWR VPWR net3657 sky130_fd_sc_hd__clkbuf_1
Xwire2912 net2913 VGND VGND VPWR VPWR net2912 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2923 net2924 VGND VGND VPWR VPWR net2923 sky130_fd_sc_hd__buf_1
Xwire3668 _06505_ VGND VGND VPWR VPWR net3668 sky130_fd_sc_hd__buf_1
Xwire3679 net3680 VGND VGND VPWR VPWR net3679 sky130_fd_sc_hd__buf_1
Xwire2934 net2935 VGND VGND VPWR VPWR net2934 sky130_fd_sc_hd__clkbuf_1
Xwire2945 _05689_ VGND VGND VPWR VPWR net2945 sky130_fd_sc_hd__clkbuf_1
X_20159_ _11980_ _11981_ _11983_ _11985_ VGND VGND VPWR VPWR _11986_ sky130_fd_sc_hd__o211a_1
Xwire2967 net2968 VGND VGND VPWR VPWR net2967 sky130_fd_sc_hd__buf_1
Xwire2978 net2979 VGND VGND VPWR VPWR net2978 sky130_fd_sc_hd__buf_1
Xwire2989 _04906_ VGND VGND VPWR VPWR net2989 sky130_fd_sc_hd__buf_1
X_12981_ _05171_ _05172_ net7738 net1617 VGND VGND VPWR VPWR _05254_ sky130_fd_sc_hd__o211a_1
X_24967_ _04738_ VGND VGND VPWR VPWR _00763_ sky130_fd_sc_hd__clkbuf_1
X_14720_ net7148 _06858_ net7457 VGND VGND VPWR VPWR _06860_ sky130_fd_sc_hd__and3b_1
XFILLER_0_169_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23918_ net4611 net4880 VGND VGND VPWR VPWR _03782_ sky130_fd_sc_hd__nand2_1
Xmax_length8342 net8338 VGND VGND VPWR VPWR net8342 sky130_fd_sc_hd__buf_1
X_24898_ pid_q.ki\[14\] net3711 net3701 pid_q.kp\[14\] VGND VGND VPWR VPWR _04690_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14651_ net7440 net7175 net2874 VGND VGND VPWR VPWR _06810_ sky130_fd_sc_hd__and3_1
X_23849_ _03623_ _03625_ _03624_ VGND VGND VPWR VPWR _03714_ sky130_fd_sc_hd__o21ai_1
Xmax_length8397 net8394 VGND VGND VPWR VPWR net8397 sky130_fd_sc_hd__buf_1
XFILLER_0_19_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13602_ _05783_ _05870_ _05871_ VGND VGND VPWR VPWR _05872_ sky130_fd_sc_hd__a21o_2
X_17370_ svm0.delta\[3\] VGND VGND VPWR VPWR _09281_ sky130_fd_sc_hd__inv_2
X_14582_ net9115 _06652_ net318 net2886 VGND VGND VPWR VPWR _00113_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6984 net6981 VGND VGND VPWR VPWR net6984 sky130_fd_sc_hd__buf_1
X_16321_ net2815 net2682 net1250 _08383_ VGND VGND VPWR VPWR _08384_ sky130_fd_sc_hd__o211a_1
X_25519_ clknet_leaf_42_clk _00399_ net8777 VGND VGND VPWR VPWR svm0.counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13533_ _05801_ _05802_ _05799_ _05800_ VGND VGND VPWR VPWR _05804_ sky130_fd_sc_hd__a211o_1
XFILLER_0_54_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout6100 net6108 VGND VGND VPWR VPWR net6100 sky130_fd_sc_hd__buf_1
XFILLER_0_82_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19040_ _10876_ net3904 VGND VGND VPWR VPWR _10877_ sky130_fd_sc_hd__xnor2_1
X_13464_ _05585_ _05586_ _05736_ VGND VGND VPWR VPWR _05737_ sky130_fd_sc_hd__o21a_1
X_16252_ net2691 _08314_ _08315_ VGND VGND VPWR VPWR _08316_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_180_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6122 cordic0.vec\[0\]\[11\] VGND VGND VPWR VPWR net6122 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15203_ _07272_ _07273_ _07276_ VGND VGND VPWR VPWR _07277_ sky130_fd_sc_hd__o21a_1
XFILLER_0_168_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13395_ _05401_ _05662_ VGND VGND VPWR VPWR _05668_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16183_ net1089 net983 _08200_ VGND VGND VPWR VPWR _08248_ sky130_fd_sc_hd__a21o_1
Xfanout6177 net6185 VGND VGND VPWR VPWR net6177 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_180_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15134_ net2777 net2743 VGND VGND VPWR VPWR _07208_ sky130_fd_sc_hd__nor2_1
Xwire6272 net6274 VGND VGND VPWR VPWR net6272 sky130_fd_sc_hd__buf_1
Xwire6283 net6284 VGND VGND VPWR VPWR net6283 sky130_fd_sc_hd__buf_1
Xfanout4753 net4762 VGND VGND VPWR VPWR net4753 sky130_fd_sc_hd__buf_1
Xwire5560 net5561 VGND VGND VPWR VPWR net5560 sky130_fd_sc_hd__clkbuf_1
X_15065_ net4120 net4115 VGND VGND VPWR VPWR _07139_ sky130_fd_sc_hd__or2_1
X_19942_ net6009 _11773_ VGND VGND VPWR VPWR _11774_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5571 net5572 VGND VGND VPWR VPWR net5571 sky130_fd_sc_hd__clkbuf_1
Xwire5582 net5583 VGND VGND VPWR VPWR net5582 sky130_fd_sc_hd__clkbuf_1
Xwire5593 net5594 VGND VGND VPWR VPWR net5593 sky130_fd_sc_hd__buf_1
X_14016_ _06278_ _06263_ _06279_ VGND VGND VPWR VPWR _06280_ sky130_fd_sc_hd__o21ai_1
Xwire4870 net4862 VGND VGND VPWR VPWR net4870 sky130_fd_sc_hd__clkbuf_1
X_19873_ net3141 net2100 _11625_ net6064 VGND VGND VPWR VPWR _11706_ sky130_fd_sc_hd__a22o_1
Xwire4881 net4882 VGND VGND VPWR VPWR net4881 sky130_fd_sc_hd__buf_1
Xwire4892 net4893 VGND VGND VPWR VPWR net4892 sky130_fd_sc_hd__clkbuf_1
X_18824_ net6837 net3920 net3983 VGND VGND VPWR VPWR _10667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18755_ _10595_ _10599_ VGND VGND VPWR VPWR _10600_ sky130_fd_sc_hd__xor2_1
X_15967_ _07940_ _07947_ _07946_ VGND VGND VPWR VPWR _08035_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17706_ _09576_ net8864 pid_q.state\[4\] _09581_ VGND VGND VPWR VPWR _09582_ sky130_fd_sc_hd__and4b_1
XFILLER_0_136_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14918_ net6619 net6644 net7385 VGND VGND VPWR VPWR _06992_ sky130_fd_sc_hd__o21a_1
XFILLER_0_188_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18686_ _10530_ _10531_ VGND VGND VPWR VPWR _10532_ sky130_fd_sc_hd__xor2_1
X_15898_ _07963_ _07966_ VGND VGND VPWR VPWR _07967_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17637_ net2153 _09515_ net2566 VGND VGND VPWR VPWR _09518_ sky130_fd_sc_hd__a21oi_1
X_14849_ net9183 matmul0.matmul_stage_inst.e\[13\] net3608 VGND VGND VPWR VPWR _06942_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17568_ net6737 _09446_ _09447_ _09448_ _09449_ VGND VGND VPWR VPWR _09450_ sky130_fd_sc_hd__o221a_1
XFILLER_0_14_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19307_ net3207 _10823_ _11141_ _11143_ VGND VGND VPWR VPWR _11144_ sky130_fd_sc_hd__a31o_1
X_16519_ _08529_ net1243 VGND VGND VPWR VPWR _08579_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17499_ _09307_ _09383_ net6705 VGND VGND VPWR VPWR _09387_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_184_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19238_ net6323 net6221 VGND VGND VPWR VPWR _11075_ sky130_fd_sc_hd__or2b_1
XPHY_EDGE_ROW_12_Left_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap3360 net9246 VGND VGND VPWR VPWR net3360 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19169_ _10940_ _11003_ _11005_ VGND VGND VPWR VPWR _11006_ sky130_fd_sc_hd__o21a_1
XFILLER_0_83_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21200_ _01115_ _01116_ net807 VGND VGND VPWR VPWR _01216_ sky130_fd_sc_hd__o21bai_1
X_22180_ _02182_ _02111_ _02184_ VGND VGND VPWR VPWR _02185_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21131_ _01145_ _01146_ VGND VGND VPWR VPWR _01147_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21062_ net862 _01077_ VGND VGND VPWR VPWR _01078_ sky130_fd_sc_hd__xnor2_1
Xwire2219 net2220 VGND VGND VPWR VPWR net2219 sky130_fd_sc_hd__buf_1
X_20013_ _11740_ _11835_ _11842_ VGND VGND VPWR VPWR _11843_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_21_Left_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25870_ clknet_leaf_17_clk _00743_ net8631 VGND VGND VPWR VPWR pid_q.mult0.a\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1507 _08417_ VGND VGND VPWR VPWR net1507 sky130_fd_sc_hd__buf_1
Xwire1518 net1519 VGND VGND VPWR VPWR net1518 sky130_fd_sc_hd__buf_1
Xwire1529 _07809_ VGND VGND VPWR VPWR net1529 sky130_fd_sc_hd__buf_1
X_24821_ _04540_ VGND VGND VPWR VPWR _04643_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24752_ net5254 net3031 VGND VGND VPWR VPWR _04583_ sky130_fd_sc_hd__nand2_1
X_21964_ _01969_ net1170 VGND VGND VPWR VPWR _01972_ sky130_fd_sc_hd__xor2_2
XFILLER_0_154_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23703_ _03567_ _03475_ _03476_ _03569_ VGND VGND VPWR VPWR _03570_ sky130_fd_sc_hd__a31o_1
X_20915_ _00927_ net1186 _00930_ VGND VGND VPWR VPWR _00931_ sky130_fd_sc_hd__o21ba_1
X_24683_ net5166 net3021 _04509_ VGND VGND VPWR VPWR _04524_ sky130_fd_sc_hd__and3_1
Xmax_length6203 net6200 VGND VGND VPWR VPWR net6203 sky130_fd_sc_hd__buf_1
X_21895_ _01742_ _01802_ _01714_ VGND VGND VPWR VPWR _01904_ sky130_fd_sc_hd__a21bo_1
X_23634_ _03499_ _03500_ VGND VGND VPWR VPWR _03501_ sky130_fd_sc_hd__xor2_1
X_20846_ _12520_ _12547_ _00861_ VGND VGND VPWR VPWR _00862_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_7_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23565_ net4749 net4826 VGND VGND VPWR VPWR _03433_ sky130_fd_sc_hd__nand2_2
XFILLER_0_119_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_30_Left_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20777_ net5557 net5795 VGND VGND VPWR VPWR _12548_ sky130_fd_sc_hd__nand2_2
X_22516_ net380 net204 net4315 net2489 VGND VGND VPWR VPWR _02517_ sky130_fd_sc_hd__o211a_1
X_25304_ clknet_leaf_69_clk _00187_ net8451 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.e\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire804 _01816_ VGND VGND VPWR VPWR net804 sky130_fd_sc_hd__clkbuf_1
Xwire815 net816 VGND VGND VPWR VPWR net815 sky130_fd_sc_hd__dlymetal6s2s_1
X_23496_ _03289_ _03291_ _03287_ VGND VGND VPWR VPWR _03365_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_174_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4878 net4874 VGND VGND VPWR VPWR net4878 sky130_fd_sc_hd__clkbuf_1
Xwire826 _07961_ VGND VGND VPWR VPWR net826 sky130_fd_sc_hd__buf_1
XFILLER_0_88_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire837 net838 VGND VGND VPWR VPWR net837 sky130_fd_sc_hd__buf_1
XFILLER_0_162_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire848 _05402_ VGND VGND VPWR VPWR net848 sky130_fd_sc_hd__buf_1
XFILLER_0_107_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25235_ clknet_leaf_17_clk net3007 net8631 VGND VGND VPWR VPWR pid_q.state\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22447_ _02440_ _02448_ VGND VGND VPWR VPWR _02449_ sky130_fd_sc_hd__xnor2_1
Xwire859 _02158_ VGND VGND VPWR VPWR net859 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13180_ _05451_ _05452_ VGND VGND VPWR VPWR _05453_ sky130_fd_sc_hd__xor2_1
X_25166_ clknet_leaf_55_clk _00055_ net8728 VGND VGND VPWR VPWR svm0.periodTop\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_22378_ _02313_ _02316_ _02281_ VGND VGND VPWR VPWR _02381_ sky130_fd_sc_hd__o21a_1
Xwire4100 _07143_ VGND VGND VPWR VPWR net4100 sky130_fd_sc_hd__clkbuf_1
X_24117_ net4590 net4852 VGND VGND VPWR VPWR _03979_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4111 net4112 VGND VGND VPWR VPWR net4111 sky130_fd_sc_hd__buf_1
X_21329_ net5739 net5560 VGND VGND VPWR VPWR _01343_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4122 net4123 VGND VGND VPWR VPWR net4122 sky130_fd_sc_hd__buf_1
X_25097_ net4400 VGND VGND VPWR VPWR _04841_ sky130_fd_sc_hd__inv_2
Xwire4133 net4134 VGND VGND VPWR VPWR net4133 sky130_fd_sc_hd__clkbuf_1
Xwire4144 net4145 VGND VGND VPWR VPWR net4144 sky130_fd_sc_hd__clkbuf_1
Xwire3410 net3411 VGND VGND VPWR VPWR net3410 sky130_fd_sc_hd__clkbuf_1
Xwire4155 _07013_ VGND VGND VPWR VPWR net4155 sky130_fd_sc_hd__clkbuf_1
X_24048_ _03813_ _03815_ _03910_ VGND VGND VPWR VPWR _03911_ sky130_fd_sc_hd__o21ai_1
Xwire3421 net3422 VGND VGND VPWR VPWR net3421 sky130_fd_sc_hd__buf_1
Xwire4166 net4167 VGND VGND VPWR VPWR net4166 sky130_fd_sc_hd__buf_1
Xwire3432 net3433 VGND VGND VPWR VPWR net3432 sky130_fd_sc_hd__buf_1
Xwire4177 _06999_ VGND VGND VPWR VPWR net4177 sky130_fd_sc_hd__clkbuf_1
Xwire3443 _07303_ VGND VGND VPWR VPWR net3443 sky130_fd_sc_hd__buf_1
Xwire4188 net4189 VGND VGND VPWR VPWR net4188 sky130_fd_sc_hd__clkbuf_1
Xwire3454 net3455 VGND VGND VPWR VPWR net3454 sky130_fd_sc_hd__clkbuf_1
Xwire4199 net4200 VGND VGND VPWR VPWR net4199 sky130_fd_sc_hd__buf_1
Xwire3465 net3466 VGND VGND VPWR VPWR net3465 sky130_fd_sc_hd__buf_1
Xwire2720 _07287_ VGND VGND VPWR VPWR net2720 sky130_fd_sc_hd__buf_1
X_16870_ net6495 net6477 VGND VGND VPWR VPWR _08835_ sky130_fd_sc_hd__or2_1
Xwire3476 net3477 VGND VGND VPWR VPWR net3476 sky130_fd_sc_hd__clkbuf_1
Xwire3487 _07141_ VGND VGND VPWR VPWR net3487 sky130_fd_sc_hd__buf_1
Xwire2742 _07226_ VGND VGND VPWR VPWR net2742 sky130_fd_sc_hd__buf_1
Xwire2753 net2754 VGND VGND VPWR VPWR net2753 sky130_fd_sc_hd__buf_1
Xwire3498 net3499 VGND VGND VPWR VPWR net3498 sky130_fd_sc_hd__buf_1
Xwire2764 net2765 VGND VGND VPWR VPWR net2764 sky130_fd_sc_hd__buf_1
X_15821_ _07775_ _07798_ net887 VGND VGND VPWR VPWR _07891_ sky130_fd_sc_hd__o21a_1
Xwire2775 _07146_ VGND VGND VPWR VPWR net2775 sky130_fd_sc_hd__clkbuf_1
Xwire2786 net2787 VGND VGND VPWR VPWR net2786 sky130_fd_sc_hd__buf_1
Xwire2797 net2798 VGND VGND VPWR VPWR net2797 sky130_fd_sc_hd__buf_1
XFILLER_0_99_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18540_ _10387_ net2541 _10388_ net6815 VGND VGND VPWR VPWR _10389_ sky130_fd_sc_hd__a211o_1
X_15752_ _07730_ _07822_ VGND VGND VPWR VPWR _07823_ sky130_fd_sc_hd__xnor2_1
X_12964_ _05030_ _05236_ VGND VGND VPWR VPWR _05237_ sky130_fd_sc_hd__or2_1
X_14703_ net7152 net7151 _06842_ VGND VGND VPWR VPWR _06847_ sky130_fd_sc_hd__or3_1
X_18471_ _10309_ _10314_ VGND VGND VPWR VPWR _10321_ sky130_fd_sc_hd__or2_1
X_15683_ net2717 net3434 VGND VGND VPWR VPWR _07754_ sky130_fd_sc_hd__nor2_1
XFILLER_0_169_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12895_ _05153_ _05154_ _05166_ _05167_ VGND VGND VPWR VPWR _05168_ sky130_fd_sc_hd__o22ai_2
X_17422_ svm0.delta\[12\] _09320_ net668 VGND VGND VPWR VPWR _09323_ sky130_fd_sc_hd__o21a_1
XFILLER_0_135_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length7471 net7472 VGND VGND VPWR VPWR net7471 sky130_fd_sc_hd__clkbuf_1
X_14634_ _06799_ VGND VGND VPWR VPWR _00123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17353_ net6658 net771 svm0.rising VGND VGND VPWR VPWR _09267_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_51_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14565_ _06737_ _06740_ _06741_ VGND VGND VPWR VPWR _06742_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16304_ _08366_ _08367_ _08241_ VGND VGND VPWR VPWR _08368_ sky130_fd_sc_hd__mux2_1
X_13516_ net7770 net1942 net2291 VGND VGND VPWR VPWR _05787_ sky130_fd_sc_hd__and3_1
X_17284_ svm0.counter\[8\] svm0.counter\[11\] svm0.counter\[10\] net6693 VGND VGND
+ VPWR VPWR _09199_ sky130_fd_sc_hd__or4_1
XFILLER_0_126_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14496_ _06673_ _06675_ _06678_ VGND VGND VPWR VPWR _06679_ sky130_fd_sc_hd__a21o_1
X_19023_ net1759 _10859_ VGND VGND VPWR VPWR _10860_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_181_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16235_ _08297_ _08299_ VGND VGND VPWR VPWR _08300_ sky130_fd_sc_hd__xor2_1
X_13447_ _05520_ _05522_ VGND VGND VPWR VPWR _05720_ sky130_fd_sc_hd__or2_1
XFILLER_0_140_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13378_ _05636_ _05650_ VGND VGND VPWR VPWR _05651_ sky130_fd_sc_hd__xor2_1
X_16166_ _08150_ _08155_ _08153_ VGND VGND VPWR VPWR _08232_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15117_ net3462 net2760 VGND VGND VPWR VPWR _07191_ sky130_fd_sc_hd__nor2_1
X_16097_ net2699 net2727 net1260 VGND VGND VPWR VPWR _08163_ sky130_fd_sc_hd__a21o_1
Xfanout4594 pid_q.mult0.a\[9\] VGND VGND VPWR VPWR net4594 sky130_fd_sc_hd__buf_1
Xwire5390 net5388 VGND VGND VPWR VPWR net5390 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_103_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19925_ _11377_ _11756_ net6174 VGND VGND VPWR VPWR _11757_ sky130_fd_sc_hd__mux2_1
X_15048_ _07111_ _07115_ _07121_ VGND VGND VPWR VPWR _07122_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19856_ _11687_ _11688_ VGND VGND VPWR VPWR _11689_ sky130_fd_sc_hd__nand2_1
X_18807_ _10649_ _10650_ VGND VGND VPWR VPWR _10651_ sky130_fd_sc_hd__xor2_1
X_19787_ net568 net488 _11620_ VGND VGND VPWR VPWR _11621_ sky130_fd_sc_hd__a21oi_1
X_16999_ _08923_ _08936_ _08938_ net7113 VGND VGND VPWR VPWR _08961_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18738_ net3231 net6826 VGND VGND VPWR VPWR _10583_ sky130_fd_sc_hd__and2_1
XFILLER_0_183_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18669_ net714 _10513_ _10514_ _10457_ VGND VGND VPWR VPWR _10515_ sky130_fd_sc_hd__o22a_1
X_20700_ _12463_ _12464_ _08993_ VGND VGND VPWR VPWR _12474_ sky130_fd_sc_hd__o21ai_1
X_21680_ net5842 net5413 VGND VGND VPWR VPWR _01691_ sky130_fd_sc_hd__nand2_1
X_20631_ _12406_ _12410_ VGND VGND VPWR VPWR _12411_ sky130_fd_sc_hd__and2b_1
XFILLER_0_18_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4119 net4120 VGND VGND VPWR VPWR net4119 sky130_fd_sc_hd__clkbuf_1
Xwire7709 net7710 VGND VGND VPWR VPWR net7709 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_178_Right_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23350_ _03218_ _03219_ VGND VGND VPWR VPWR _03220_ sky130_fd_sc_hd__xnor2_1
X_20562_ net1237 _12345_ net2516 VGND VGND VPWR VPWR _12347_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22301_ net5762 _02228_ VGND VGND VPWR VPWR _02305_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23281_ _03104_ _03112_ _03150_ VGND VGND VPWR VPWR _03151_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20493_ net3169 net1499 VGND VGND VPWR VPWR _12281_ sky130_fd_sc_hd__nand2_1
X_25020_ _03578_ _04768_ _04773_ VGND VGND VPWR VPWR _04774_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22232_ _02207_ _02236_ VGND VGND VPWR VPWR _02237_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22163_ _02116_ _02168_ VGND VGND VPWR VPWR _02169_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21114_ _01126_ _01129_ VGND VGND VPWR VPWR _01130_ sky130_fd_sc_hd__or2b_1
X_22094_ _02100_ _02010_ pid_d.prev_error\[8\] VGND VGND VPWR VPWR _02101_ sky130_fd_sc_hd__o21ba_1
Xwire2005 net2006 VGND VGND VPWR VPWR net2005 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2016 net2017 VGND VGND VPWR VPWR net2016 sky130_fd_sc_hd__buf_1
XFILLER_0_121_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2027 _02870_ VGND VGND VPWR VPWR net2027 sky130_fd_sc_hd__buf_1
X_25922_ clknet_leaf_96_clk _00795_ net8412 VGND VGND VPWR VPWR pid_d.prev_int\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_21045_ net2075 net2074 net2480 VGND VGND VPWR VPWR _01061_ sky130_fd_sc_hd__a21o_1
Xwire1304 _06374_ VGND VGND VPWR VPWR net1304 sky130_fd_sc_hd__clkbuf_2
Xwire2049 _02521_ VGND VGND VPWR VPWR net2049 sky130_fd_sc_hd__buf_1
Xwire1315 net1316 VGND VGND VPWR VPWR net1315 sky130_fd_sc_hd__buf_1
XFILLER_0_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1326 net1327 VGND VGND VPWR VPWR net1326 sky130_fd_sc_hd__buf_1
X_25853_ clknet_leaf_38_clk _00726_ net8745 VGND VGND VPWR VPWR pid_q.mult0.b\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1348 net1349 VGND VGND VPWR VPWR net1348 sky130_fd_sc_hd__clkbuf_1
Xwire1359 _04735_ VGND VGND VPWR VPWR net1359 sky130_fd_sc_hd__buf_1
X_24804_ net7961 _04620_ _04626_ _04627_ VGND VGND VPWR VPWR _04628_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25784_ clknet_leaf_57_clk _00657_ net8709 VGND VGND VPWR VPWR matmul0.beta_pass\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_22996_ net7470 pid_q.state\[0\] net7489 net8865 VGND VGND VPWR VPWR _02866_ sky130_fd_sc_hd__o31a_1
XFILLER_0_119_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24735_ net8007 net4272 VGND VGND VPWR VPWR _04568_ sky130_fd_sc_hd__xor2_1
XFILLER_0_179_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21947_ net5839 net5394 net5406 VGND VGND VPWR VPWR _01955_ sky130_fd_sc_hd__or3b_1
X_12680_ _04949_ _04952_ VGND VGND VPWR VPWR _04953_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_16_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24666_ net9139 net1375 _04515_ VGND VGND VPWR VPWR _00685_ sky130_fd_sc_hd__a21o_1
X_21878_ net2064 VGND VGND VPWR VPWR _01887_ sky130_fd_sc_hd__buf_1
XFILLER_0_49_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23617_ pid_q.curr_int\[3\] pid_q.prev_int\[3\] VGND VGND VPWR VPWR _03484_ sky130_fd_sc_hd__xor2_1
X_20829_ _12560_ _12561_ _12562_ VGND VGND VPWR VPWR _00845_ sky130_fd_sc_hd__o21a_1
Xwire8911 net8912 VGND VGND VPWR VPWR net8911 sky130_fd_sc_hd__buf_1
Xwire8922 net8923 VGND VGND VPWR VPWR net8922 sky130_fd_sc_hd__clkbuf_1
X_24597_ _09581_ _04452_ VGND VGND VPWR VPWR _04453_ sky130_fd_sc_hd__nor2_1
Xmax_length5354 pid_d.out\[9\] VGND VGND VPWR VPWR net5354 sky130_fd_sc_hd__buf_1
Xwire8933 net8934 VGND VGND VPWR VPWR net8933 sky130_fd_sc_hd__clkbuf_1
Xwire8944 net8945 VGND VGND VPWR VPWR net8944 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_145_Right_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14350_ _06564_ matmul0.a_in\[7\] net903 VGND VGND VPWR VPWR _06565_ sky130_fd_sc_hd__mux2_1
X_23548_ _03337_ _03338_ _03339_ VGND VGND VPWR VPWR _03416_ sky130_fd_sc_hd__o21a_1
Xwire601 net602 VGND VGND VPWR VPWR net601 sky130_fd_sc_hd__clkbuf_1
Xwire612 _09282_ VGND VGND VPWR VPWR net612 sky130_fd_sc_hd__buf_1
XFILLER_0_107_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire623 net624 VGND VGND VPWR VPWR net623 sky130_fd_sc_hd__clkbuf_1
X_13301_ net1135 _05499_ VGND VGND VPWR VPWR _05574_ sky130_fd_sc_hd__or2b_1
Xwire634 net635 VGND VGND VPWR VPWR net634 sky130_fd_sc_hd__clkbuf_2
X_14281_ net72 net2902 net2265 net7914 VGND VGND VPWR VPWR _00052_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23479_ _03336_ _03347_ VGND VGND VPWR VPWR _03348_ sky130_fd_sc_hd__xnor2_1
Xwire645 _03238_ VGND VGND VPWR VPWR net645 sky130_fd_sc_hd__clkbuf_1
Xwire656 _11368_ VGND VGND VPWR VPWR net656 sky130_fd_sc_hd__clkbuf_1
Xmax_length3963 _09795_ VGND VGND VPWR VPWR net3963 sky130_fd_sc_hd__buf_1
Xwire667 net668 VGND VGND VPWR VPWR net667 sky130_fd_sc_hd__buf_1
XFILLER_0_134_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire678 _06079_ VGND VGND VPWR VPWR net678 sky130_fd_sc_hd__clkbuf_1
X_13232_ net7755 _05504_ VGND VGND VPWR VPWR _05505_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16020_ _08087_ VGND VGND VPWR VPWR _00221_ sky130_fd_sc_hd__clkbuf_1
Xwire689 _04650_ VGND VGND VPWR VPWR net689 sky130_fd_sc_hd__clkbuf_1
X_25218_ clknet_leaf_59_clk _00107_ net8689 VGND VGND VPWR VPWR svm0.vC\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length265 _04388_ VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__clkbuf_1
X_13163_ _05374_ _05375_ VGND VGND VPWR VPWR _05436_ sky130_fd_sc_hd__and2_1
X_25149_ clknet_leaf_44_clk _00038_ net8781 VGND VGND VPWR VPWR pid_q.target\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13094_ net7672 net2339 net1967 VGND VGND VPWR VPWR _05367_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17971_ _09820_ _09821_ VGND VGND VPWR VPWR _09822_ sky130_fd_sc_hd__or2b_1
X_19710_ _11544_ _11545_ VGND VGND VPWR VPWR _11546_ sky130_fd_sc_hd__nor2_1
X_16922_ cordic0.slte0.opA\[1\] cordic0.slte0.opA\[0\] cordic0.slte0.opA\[2\] VGND
+ VGND VPWR VPWR _08886_ sky130_fd_sc_hd__o21ai_1
Xwire3251 net3252 VGND VGND VPWR VPWR net3251 sky130_fd_sc_hd__clkbuf_1
Xwire3273 net3274 VGND VGND VPWR VPWR net3273 sky130_fd_sc_hd__buf_1
Xwire2550 _09865_ VGND VGND VPWR VPWR net2550 sky130_fd_sc_hd__clkbuf_2
X_19641_ _11405_ _11476_ _11477_ VGND VGND VPWR VPWR _11478_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16853_ _08817_ VGND VGND VPWR VPWR _08818_ sky130_fd_sc_hd__clkbuf_1
Xwire2561 _09677_ VGND VGND VPWR VPWR net2561 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2572 net2573 VGND VGND VPWR VPWR net2572 sky130_fd_sc_hd__buf_1
Xwire2583 net2584 VGND VGND VPWR VPWR net2583 sky130_fd_sc_hd__buf_1
Xwire2594 _09069_ VGND VGND VPWR VPWR net2594 sky130_fd_sc_hd__buf_1
XFILLER_0_172_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1860 _07537_ VGND VGND VPWR VPWR net1860 sky130_fd_sc_hd__buf_1
X_15804_ net2693 net3465 VGND VGND VPWR VPWR _07874_ sky130_fd_sc_hd__nor2_1
X_19572_ _10790_ VGND VGND VPWR VPWR _11409_ sky130_fd_sc_hd__buf_1
Xwire1871 _07385_ VGND VGND VPWR VPWR net1871 sky130_fd_sc_hd__clkbuf_1
X_16784_ net7592 matmul0.a\[11\] net3373 VGND VGND VPWR VPWR _08782_ sky130_fd_sc_hd__mux2_1
X_13996_ _06169_ _06170_ VGND VGND VPWR VPWR _06261_ sky130_fd_sc_hd__and2b_1
Xwire1882 _07271_ VGND VGND VPWR VPWR net1882 sky130_fd_sc_hd__buf_1
XFILLER_0_88_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1893 _07188_ VGND VGND VPWR VPWR net1893 sky130_fd_sc_hd__clkbuf_2
X_18523_ net3285 net6793 VGND VGND VPWR VPWR _10372_ sky130_fd_sc_hd__nand2_2
XFILLER_0_153_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15735_ net2250 _07720_ _07717_ VGND VGND VPWR VPWR _07806_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_158_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12947_ net7940 net7917 net1350 _05216_ _05219_ VGND VGND VPWR VPWR _05220_ sky130_fd_sc_hd__a41o_1
XFILLER_0_172_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18454_ _10302_ _10303_ VGND VGND VPWR VPWR _10304_ sky130_fd_sc_hd__nor2_2
X_15666_ net574 _07642_ _07637_ VGND VGND VPWR VPWR _07738_ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12878_ _05079_ _05083_ _05143_ _05088_ VGND VGND VPWR VPWR _05151_ sky130_fd_sc_hd__o22a_1
XFILLER_0_185_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17405_ net613 _09309_ _09307_ VGND VGND VPWR VPWR _09310_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14617_ _06787_ _06788_ VGND VGND VPWR VPWR _06789_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18385_ _10234_ _10235_ net7012 VGND VGND VPWR VPWR _10236_ sky130_fd_sc_hd__a21o_1
X_15597_ net1109 _07623_ _07668_ VGND VGND VPWR VPWR _07669_ sky130_fd_sc_hd__o21a_1
X_17336_ _09210_ _09229_ _09234_ _09235_ _09249_ VGND VGND VPWR VPWR _09250_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_172_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14548_ _06711_ _06717_ VGND VGND VPWR VPWR _06726_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_112_Right_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17267_ net2160 net223 net1797 svm0.tA\[3\] VGND VGND VPWR VPWR _00361_ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14479_ _06663_ _06664_ VGND VGND VPWR VPWR _06665_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19006_ _10842_ VGND VGND VPWR VPWR _10843_ sky130_fd_sc_hd__buf_1
XFILLER_0_102_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16218_ _08274_ _08282_ VGND VGND VPWR VPWR _08283_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17198_ net6850 net618 _09147_ net6841 _09129_ VGND VGND VPWR VPWR _09148_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16149_ net2662 _08114_ _08116_ VGND VGND VPWR VPWR _08215_ sky130_fd_sc_hd__o21a_1
XFILLER_0_80_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19908_ _11712_ _11714_ VGND VGND VPWR VPWR _11740_ sky130_fd_sc_hd__nor2_1
Xhold19 cordic0.cos\[9\] VGND VGND VPWR VPWR net8972 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19839_ net8968 net1200 _11672_ net1768 VGND VGND VPWR VPWR _00456_ sky130_fd_sc_hd__a22o_1
XFILLER_0_190_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22850_ _02747_ _02748_ VGND VGND VPWR VPWR _02749_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21801_ _01810_ _01730_ pid_d.prev_error\[5\] VGND VGND VPWR VPWR _01811_ sky130_fd_sc_hd__o21ba_1
X_22781_ _02698_ VGND VGND VPWR VPWR _00617_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24520_ net792 VGND VGND VPWR VPWR _04377_ sky130_fd_sc_hd__inv_2
X_21732_ _01654_ _01716_ _01741_ VGND VGND VPWR VPWR _01742_ sky130_fd_sc_hd__o21a_2
XFILLER_0_4_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24451_ _04270_ _04308_ VGND VGND VPWR VPWR _04309_ sky130_fd_sc_hd__xnor2_1
X_21663_ net5768 net5502 VGND VGND VPWR VPWR _01674_ sky130_fd_sc_hd__nand2_1
Xwire8207 net8208 VGND VGND VPWR VPWR net8207 sky130_fd_sc_hd__clkbuf_1
Xwire8218 net8219 VGND VGND VPWR VPWR net8218 sky130_fd_sc_hd__clkbuf_1
Xwire8229 net8230 VGND VGND VPWR VPWR net8229 sky130_fd_sc_hd__clkbuf_1
X_23402_ net5033 net4614 VGND VGND VPWR VPWR _03272_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20614_ net3854 net3852 net2594 VGND VGND VPWR VPWR _12395_ sky130_fd_sc_hd__mux2_1
Xwire7506 net7501 VGND VGND VPWR VPWR net7506 sky130_fd_sc_hd__buf_1
X_24382_ _04153_ _04157_ _04158_ VGND VGND VPWR VPWR _04241_ sky130_fd_sc_hd__a21bo_1
Xwire7517 net7518 VGND VGND VPWR VPWR net7517 sky130_fd_sc_hd__clkbuf_1
Xmax_length3204 net3205 VGND VGND VPWR VPWR net3204 sky130_fd_sc_hd__clkbuf_1
X_21594_ net5892 net5400 VGND VGND VPWR VPWR _01606_ sky130_fd_sc_hd__nand2_1
Xwire7528 net7529 VGND VGND VPWR VPWR net7528 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23333_ net5162 net4540 VGND VGND VPWR VPWR _03203_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_104_Left_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire7539 net7540 VGND VGND VPWR VPWR net7539 sky130_fd_sc_hd__clkbuf_1
X_20545_ net2084 _12329_ net6310 VGND VGND VPWR VPWR _12330_ sky130_fd_sc_hd__a21o_1
Xwire6805 net6803 VGND VGND VPWR VPWR net6805 sky130_fd_sc_hd__clkbuf_1
Xwire6827 net6825 VGND VGND VPWR VPWR net6827 sky130_fd_sc_hd__buf_1
Xwire6838 net6834 VGND VGND VPWR VPWR net6838 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire6849 net6843 VGND VGND VPWR VPWR net6849 sky130_fd_sc_hd__buf_1
X_23264_ net4983 net4776 _03032_ VGND VGND VPWR VPWR _03134_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20476_ net7056 net7010 net7042 net6983 net6489 net6512 VGND VGND VPWR VPWR _12265_
+ sky130_fd_sc_hd__mux4_1
X_22215_ _02214_ _02219_ VGND VGND VPWR VPWR _02220_ sky130_fd_sc_hd__xnor2_1
X_25003_ pid_q.out\[1\] net1631 net2394 _04759_ VGND VGND VPWR VPWR _00778_ sky130_fd_sc_hd__a22o_1
X_23195_ net4757 net4777 VGND VGND VPWR VPWR _03065_ sky130_fd_sc_hd__and2_1
X_22146_ net5380 _02151_ VGND VGND VPWR VPWR _02152_ sky130_fd_sc_hd__nand2_2
XFILLER_0_30_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22077_ _01974_ _02082_ _02083_ _01978_ VGND VGND VPWR VPWR _02084_ sky130_fd_sc_hd__o22ai_2
Xwire1101 net1102 VGND VGND VPWR VPWR net1101 sky130_fd_sc_hd__clkbuf_1
X_25905_ clknet_leaf_65_clk _00778_ net8703 VGND VGND VPWR VPWR pid_q.out\[1\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_113_Left_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21028_ _00987_ _00988_ VGND VGND VPWR VPWR _01044_ sky130_fd_sc_hd__xnor2_1
Xwire1112 _07612_ VGND VGND VPWR VPWR net1112 sky130_fd_sc_hd__clkbuf_1
Xwire1123 _06326_ VGND VGND VPWR VPWR net1123 sky130_fd_sc_hd__clkbuf_2
Xwire1134 _05513_ VGND VGND VPWR VPWR net1134 sky130_fd_sc_hd__clkbuf_1
Xwire1145 net1146 VGND VGND VPWR VPWR net1145 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1156 _05023_ VGND VGND VPWR VPWR net1156 sky130_fd_sc_hd__clkbuf_1
Xwire1167 _03295_ VGND VGND VPWR VPWR net1167 sky130_fd_sc_hd__buf_1
X_13850_ net7633 VGND VGND VPWR VPWR _06117_ sky130_fd_sc_hd__inv_2
X_25836_ clknet_leaf_31_clk _00709_ net8685 VGND VGND VPWR VPWR pid_q.curr_error\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1178 _01583_ VGND VGND VPWR VPWR net1178 sky130_fd_sc_hd__buf_1
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1189 net1190 VGND VGND VPWR VPWR net1189 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12801_ _05073_ VGND VGND VPWR VPWR _05074_ sky130_fd_sc_hd__inv_2
X_13781_ net841 _06048_ VGND VGND VPWR VPWR _06049_ sky130_fd_sc_hd__xnor2_1
X_25767_ clknet_leaf_27_clk _00640_ net8646 VGND VGND VPWR VPWR pid_d.out\[8\] sky130_fd_sc_hd__dfrtp_1
X_22979_ _02857_ VGND VGND VPWR VPWR _00656_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15520_ net3497 net3600 VGND VGND VPWR VPWR _07593_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24718_ net8017 net4268 VGND VGND VPWR VPWR _04553_ sky130_fd_sc_hd__xor2_1
X_12732_ net7882 net1974 net1971 VGND VGND VPWR VPWR _05005_ sky130_fd_sc_hd__and3_1
Xfanout8602 net8607 VGND VGND VPWR VPWR net8602 sky130_fd_sc_hd__buf_1
X_25698_ clknet_leaf_120_clk _00571_ net8395 VGND VGND VPWR VPWR pid_d.mult0.b\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15451_ net1539 net1869 _07524_ VGND VGND VPWR VPWR _07525_ sky130_fd_sc_hd__o21a_1
X_24649_ net3731 _04503_ VGND VGND VPWR VPWR _04504_ sky130_fd_sc_hd__xnor2_1
X_12663_ net7813 _04924_ _04926_ VGND VGND VPWR VPWR _04936_ sky130_fd_sc_hd__and3_1
XFILLER_0_84_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14402_ net5289 net1298 net2892 net4458 _06604_ VGND VGND VPWR VPWR _06605_ sky130_fd_sc_hd__a221o_1
XFILLER_0_194_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout7934 net7942 VGND VGND VPWR VPWR net7934 sky130_fd_sc_hd__clkbuf_1
X_18170_ _09777_ _09778_ _09779_ _09673_ VGND VGND VPWR VPWR _10021_ sky130_fd_sc_hd__o31a_1
Xwire8741 net8742 VGND VGND VPWR VPWR net8741 sky130_fd_sc_hd__clkbuf_1
X_15382_ net1878 net1275 _07313_ VGND VGND VPWR VPWR _07456_ sky130_fd_sc_hd__a21o_1
X_12594_ _04865_ net4293 VGND VGND VPWR VPWR _00005_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17121_ _09064_ _09076_ VGND VGND VPWR VPWR _09077_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8774 net8775 VGND VGND VPWR VPWR net8774 sky130_fd_sc_hd__clkbuf_1
Xwire420 _11926_ VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__buf_1
X_14333_ net7332 net1299 net2896 pid_d.out\[3\] _06551_ VGND VGND VPWR VPWR _06552_
+ sky130_fd_sc_hd__a221o_1
Xwire8785 net8784 VGND VGND VPWR VPWR net8785 sky130_fd_sc_hd__clkbuf_2
Xwire431 net432 VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__clkbuf_1
Xwire8796 net8792 VGND VGND VPWR VPWR net8796 sky130_fd_sc_hd__buf_1
Xwire442 net443 VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__clkbuf_1
Xmax_length4494 net4495 VGND VGND VPWR VPWR net4494 sky130_fd_sc_hd__clkbuf_1
Xwire453 net454 VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire464 net465 VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__clkbuf_1
X_17052_ net1805 _08975_ net2172 net1807 VGND VGND VPWR VPWR _09011_ sky130_fd_sc_hd__o31a_1
X_14264_ net57 net2931 net2278 net9023 VGND VGND VPWR VPWR _00037_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire475 net476 VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire486 _01242_ VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__clkbuf_1
Xwire497 net498 VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__clkbuf_1
X_16003_ _07973_ _08069_ _08070_ VGND VGND VPWR VPWR _08071_ sky130_fd_sc_hd__a21oi_1
X_13215_ net7690 net1340 VGND VGND VPWR VPWR _05488_ sky130_fd_sc_hd__nand2_1
X_14195_ _06451_ _06416_ _06452_ _06453_ _06454_ VGND VGND VPWR VPWR _06455_ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13146_ net7215 net3029 _04894_ VGND VGND VPWR VPWR _05419_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13077_ _05290_ _05296_ _05287_ VGND VGND VPWR VPWR _05350_ sky130_fd_sc_hd__o21ai_1
X_17954_ net2552 _09803_ _09804_ VGND VGND VPWR VPWR _09805_ sky130_fd_sc_hd__or3_1
Xwire3070 net3071 VGND VGND VPWR VPWR net3070 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire3081 _02600_ VGND VGND VPWR VPWR net3081 sky130_fd_sc_hd__dlymetal6s2s_1
X_16905_ _08862_ net6371 VGND VGND VPWR VPWR _08869_ sky130_fd_sc_hd__nor2_1
Xwire3092 _02552_ VGND VGND VPWR VPWR net3092 sky130_fd_sc_hd__buf_1
X_17885_ net6994 net6947 VGND VGND VPWR VPWR _09736_ sky130_fd_sc_hd__nand2_1
Xwire2380 net2381 VGND VGND VPWR VPWR net2380 sky130_fd_sc_hd__buf_1
XFILLER_0_164_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2391 _04852_ VGND VGND VPWR VPWR net2391 sky130_fd_sc_hd__buf_1
X_19624_ _11459_ _11460_ net6221 VGND VGND VPWR VPWR _11461_ sky130_fd_sc_hd__a21o_1
X_16836_ net9245 matmul0.sin\[6\] net3366 VGND VGND VPWR VPWR _08809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1690 net1691 VGND VGND VPWR VPWR net1690 sky130_fd_sc_hd__buf_1
X_19555_ net3177 _10938_ _11324_ VGND VGND VPWR VPWR _11392_ sky130_fd_sc_hd__mux2_1
X_16767_ net9158 matmul0.a\[3\] net3378 VGND VGND VPWR VPWR _08773_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13979_ _06234_ _06243_ VGND VGND VPWR VPWR _06244_ sky130_fd_sc_hd__xnor2_1
X_18506_ net3928 _10288_ _10354_ VGND VGND VPWR VPWR _10355_ sky130_fd_sc_hd__a21oi_1
X_15718_ net2799 net3392 VGND VGND VPWR VPWR _07789_ sky130_fd_sc_hd__nor2_1
X_19486_ _11262_ _11263_ net6272 VGND VGND VPWR VPWR _11323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16698_ _08727_ VGND VGND VPWR VPWR _00259_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18437_ net6956 _10285_ _10286_ net3933 VGND VGND VPWR VPWR _10287_ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15649_ net2250 net2666 _07717_ VGND VGND VPWR VPWR _07721_ sky130_fd_sc_hd__or3_1
XFILLER_0_111_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18368_ _10169_ net3924 VGND VGND VPWR VPWR _10219_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17319_ _09209_ _09231_ _09232_ VGND VGND VPWR VPWR _09233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18299_ net815 _10147_ _10137_ _10149_ VGND VGND VPWR VPWR _10150_ sky130_fd_sc_hd__or4b_1
Xclkbuf_leaf_122_clk clknet_4_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_122_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_113_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20330_ net2607 _08990_ VGND VGND VPWR VPWR _12133_ sky130_fd_sc_hd__nand2_2
XFILLER_0_98_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_189_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20261_ net8121 _12072_ VGND VGND VPWR VPWR _12073_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22000_ pid_d.curr_error\[7\] VGND VGND VPWR VPWR _02008_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20192_ net1770 _12016_ _12017_ VGND VGND VPWR VPWR _00464_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput109 pid_d_data[6] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_1
X_23951_ _03681_ _03683_ _03814_ VGND VGND VPWR VPWR _03815_ sky130_fd_sc_hd__a21oi_2
Xmax_length8705 net8706 VGND VGND VPWR VPWR net8705 sky130_fd_sc_hd__clkbuf_1
Xmax_length8716 net8712 VGND VGND VPWR VPWR net8716 sky130_fd_sc_hd__buf_1
X_22902_ pid_d.out\[10\] net3103 VGND VGND VPWR VPWR _02795_ sky130_fd_sc_hd__nor2_1
X_23882_ _03736_ _03746_ VGND VGND VPWR VPWR _03747_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length8749 net8750 VGND VGND VPWR VPWR net8749 sky130_fd_sc_hd__clkbuf_1
X_25621_ clknet_leaf_116_clk _00494_ net8329 VGND VGND VPWR VPWR cordic0.slte0.opA\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_22833_ net5983 VGND VGND VPWR VPWR _02733_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25552_ clknet_leaf_79_clk net6592 net8490 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_22764_ _02687_ VGND VGND VPWR VPWR _00611_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_177_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24503_ _04296_ net4551 net2406 net4539 VGND VGND VPWR VPWR _04360_ sky130_fd_sc_hd__or4b_1
XFILLER_0_164_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21715_ _01724_ _01725_ VGND VGND VPWR VPWR _01726_ sky130_fd_sc_hd__and2b_1
X_25483_ clknet_leaf_45_clk _00363_ net8787 VGND VGND VPWR VPWR svm0.tA\[5\] sky130_fd_sc_hd__dfrtp_1
X_22695_ _02638_ VGND VGND VPWR VPWR _00591_ sky130_fd_sc_hd__clkbuf_1
Xwire8004 net8005 VGND VGND VPWR VPWR net8004 sky130_fd_sc_hd__clkbuf_1
Xwire8015 net8016 VGND VGND VPWR VPWR net8015 sky130_fd_sc_hd__clkbuf_1
Xwire8026 net8027 VGND VGND VPWR VPWR net8026 sky130_fd_sc_hd__clkbuf_1
Xwire8037 net8038 VGND VGND VPWR VPWR net8037 sky130_fd_sc_hd__clkbuf_1
X_24434_ net4872 net3745 net3753 VGND VGND VPWR VPWR _04292_ sky130_fd_sc_hd__a21o_1
X_21646_ _01556_ _01566_ _01561_ VGND VGND VPWR VPWR _01657_ sky130_fd_sc_hd__a21bo_1
Xwire7303 net7304 VGND VGND VPWR VPWR net7303 sky130_fd_sc_hd__buf_1
Xwire8048 net8049 VGND VGND VPWR VPWR net8048 sky130_fd_sc_hd__buf_1
Xwire7314 net7315 VGND VGND VPWR VPWR net7314 sky130_fd_sc_hd__buf_1
Xwire8059 net8061 VGND VGND VPWR VPWR net8059 sky130_fd_sc_hd__clkbuf_1
Xwire7325 net7326 VGND VGND VPWR VPWR net7325 sky130_fd_sc_hd__buf_1
Xwire7336 net7337 VGND VGND VPWR VPWR net7336 sky130_fd_sc_hd__dlymetal6s2s_1
X_24365_ net3041 _04223_ VGND VGND VPWR VPWR _04224_ sky130_fd_sc_hd__xnor2_1
Xwire6602 net6603 VGND VGND VPWR VPWR net6602 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21577_ _01585_ _01588_ VGND VGND VPWR VPWR _01589_ sky130_fd_sc_hd__xnor2_2
Xclkbuf_leaf_113_clk clknet_4_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_113_clk
+ sky130_fd_sc_hd__clkbuf_16
Xwire7347 net7348 VGND VGND VPWR VPWR net7347 sky130_fd_sc_hd__clkbuf_1
Xwire7358 net7359 VGND VGND VPWR VPWR net7358 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7369 net7370 VGND VGND VPWR VPWR net7369 sky130_fd_sc_hd__buf_1
X_23316_ net4864 net4760 VGND VGND VPWR VPWR _03186_ sky130_fd_sc_hd__nand2_1
Xfanout5839 net5848 VGND VGND VPWR VPWR net5839 sky130_fd_sc_hd__clkbuf_2
X_20528_ net6983 net6938 net6962 net6923 net6490 net6513 VGND VGND VPWR VPWR _12314_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_160_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24296_ net4803 _04056_ _04154_ VGND VGND VPWR VPWR _04156_ sky130_fd_sc_hd__a21o_1
Xwire6646 net6647 VGND VGND VPWR VPWR net6646 sky130_fd_sc_hd__clkbuf_1
Xwire5901 net5902 VGND VGND VPWR VPWR net5901 sky130_fd_sc_hd__clkbuf_1
Xwire6657 net6659 VGND VGND VPWR VPWR net6657 sky130_fd_sc_hd__buf_1
XFILLER_0_162_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6668 net6669 VGND VGND VPWR VPWR net6668 sky130_fd_sc_hd__clkbuf_1
Xmax_length1610 _05015_ VGND VGND VPWR VPWR net1610 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire5923 net5924 VGND VGND VPWR VPWR net5923 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5934 net5931 VGND VGND VPWR VPWR net5934 sky130_fd_sc_hd__clkbuf_1
Xwire6679 net6680 VGND VGND VPWR VPWR net6679 sky130_fd_sc_hd__clkbuf_1
X_23247_ net4966 net4776 VGND VGND VPWR VPWR _03117_ sky130_fd_sc_hd__nand2_1
X_20459_ _12244_ net809 cordic0.slte0.opA\[14\] VGND VGND VPWR VPWR _12251_ sky130_fd_sc_hd__a21bo_1
Xwire5945 net5946 VGND VGND VPWR VPWR net5945 sky130_fd_sc_hd__buf_1
Xwire5956 net5957 VGND VGND VPWR VPWR net5956 sky130_fd_sc_hd__clkbuf_1
Xwire5967 pid_d.curr_error\[9\] VGND VGND VPWR VPWR net5967 sky130_fd_sc_hd__buf_1
Xmax_length1665 _03575_ VGND VGND VPWR VPWR net1665 sky130_fd_sc_hd__clkbuf_1
X_13000_ _05156_ _05157_ net7874 net1959 VGND VGND VPWR VPWR _05273_ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5978 pid_d.curr_int\[7\] VGND VGND VPWR VPWR net5978 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_162_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5989 net5990 VGND VGND VPWR VPWR net5989 sky130_fd_sc_hd__dlymetal6s2s_1
X_23178_ _03046_ _03047_ VGND VGND VPWR VPWR _03048_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22129_ _02126_ _02134_ VGND VGND VPWR VPWR _02135_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14951_ net6630 matmul0.matmul_stage_inst.d\[4\] net7414 net6532 VGND VGND VPWR VPWR
+ _07025_ sky130_fd_sc_hd__a22o_1
X_13902_ net7744 net1326 _06101_ _06100_ VGND VGND VPWR VPWR _06168_ sky130_fd_sc_hd__a31o_1
X_17670_ net4013 svm0.tA\[1\] VGND VGND VPWR VPWR _09550_ sky130_fd_sc_hd__nand2_1
X_14882_ net9237 matmul0.matmul_stage_inst.f\[13\] net3606 VGND VGND VPWR VPWR _06959_
+ sky130_fd_sc_hd__mux2_1
X_16621_ matmul0.matmul_stage_inst.mult2\[0\] matmul0.matmul_stage_inst.mult1\[0\]
+ VGND VGND VPWR VPWR _08661_ sky130_fd_sc_hd__nand2_1
X_13833_ net7766 net2948 net1940 VGND VGND VPWR VPWR _06100_ sky130_fd_sc_hd__and3_1
X_25819_ clknet_leaf_32_clk _00692_ net8685 VGND VGND VPWR VPWR pid_q.prev_error\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19340_ net6227 net6289 VGND VGND VPWR VPWR _11177_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16552_ _08562_ _08610_ VGND VGND VPWR VPWR _08611_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13764_ _06029_ _06030_ _06027_ VGND VGND VPWR VPWR _06032_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15503_ net2228 _07575_ VGND VGND VPWR VPWR _07576_ sky130_fd_sc_hd__xnor2_2
X_12715_ _04986_ _04987_ VGND VGND VPWR VPWR _04988_ sky130_fd_sc_hd__xor2_2
X_19271_ _11094_ _11096_ _11107_ VGND VGND VPWR VPWR _11108_ sky130_fd_sc_hd__and3b_1
Xfanout8410 net8418 VGND VGND VPWR VPWR net8410 sky130_fd_sc_hd__clkbuf_1
X_16483_ _08542_ _08543_ VGND VGND VPWR VPWR _08544_ sky130_fd_sc_hd__or2b_1
X_13695_ _05962_ _05963_ VGND VGND VPWR VPWR _05964_ sky130_fd_sc_hd__xnor2_1
Xfanout8432 net8522 VGND VGND VPWR VPWR net8432 sky130_fd_sc_hd__buf_1
XFILLER_0_31_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18222_ _10055_ _10072_ VGND VGND VPWR VPWR _10073_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_182_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15434_ net3510 net3505 net4210 net4208 VGND VGND VPWR VPWR _07508_ sky130_fd_sc_hd__o22a_1
X_12646_ net2353 net2348 VGND VGND VPWR VPWR _04919_ sky130_fd_sc_hd__and2_1
Xfanout8465 net8483 VGND VGND VPWR VPWR net8465 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8560 net8555 VGND VGND VPWR VPWR net8560 sky130_fd_sc_hd__clkbuf_2
X_18153_ _09751_ _09755_ VGND VGND VPWR VPWR _10004_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_104_clk clknet_4_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_104_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15365_ net2233 net2824 net2249 _07438_ VGND VGND VPWR VPWR _07439_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8582 net8583 VGND VGND VPWR VPWR net8582 sky130_fd_sc_hd__buf_1
XFILLER_0_4_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12577_ net6597 VGND VGND VPWR VPWR _04864_ sky130_fd_sc_hd__inv_2
Xfanout7786 net7793 VGND VGND VPWR VPWR net7786 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8593 net8594 VGND VGND VPWR VPWR net8593 sky130_fd_sc_hd__buf_1
X_17104_ _09039_ net772 net6981 VGND VGND VPWR VPWR _09061_ sky130_fd_sc_hd__a21o_1
X_14316_ clarke_done net2386 _06537_ VGND VGND VPWR VPWR _06538_ sky130_fd_sc_hd__o21a_1
Xwire250 net251 VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7870 net7871 VGND VGND VPWR VPWR net7870 sky130_fd_sc_hd__clkbuf_1
Xwire261 net262 VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__clkbuf_1
X_18084_ net7062 _09933_ net3940 VGND VGND VPWR VPWR _09935_ sky130_fd_sc_hd__o21a_1
Xwire272 net273 VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__buf_1
Xwire7881 net7882 VGND VGND VPWR VPWR net7881 sky130_fd_sc_hd__buf_1
X_15296_ net6631 matmul0.matmul_stage_inst.d\[12\] matmul0.matmul_stage_inst.c\[12\]
+ net6533 VGND VGND VPWR VPWR _07370_ sky130_fd_sc_hd__a22o_1
Xwire7892 net7893 VGND VGND VPWR VPWR net7892 sky130_fd_sc_hd__clkbuf_1
Xwire283 _06020_ VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3590 net3591 VGND VGND VPWR VPWR net3590 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire294 _02614_ VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__clkbuf_1
X_17035_ _08976_ _08980_ VGND VGND VPWR VPWR _08995_ sky130_fd_sc_hd__nor2_1
X_14247_ _06501_ VGND VGND VPWR VPWR _06502_ sky130_fd_sc_hd__buf_1
XFILLER_0_110_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14178_ _06434_ _06436_ _06437_ VGND VGND VPWR VPWR _06438_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13129_ net920 _05302_ VGND VGND VPWR VPWR _05402_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18986_ net6312 net6352 VGND VGND VPWR VPWR _10823_ sky130_fd_sc_hd__or2b_1
X_17937_ _09780_ _09787_ VGND VGND VPWR VPWR _09788_ sky130_fd_sc_hd__nand2_1
X_17868_ _09715_ _09716_ _09717_ _09718_ VGND VGND VPWR VPWR _09719_ sky130_fd_sc_hd__o22a_1
X_19607_ net6097 net6085 VGND VGND VPWR VPWR _11444_ sky130_fd_sc_hd__and2b_1
X_16819_ cordic0.cos\[12\] matmul0.cos\[12\] _08792_ VGND VGND VPWR VPWR _08800_ sky130_fd_sc_hd__mux2_1
X_17799_ net7104 net7119 net7091 VGND VGND VPWR VPWR _09650_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_191_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19538_ _11346_ net3155 _11374_ VGND VGND VPWR VPWR _11375_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_177_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19469_ net960 net1420 VGND VGND VPWR VPWR _11306_ sky130_fd_sc_hd__or2_1
XFILLER_0_192_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21500_ _01381_ _01382_ _01512_ VGND VGND VPWR VPWR _01513_ sky130_fd_sc_hd__a21oi_1
X_22480_ _02477_ _02480_ VGND VGND VPWR VPWR _02481_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21431_ _01403_ _01443_ VGND VGND VPWR VPWR _01444_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24150_ net4675 net3043 _03924_ VGND VGND VPWR VPWR _04012_ sky130_fd_sc_hd__or3b_1
XFILLER_0_140_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21362_ _01374_ _01375_ VGND VGND VPWR VPWR _01376_ sky130_fd_sc_hd__xnor2_1
Xwire5208 net5209 VGND VGND VPWR VPWR net5208 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23101_ _02969_ _02970_ VGND VGND VPWR VPWR _02971_ sky130_fd_sc_hd__nand2_1
X_20313_ net9187 _12116_ _12117_ VGND VGND VPWR VPWR _00485_ sky130_fd_sc_hd__a21bo_1
X_24081_ _03941_ _03943_ VGND VGND VPWR VPWR _03944_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput80 periodTop[9] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21293_ net3811 _12515_ _01307_ VGND VGND VPWR VPWR _01308_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_102_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput91 pid_d_addr[4] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_1
Xwire4518 net4519 VGND VGND VPWR VPWR net4518 sky130_fd_sc_hd__clkbuf_1
Xwire4529 net4531 VGND VGND VPWR VPWR net4529 sky130_fd_sc_hd__clkbuf_1
X_23032_ _02900_ _02901_ VGND VGND VPWR VPWR _02902_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20244_ _12059_ cordic0.slte0.opB\[9\] net2532 VGND VGND VPWR VPWR _12060_ sky130_fd_sc_hd__mux2_1
Xwire3806 _01054_ VGND VGND VPWR VPWR net3806 sky130_fd_sc_hd__buf_1
Xwire3817 net3818 VGND VGND VPWR VPWR net3817 sky130_fd_sc_hd__clkbuf_1
Xwire3828 _00960_ VGND VGND VPWR VPWR net3828 sky130_fd_sc_hd__clkbuf_1
Xwire3839 _00881_ VGND VGND VPWR VPWR net3839 sky130_fd_sc_hd__buf_1
XFILLER_0_149_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20175_ net6059 net6100 net2580 net6024 VGND VGND VPWR VPWR _12001_ sky130_fd_sc_hd__or4_1
X_24983_ _04746_ VGND VGND VPWR VPWR _00771_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23934_ _03715_ _03720_ _03713_ VGND VGND VPWR VPWR _03798_ sky130_fd_sc_hd__o21a_1
XFILLER_0_192_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length7801 net7802 VGND VGND VPWR VPWR net7801 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23865_ _03727_ _03729_ VGND VGND VPWR VPWR _03730_ sky130_fd_sc_hd__nand2_1
XFILLER_0_168_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25604_ clknet_leaf_108_clk _00477_ net8344 VGND VGND VPWR VPWR cordic0.slte0.opB\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_22816_ _02718_ net4336 VGND VGND VPWR VPWR _02719_ sky130_fd_sc_hd__and2b_1
XFILLER_0_79_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23796_ pid_q.prev_error\[3\] VGND VGND VPWR VPWR _03662_ sky130_fd_sc_hd__inv_2
XFILLER_0_196_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25535_ clknet_4_12__leaf_clk _00415_ net8695 VGND VGND VPWR VPWR pid_q.prev_int\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22747_ net3719 net110 VGND VGND VPWR VPWR _02676_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25466_ clknet_leaf_52_clk _00346_ net8807 VGND VGND VPWR VPWR svm0.tB\[4\] sky130_fd_sc_hd__dfrtp_1
X_13480_ _05751_ _05752_ VGND VGND VPWR VPWR _05753_ sky130_fd_sc_hd__xor2_1
Xfanout7027 net7031 VGND VGND VPWR VPWR net7027 sky130_fd_sc_hd__buf_2
X_22678_ pid_d.ki\[3\] net2439 net2994 pid_d.kp\[3\] VGND VGND VPWR VPWR _02627_ sky130_fd_sc_hd__a22o_1
Xwire7100 net7101 VGND VGND VPWR VPWR net7100 sky130_fd_sc_hd__clkbuf_1
X_24417_ net4798 _04209_ _04273_ VGND VGND VPWR VPWR _04275_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21629_ _01638_ _01639_ VGND VGND VPWR VPWR _01641_ sky130_fd_sc_hd__or2_1
Xfanout6337 net6341 VGND VGND VPWR VPWR net6337 sky130_fd_sc_hd__clkbuf_1
Xwire7133 net7131 VGND VGND VPWR VPWR net7133 sky130_fd_sc_hd__clkbuf_4
X_25397_ clknet_leaf_71_clk _00280_ net8461 VGND VGND VPWR VPWR matmul0.a\[0\] sky130_fd_sc_hd__dfrtp_1
Xwire7144 net7145 VGND VGND VPWR VPWR net7144 sky130_fd_sc_hd__buf_1
Xfanout5614 net5619 VGND VGND VPWR VPWR net5614 sky130_fd_sc_hd__clkbuf_1
Xwire6410 net6411 VGND VGND VPWR VPWR net6410 sky130_fd_sc_hd__buf_1
Xwire7155 matmul0.sin\[5\] VGND VGND VPWR VPWR net7155 sky130_fd_sc_hd__buf_1
Xfanout5625 net5629 VGND VGND VPWR VPWR net5625 sky130_fd_sc_hd__buf_1
X_15150_ net2757 _07142_ VGND VGND VPWR VPWR _07224_ sky130_fd_sc_hd__nor2_1
Xwire7166 matmul0.cos\[13\] VGND VGND VPWR VPWR net7166 sky130_fd_sc_hd__buf_1
Xwire6421 cordic0.sin\[11\] VGND VGND VPWR VPWR net6421 sky130_fd_sc_hd__clkbuf_1
X_24348_ net4536 net4857 VGND VGND VPWR VPWR _04207_ sky130_fd_sc_hd__nand2_1
Xwire7177 matmul0.cos\[7\] VGND VGND VPWR VPWR net7177 sky130_fd_sc_hd__clkbuf_1
Xwire6432 net6433 VGND VGND VPWR VPWR net6432 sky130_fd_sc_hd__buf_1
Xfanout5636 net5643 VGND VGND VPWR VPWR net5636 sky130_fd_sc_hd__buf_1
Xwire7188 net7189 VGND VGND VPWR VPWR net7188 sky130_fd_sc_hd__clkbuf_1
X_14101_ net9112 _05780_ net188 net2374 VGND VGND VPWR VPWR _00026_ sky130_fd_sc_hd__a22o_1
Xwire7199 net7200 VGND VGND VPWR VPWR net7199 sky130_fd_sc_hd__buf_1
Xwire6454 net6452 VGND VGND VPWR VPWR net6454 sky130_fd_sc_hd__clkbuf_2
Xwire5720 net5721 VGND VGND VPWR VPWR net5720 sky130_fd_sc_hd__buf_1
Xfanout5669 net5678 VGND VGND VPWR VPWR net5669 sky130_fd_sc_hd__buf_1
XFILLER_0_121_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6465 net6463 VGND VGND VPWR VPWR net6465 sky130_fd_sc_hd__buf_1
Xwire5731 net5724 VGND VGND VPWR VPWR net5731 sky130_fd_sc_hd__buf_1
X_15081_ net2781 net2795 _07145_ net3489 VGND VGND VPWR VPWR _07155_ sky130_fd_sc_hd__and4_1
X_24279_ _04081_ _04083_ _04138_ VGND VGND VPWR VPWR _04139_ sky130_fd_sc_hd__o21ai_1
Xwire5742 net5743 VGND VGND VPWR VPWR net5742 sky130_fd_sc_hd__clkbuf_1
Xwire6487 cordic0.gm0.iter\[2\] VGND VGND VPWR VPWR net6487 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5753 net5754 VGND VGND VPWR VPWR net5753 sky130_fd_sc_hd__buf_1
Xmax_length1451 net1452 VGND VGND VPWR VPWR net1451 sky130_fd_sc_hd__buf_1
X_14032_ net7642 _05608_ _05609_ VGND VGND VPWR VPWR _06296_ sky130_fd_sc_hd__and3_1
Xwire5764 net5762 VGND VGND VPWR VPWR net5764 sky130_fd_sc_hd__buf_1
Xwire5786 net5787 VGND VGND VPWR VPWR net5786 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5797 net5795 VGND VGND VPWR VPWR net5797 sky130_fd_sc_hd__buf_1
X_18840_ _10641_ _10349_ VGND VGND VPWR VPWR _10683_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18771_ _10603_ _10615_ VGND VGND VPWR VPWR _10616_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15983_ net2762 _07932_ net3444 VGND VGND VPWR VPWR _08051_ sky130_fd_sc_hd__or3b_1
X_17722_ net9125 net1456 net1789 net5173 VGND VGND VPWR VPWR _00427_ sky130_fd_sc_hd__a22o_1
X_14934_ net2256 _07007_ VGND VGND VPWR VPWR _07008_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_54_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17653_ _09525_ _09526_ _09527_ _09532_ VGND VGND VPWR VPWR _09533_ sky130_fd_sc_hd__or4_1
X_14865_ net4284 VGND VGND VPWR VPWR _06950_ sky130_fd_sc_hd__buf_1
X_16604_ matmul0.matmul_stage_inst.mult2\[9\] net305 net2618 VGND VGND VPWR VPWR _08652_
+ sky130_fd_sc_hd__mux2_1
X_13816_ net532 _06083_ VGND VGND VPWR VPWR _06084_ sky130_fd_sc_hd__xor2_1
X_17584_ svm0.tC\[11\] _09439_ _09465_ VGND VGND VPWR VPWR _09466_ sky130_fd_sc_hd__o21a_1
X_14796_ net7438 net7181 net2856 VGND VGND VPWR VPWR _06915_ sky130_fd_sc_hd__a21o_1
XFILLER_0_159_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19323_ net2107 _11159_ VGND VGND VPWR VPWR _11160_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_175_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16535_ _08522_ net880 VGND VGND VPWR VPWR _08594_ sky130_fd_sc_hd__nand2_1
X_13747_ _05866_ _05868_ net404 VGND VGND VPWR VPWR _06015_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19254_ net1753 _11089_ VGND VGND VPWR VPWR _11091_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16466_ net2625 net2209 VGND VGND VPWR VPWR _08527_ sky130_fd_sc_hd__nand2_1
X_13678_ net7768 net3670 VGND VGND VPWR VPWR _05947_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18205_ net2139 _09805_ _09806_ _09812_ VGND VGND VPWR VPWR _10056_ sky130_fd_sc_hd__a31o_1
X_15417_ _07487_ _07490_ VGND VGND VPWR VPWR _07491_ sky130_fd_sc_hd__nor2_1
X_12629_ net1618 VGND VGND VPWR VPWR _04902_ sky130_fd_sc_hd__clkbuf_1
X_19185_ net1064 _11021_ VGND VGND VPWR VPWR _11022_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16397_ net2783 _08455_ _08456_ _08458_ net2744 VGND VGND VPWR VPWR _08459_ sky130_fd_sc_hd__o32a_1
XFILLER_0_53_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18136_ _09914_ _09923_ _09929_ VGND VGND VPWR VPWR _09987_ sky130_fd_sc_hd__a21o_1
Xwire8390 net8391 VGND VGND VPWR VPWR net8390 sky130_fd_sc_hd__clkbuf_2
X_15348_ net2726 net2782 net2704 VGND VGND VPWR VPWR _07422_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold105 svm0.vC\[5\] VGND VGND VPWR VPWR net9058 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18067_ net7041 net7112 net7134 VGND VGND VPWR VPWR _09918_ sky130_fd_sc_hd__and3_1
XFILLER_0_124_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15279_ net4095 net4094 VGND VGND VPWR VPWR _07353_ sky130_fd_sc_hd__nor2_1
Xhold116 matmul0.matmul_stage_inst.d\[2\] VGND VGND VPWR VPWR net9069 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 svm0.tB\[9\] VGND VGND VPWR VPWR net9080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 svm0.tC\[14\] VGND VGND VPWR VPWR net9091 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 cordic0.in_valid VGND VGND VPWR VPWR net9102 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17018_ net7086 _08959_ VGND VGND VPWR VPWR _08979_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18969_ net2530 net3214 VGND VGND VPWR VPWR _10806_ sky130_fd_sc_hd__or2_1
X_21980_ net1717 _01878_ VGND VGND VPWR VPWR _01988_ sky130_fd_sc_hd__xnor2_1
Xmax_length7108 net7109 VGND VGND VPWR VPWR net7108 sky130_fd_sc_hd__clkbuf_2
X_20931_ _00945_ _00946_ VGND VGND VPWR VPWR _00947_ sky130_fd_sc_hd__nand2_1
Xmax_length7119 net7121 VGND VGND VPWR VPWR net7119 sky130_fd_sc_hd__buf_1
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23650_ net3748 _03395_ _03394_ VGND VGND VPWR VPWR _03517_ sky130_fd_sc_hd__o21ai_1
X_20862_ net5642 net5740 VGND VGND VPWR VPWR _00878_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22601_ net7265 _02574_ VGND VGND VPWR VPWR _02576_ sky130_fd_sc_hd__or2_2
X_23581_ _03423_ _03448_ VGND VGND VPWR VPWR _03449_ sky130_fd_sc_hd__xnor2_2
X_20793_ _12560_ _12563_ VGND VGND VPWR VPWR _00809_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_159_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25320_ clknet_leaf_75_clk _00203_ net8463 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.f\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22532_ net9106 net1699 _02528_ VGND VGND VPWR VPWR _00538_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25251_ clknet_leaf_88_clk _00134_ net8431 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.a\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22463_ pid_d.curr_int\[15\] pid_d.prev_int\[15\] VGND VGND VPWR VPWR _02464_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24202_ net4535 net4890 VGND VGND VPWR VPWR _04063_ sky130_fd_sc_hd__nand2_1
X_21414_ pid_d.prev_error\[1\] net5972 VGND VGND VPWR VPWR _01428_ sky130_fd_sc_hd__or2_1
X_22394_ pid_d.curr_int\[13\] net3844 net2488 _02396_ VGND VGND VPWR VPWR _00532_
+ sky130_fd_sc_hd__a22o_1
X_25182_ clknet_leaf_68_clk _00071_ net8450 VGND VGND VPWR VPWR matmul0.a_in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire5005 net5006 VGND VGND VPWR VPWR net5005 sky130_fd_sc_hd__buf_1
Xwire5016 net5017 VGND VGND VPWR VPWR net5016 sky130_fd_sc_hd__buf_1
XFILLER_0_161_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5027 net5028 VGND VGND VPWR VPWR net5027 sky130_fd_sc_hd__buf_1
X_24133_ _03878_ _03883_ _03876_ VGND VGND VPWR VPWR _03995_ sky130_fd_sc_hd__o21a_1
XFILLER_0_114_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21345_ _01292_ _01297_ VGND VGND VPWR VPWR _01359_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5038 net5039 VGND VGND VPWR VPWR net5038 sky130_fd_sc_hd__buf_1
Xwire5049 net5050 VGND VGND VPWR VPWR net5049 sky130_fd_sc_hd__clkbuf_1
Xwire4304 net4305 VGND VGND VPWR VPWR net4304 sky130_fd_sc_hd__clkbuf_1
Xwire4315 net4316 VGND VGND VPWR VPWR net4315 sky130_fd_sc_hd__buf_1
X_24064_ _03925_ _03926_ net4675 VGND VGND VPWR VPWR _03927_ sky130_fd_sc_hd__mux2_1
Xwire4337 net4338 VGND VGND VPWR VPWR net4337 sky130_fd_sc_hd__buf_1
X_21276_ net5687 net5626 VGND VGND VPWR VPWR _01291_ sky130_fd_sc_hd__nand2_1
Xwire4348 net4349 VGND VGND VPWR VPWR net4348 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3614 net3615 VGND VGND VPWR VPWR net3614 sky130_fd_sc_hd__buf_1
X_23015_ _02881_ _02882_ _02884_ VGND VGND VPWR VPWR _02885_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20227_ _12046_ VGND VGND VPWR VPWR _00470_ sky130_fd_sc_hd__clkbuf_1
Xwire3625 _06818_ VGND VGND VPWR VPWR net3625 sky130_fd_sc_hd__buf_1
XFILLER_0_102_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3636 _06575_ VGND VGND VPWR VPWR net3636 sky130_fd_sc_hd__buf_1
Xwire2902 net2903 VGND VGND VPWR VPWR net2902 sky130_fd_sc_hd__clkbuf_2
Xwire3647 net3648 VGND VGND VPWR VPWR net3647 sky130_fd_sc_hd__buf_1
Xwire2913 _06516_ VGND VGND VPWR VPWR net2913 sky130_fd_sc_hd__clkbuf_1
Xwire3658 net3659 VGND VGND VPWR VPWR net3658 sky130_fd_sc_hd__buf_1
Xwire2924 net2925 VGND VGND VPWR VPWR net2924 sky130_fd_sc_hd__clkbuf_1
Xwire3669 net3670 VGND VGND VPWR VPWR net3669 sky130_fd_sc_hd__buf_1
X_20158_ _11984_ _11980_ VGND VGND VPWR VPWR _11985_ sky130_fd_sc_hd__or2_1
Xwire2946 net2947 VGND VGND VPWR VPWR net2946 sky130_fd_sc_hd__buf_1
Xwire2957 net2958 VGND VGND VPWR VPWR net2957 sky130_fd_sc_hd__clkbuf_1
Xwire2968 net2969 VGND VGND VPWR VPWR net2968 sky130_fd_sc_hd__buf_1
Xwire2979 net2980 VGND VGND VPWR VPWR net2979 sky130_fd_sc_hd__clkbuf_1
X_24966_ pid_q.kp\[2\] _04706_ net1357 VGND VGND VPWR VPWR _04738_ sky130_fd_sc_hd__mux2_1
X_12980_ _05249_ _05252_ VGND VGND VPWR VPWR _05253_ sky130_fd_sc_hd__xnor2_2
X_20089_ _11914_ _11916_ _11917_ _11846_ net3861 VGND VGND VPWR VPWR _11918_ sky130_fd_sc_hd__a221oi_1
X_23917_ _03731_ _03732_ _03780_ VGND VGND VPWR VPWR _03781_ sky130_fd_sc_hd__o21a_1
X_24897_ _04689_ VGND VGND VPWR VPWR _00742_ sky130_fd_sc_hd__clkbuf_1
X_14650_ net8989 net2880 _06809_ VGND VGND VPWR VPWR _00129_ sky130_fd_sc_hd__a21o_1
X_23848_ _03711_ _03712_ VGND VGND VPWR VPWR _03713_ sky130_fd_sc_hd__xor2_2
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length7653 net7654 VGND VGND VPWR VPWR net7653 sky130_fd_sc_hd__buf_1
XFILLER_0_79_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13601_ _05784_ net533 VGND VGND VPWR VPWR _05871_ sky130_fd_sc_hd__nor2_1
Xmax_length6930 net6923 VGND VGND VPWR VPWR net6930 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14581_ _06752_ _06756_ VGND VGND VPWR VPWR _06757_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_184_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23779_ net4796 net3049 VGND VGND VPWR VPWR _03645_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16320_ net2721 net2707 net2648 _08258_ VGND VGND VPWR VPWR _08383_ sky130_fd_sc_hd__a211o_1
X_25518_ clknet_leaf_44_clk _00398_ net8785 VGND VGND VPWR VPWR svm0.counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13532_ _05799_ _05800_ _05801_ _05802_ VGND VGND VPWR VPWR _05803_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_82_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16251_ net2220 _08279_ _08312_ net2651 net3492 VGND VGND VPWR VPWR _08315_ sky130_fd_sc_hd__o221a_1
X_13463_ net7705 net1151 _05585_ _05586_ VGND VGND VPWR VPWR _05736_ sky130_fd_sc_hd__a22o_1
X_25449_ clknet_leaf_119_clk _00332_ net8338 VGND VGND VPWR VPWR cordic0.vec\[1\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15202_ net2238 _07087_ _07272_ _07273_ VGND VGND VPWR VPWR _07276_ sky130_fd_sc_hd__a22o_1
Xfanout6156 net6159 VGND VGND VPWR VPWR net6156 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16182_ net774 _08246_ _08207_ VGND VGND VPWR VPWR _08247_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_180_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13394_ net583 _05663_ net581 VGND VGND VPWR VPWR _05667_ sky130_fd_sc_hd__nand3_1
Xwire6251 net6252 VGND VGND VPWR VPWR net6251 sky130_fd_sc_hd__buf_1
X_15133_ net3481 VGND VGND VPWR VPWR _07207_ sky130_fd_sc_hd__clkbuf_1
Xwire6262 net6261 VGND VGND VPWR VPWR net6262 sky130_fd_sc_hd__buf_1
Xfanout4721 net4732 VGND VGND VPWR VPWR net4721 sky130_fd_sc_hd__clkbuf_1
Xwire6273 net6274 VGND VGND VPWR VPWR net6273 sky130_fd_sc_hd__buf_1
Xwire6284 net6285 VGND VGND VPWR VPWR net6284 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5550 net5551 VGND VGND VPWR VPWR net5550 sky130_fd_sc_hd__buf_1
Xwire5561 net5562 VGND VGND VPWR VPWR net5561 sky130_fd_sc_hd__clkbuf_1
X_15064_ net3488 VGND VGND VPWR VPWR _07138_ sky130_fd_sc_hd__clkbuf_1
X_19941_ net6033 net2501 _11699_ net6044 VGND VGND VPWR VPWR _11773_ sky130_fd_sc_hd__a2bb2o_1
Xwire5572 net5573 VGND VGND VPWR VPWR net5572 sky130_fd_sc_hd__buf_1
XFILLER_0_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout4787 pid_q.mult0.b\[15\] VGND VGND VPWR VPWR net4787 sky130_fd_sc_hd__buf_1
Xwire5583 net5584 VGND VGND VPWR VPWR net5583 sky130_fd_sc_hd__buf_1
X_14015_ _06278_ _06263_ net529 VGND VGND VPWR VPWR _06279_ sky130_fd_sc_hd__a21o_1
Xfanout4798 net4817 VGND VGND VPWR VPWR net4798 sky130_fd_sc_hd__buf_1
Xwire5594 net5586 VGND VGND VPWR VPWR net5594 sky130_fd_sc_hd__clkbuf_1
Xwire4860 net4861 VGND VGND VPWR VPWR net4860 sky130_fd_sc_hd__clkbuf_1
X_19872_ _11677_ _11704_ VGND VGND VPWR VPWR _11705_ sky130_fd_sc_hd__xnor2_1
Xwire4882 net4883 VGND VGND VPWR VPWR net4882 sky130_fd_sc_hd__clkbuf_1
Xwire4893 net4885 VGND VGND VPWR VPWR net4893 sky130_fd_sc_hd__clkbuf_1
X_18823_ _10636_ _10645_ _10644_ VGND VGND VPWR VPWR _10666_ sky130_fd_sc_hd__a21o_1
X_15966_ _07970_ net1522 _08033_ VGND VGND VPWR VPWR _08034_ sky130_fd_sc_hd__a21o_1
X_18754_ _10596_ _10598_ VGND VGND VPWR VPWR _10599_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_175_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17705_ net7496 VGND VGND VPWR VPWR _09581_ sky130_fd_sc_hd__inv_2
X_14917_ _06981_ _06986_ _06990_ VGND VGND VPWR VPWR _06991_ sky130_fd_sc_hd__o21a_1
XFILLER_0_175_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15897_ _07964_ _07965_ VGND VGND VPWR VPWR _07966_ sky130_fd_sc_hd__xor2_1
X_18685_ net6838 net3287 VGND VGND VPWR VPWR _10531_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_159_Right_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17636_ svm0.tB\[15\] _09472_ _09516_ VGND VGND VPWR VPWR _09517_ sky130_fd_sc_hd__o21a_1
XFILLER_0_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14848_ _06941_ VGND VGND VPWR VPWR _00195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17567_ net6706 _09442_ VGND VGND VPWR VPWR _09449_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14779_ net2866 _06903_ net9116 net3001 VGND VGND VPWR VPWR _00164_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_147_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19306_ net6312 net6352 _11142_ net6262 VGND VGND VPWR VPWR _11143_ sky130_fd_sc_hd__o211a_1
X_16518_ net3420 _08574_ _08576_ _08577_ VGND VGND VPWR VPWR _08578_ sky130_fd_sc_hd__a211o_1
X_17498_ net6705 _09385_ _09386_ _09384_ VGND VGND VPWR VPWR _00400_ sky130_fd_sc_hd__a22o_1
XFILLER_0_162_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19237_ _11071_ _11073_ net3198 VGND VGND VPWR VPWR _11074_ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16449_ _08505_ net1246 net1245 VGND VGND VPWR VPWR _08510_ sky130_fd_sc_hd__o21a_1
XFILLER_0_54_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19168_ _10940_ _11003_ _11004_ VGND VGND VPWR VPWR _11005_ sky130_fd_sc_hd__a21o_1
XFILLER_0_182_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18119_ _09968_ _09969_ VGND VGND VPWR VPWR _09970_ sky130_fd_sc_hd__and2b_1
XFILLER_0_124_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout6690 svm0.counter\[13\] VGND VGND VPWR VPWR net6690 sky130_fd_sc_hd__buf_1
X_19099_ _10922_ _10935_ VGND VGND VPWR VPWR _10936_ sky130_fd_sc_hd__or2b_1
XFILLER_0_30_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21130_ _01104_ _01111_ _01110_ VGND VGND VPWR VPWR _01146_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21061_ net1185 _01024_ VGND VGND VPWR VPWR _01077_ sky130_fd_sc_hd__xor2_1
Xwire2209 net2210 VGND VGND VPWR VPWR net2209 sky130_fd_sc_hd__buf_1
X_20012_ _11823_ _11836_ VGND VGND VPWR VPWR _11842_ sky130_fd_sc_hd__nor2_1
Xwire1508 _08254_ VGND VGND VPWR VPWR net1508 sky130_fd_sc_hd__buf_1
Xwire1519 _08045_ VGND VGND VPWR VPWR net1519 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24820_ net2008 VGND VGND VPWR VPWR _04642_ sky130_fd_sc_hd__buf_2
XFILLER_0_154_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24751_ _04580_ _04581_ VGND VGND VPWR VPWR _04582_ sky130_fd_sc_hd__nand2_1
X_21963_ _01845_ _01856_ _01970_ VGND VGND VPWR VPWR _01971_ sky130_fd_sc_hd__o21a_1
XFILLER_0_146_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_93_clk clknet_4_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_93_clk sky130_fd_sc_hd__clkbuf_16
X_23702_ pid_q.prev_error\[2\] VGND VGND VPWR VPWR _03569_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_126_Right_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20914_ _00926_ net1392 net1187 VGND VGND VPWR VPWR _00930_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_169_Left_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24682_ net9032 net1647 _04523_ VGND VGND VPWR VPWR _00693_ sky130_fd_sc_hd__a21o_1
XFILLER_0_178_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21894_ _01893_ _01902_ VGND VGND VPWR VPWR _01903_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23633_ net4748 net4812 VGND VGND VPWR VPWR _03500_ sky130_fd_sc_hd__nand2_1
Xmax_length6237 net6238 VGND VGND VPWR VPWR net6237 sky130_fd_sc_hd__clkbuf_1
X_20845_ _12520_ _12547_ _12535_ VGND VGND VPWR VPWR _00861_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_65_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23564_ _03350_ _03352_ _03431_ VGND VGND VPWR VPWR _03432_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_37_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length5558 net5559 VGND VGND VPWR VPWR net5558 sky130_fd_sc_hd__buf_1
X_20776_ _12541_ _12546_ VGND VGND VPWR VPWR _12547_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length4835 net4836 VGND VGND VPWR VPWR net4835 sky130_fd_sc_hd__buf_1
X_25303_ clknet_leaf_70_clk _00186_ net8459 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.e\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_193_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22515_ _02514_ _02515_ _02411_ VGND VGND VPWR VPWR _02516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23495_ _03245_ _03252_ _03251_ VGND VGND VPWR VPWR _03364_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire816 _10146_ VGND VGND VPWR VPWR net816 sky130_fd_sc_hd__clkbuf_1
Xwire827 net828 VGND VGND VPWR VPWR net827 sky130_fd_sc_hd__clkbuf_2
Xwire838 _06114_ VGND VGND VPWR VPWR net838 sky130_fd_sc_hd__clkbuf_1
X_25234_ clknet_leaf_23_clk _00007_ net8582 VGND VGND VPWR VPWR pid_q.state\[1\] sky130_fd_sc_hd__dfrtp_1
X_22446_ _02443_ _02447_ VGND VGND VPWR VPWR _02448_ sky130_fd_sc_hd__xor2_1
Xwire849 _05395_ VGND VGND VPWR VPWR net849 sky130_fd_sc_hd__buf_1
XFILLER_0_44_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25165_ clknet_leaf_54_clk _00054_ net8730 VGND VGND VPWR VPWR svm0.periodTop\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_178_Left_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22377_ _02341_ _02379_ VGND VGND VPWR VPWR _02380_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4101 net4102 VGND VGND VPWR VPWR net4101 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_102_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24116_ _03885_ _03888_ _03977_ VGND VGND VPWR VPWR _03978_ sky130_fd_sc_hd__a21o_1
XFILLER_0_130_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4112 net4113 VGND VGND VPWR VPWR net4112 sky130_fd_sc_hd__clkbuf_1
X_21328_ net759 _01253_ _01328_ _01329_ VGND VGND VPWR VPWR _01342_ sky130_fd_sc_hd__o31ai_2
X_25096_ _04836_ _04839_ VGND VGND VPWR VPWR _04840_ sky130_fd_sc_hd__xnor2_1
Xwire4123 _07088_ VGND VGND VPWR VPWR net4123 sky130_fd_sc_hd__buf_1
Xwire4134 _07030_ VGND VGND VPWR VPWR net4134 sky130_fd_sc_hd__clkbuf_1
Xwire3400 _07603_ VGND VGND VPWR VPWR net3400 sky130_fd_sc_hd__buf_1
Xwire4145 _07022_ VGND VGND VPWR VPWR net4145 sky130_fd_sc_hd__clkbuf_1
Xwire3411 net3412 VGND VGND VPWR VPWR net3411 sky130_fd_sc_hd__buf_1
Xwire4156 net4157 VGND VGND VPWR VPWR net4156 sky130_fd_sc_hd__buf_1
X_24047_ _03813_ _03815_ _03811_ VGND VGND VPWR VPWR _03910_ sky130_fd_sc_hd__a21bo_1
Xwire3422 _07511_ VGND VGND VPWR VPWR net3422 sky130_fd_sc_hd__buf_1
Xwire4167 net4168 VGND VGND VPWR VPWR net4167 sky130_fd_sc_hd__buf_1
X_21259_ _00825_ _00830_ _01273_ VGND VGND VPWR VPWR _01274_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3433 _07378_ VGND VGND VPWR VPWR net3433 sky130_fd_sc_hd__clkbuf_1
Xwire4178 _06997_ VGND VGND VPWR VPWR net4178 sky130_fd_sc_hd__buf_1
Xwire3444 _07245_ VGND VGND VPWR VPWR net3444 sky130_fd_sc_hd__buf_1
Xwire4189 _06993_ VGND VGND VPWR VPWR net4189 sky130_fd_sc_hd__clkbuf_1
Xwire3455 net3456 VGND VGND VPWR VPWR net3455 sky130_fd_sc_hd__buf_1
Xwire3466 _07157_ VGND VGND VPWR VPWR net3466 sky130_fd_sc_hd__buf_1
Xwire2721 net2722 VGND VGND VPWR VPWR net2721 sky130_fd_sc_hd__clkbuf_2
Xwire3477 _07151_ VGND VGND VPWR VPWR net3477 sky130_fd_sc_hd__clkbuf_1
Xwire2743 _07207_ VGND VGND VPWR VPWR net2743 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15820_ net827 _07889_ VGND VGND VPWR VPWR _07890_ sky130_fd_sc_hd__xnor2_2
Xwire3499 net3500 VGND VGND VPWR VPWR net3499 sky130_fd_sc_hd__clkbuf_2
Xwire2765 net2766 VGND VGND VPWR VPWR net2765 sky130_fd_sc_hd__buf_1
Xwire2787 net2788 VGND VGND VPWR VPWR net2787 sky130_fd_sc_hd__clkbuf_1
X_15751_ _07819_ _07821_ VGND VGND VPWR VPWR _07822_ sky130_fd_sc_hd__xnor2_1
X_24949_ pid_q.ki\[12\] _04726_ net1636 VGND VGND VPWR VPWR _04727_ sky130_fd_sc_hd__mux2_1
X_12963_ _05004_ net851 VGND VGND VPWR VPWR _05236_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_187_Left_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_84_clk clknet_4_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_84_clk sky130_fd_sc_hd__clkbuf_16
X_14702_ net9113 net2862 net2262 net1909 VGND VGND VPWR VPWR _00144_ sky130_fd_sc_hd__a22o_1
X_18470_ _10309_ _10318_ _10319_ _10315_ net6771 VGND VGND VPWR VPWR _10320_ sky130_fd_sc_hd__a311o_1
X_15682_ net3447 net3600 VGND VGND VPWR VPWR _07753_ sky130_fd_sc_hd__nor2_1
X_12894_ _05164_ _05165_ _05159_ VGND VGND VPWR VPWR _05167_ sky130_fd_sc_hd__a21oi_2
X_17421_ _09319_ net615 _09320_ _09322_ VGND VGND VPWR VPWR _00387_ sky130_fd_sc_hd__a31o_1
X_14633_ net7550 matmul0.op\[1\] net3704 VGND VGND VPWR VPWR _06799_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17352_ _09216_ _09256_ _09263_ _09265_ VGND VGND VPWR VPWR _09266_ sky130_fd_sc_hd__and4bb_1
X_14564_ net7244 net5213 VGND VGND VPWR VPWR _06741_ sky130_fd_sc_hd__xor2_2
XFILLER_0_67_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16303_ _08245_ _08365_ _08362_ VGND VGND VPWR VPWR _08367_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13515_ net7746 net2307 net1952 VGND VGND VPWR VPWR _05786_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17283_ net6732 net6716 net6708 net6745 VGND VGND VPWR VPWR _09198_ sky130_fd_sc_hd__or4_1
XFILLER_0_55_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14495_ _06673_ _06675_ _06674_ VGND VGND VPWR VPWR _06678_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_71_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19022_ net2527 _10858_ VGND VGND VPWR VPWR _10859_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16234_ net1088 net1511 _08298_ VGND VGND VPWR VPWR _08299_ sky130_fd_sc_hd__o21a_2
X_13446_ net7860 net1590 _05520_ _05522_ VGND VGND VPWR VPWR _05719_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_196_Left_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16165_ _08224_ _08230_ VGND VGND VPWR VPWR _08231_ sky130_fd_sc_hd__xnor2_1
X_13377_ _05538_ _05638_ _05644_ _05648_ _05649_ VGND VGND VPWR VPWR _05650_ sky130_fd_sc_hd__a311o_1
XFILLER_0_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6081 net6080 VGND VGND VPWR VPWR net6081 sky130_fd_sc_hd__clkbuf_2
X_15116_ net3597 net3591 VGND VGND VPWR VPWR _07190_ sky130_fd_sc_hd__nor2_1
Xfanout4540 net4550 VGND VGND VPWR VPWR net4540 sky130_fd_sc_hd__buf_1
Xfanout4551 net4565 VGND VGND VPWR VPWR net4551 sky130_fd_sc_hd__clkbuf_1
Xwire6092 net6091 VGND VGND VPWR VPWR net6092 sky130_fd_sc_hd__buf_1
X_16096_ _08162_ VGND VGND VPWR VPWR _00222_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19924_ net6111 net3200 VGND VGND VPWR VPWR _11756_ sky130_fd_sc_hd__nand2_1
X_15047_ _07111_ _07115_ _07120_ VGND VGND VPWR VPWR _07121_ sky130_fd_sc_hd__o21a_1
Xwire4690 net4691 VGND VGND VPWR VPWR net4690 sky130_fd_sc_hd__clkbuf_1
X_19855_ net6212 net6135 net6110 VGND VGND VPWR VPWR _11688_ sky130_fd_sc_hd__or3b_1
XFILLER_0_177_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18806_ net3221 net1760 VGND VGND VPWR VPWR _10650_ sky130_fd_sc_hd__nor2_1
X_19786_ net3859 VGND VGND VPWR VPWR _11620_ sky130_fd_sc_hd__buf_1
X_16998_ _08936_ _08938_ _08923_ VGND VGND VPWR VPWR _08960_ sky130_fd_sc_hd__a21o_1
X_18737_ net3231 net6826 VGND VGND VPWR VPWR _10582_ sky130_fd_sc_hd__nor2_1
X_15949_ _07958_ VGND VGND VPWR VPWR _08017_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_75_clk clknet_4_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_75_clk sky130_fd_sc_hd__clkbuf_16
X_18668_ net714 _10502_ VGND VGND VPWR VPWR _10514_ sky130_fd_sc_hd__nand2_1
X_17619_ net4012 svm0.tB\[1\] VGND VGND VPWR VPWR _09500_ sky130_fd_sc_hd__and2_1
X_18599_ net6860 _10369_ _10371_ net2129 VGND VGND VPWR VPWR _10447_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20630_ net1739 _12409_ VGND VGND VPWR VPWR _12410_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20561_ net2192 _12345_ VGND VGND VPWR VPWR _12346_ sky130_fd_sc_hd__or2_1
XFILLER_0_190_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22300_ _02283_ _02303_ VGND VGND VPWR VPWR _02304_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_41_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23280_ _03104_ _03112_ _03092_ VGND VGND VPWR VPWR _03150_ sky130_fd_sc_hd__o21a_1
X_20492_ net6363 net970 VGND VGND VPWR VPWR _12280_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length2718 net2719 VGND VGND VPWR VPWR net2718 sky130_fd_sc_hd__buf_1
Xmax_length2729 _07241_ VGND VGND VPWR VPWR net2729 sky130_fd_sc_hd__buf_1
XFILLER_0_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22231_ _02233_ net1033 VGND VGND VPWR VPWR _02236_ sky130_fd_sc_hd__xor2_1
XFILLER_0_48_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22162_ _02118_ _02167_ VGND VGND VPWR VPWR _02168_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_160_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21113_ _01127_ _01128_ VGND VGND VPWR VPWR _01129_ sky130_fd_sc_hd__xor2_2
XFILLER_0_140_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22093_ pid_d.curr_error\[8\] VGND VGND VPWR VPWR _02100_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2006 net2008 VGND VGND VPWR VPWR net2006 sky130_fd_sc_hd__clkbuf_1
Xwire2017 _04360_ VGND VGND VPWR VPWR net2017 sky130_fd_sc_hd__buf_1
X_25921_ clknet_leaf_97_clk _00794_ net8412 VGND VGND VPWR VPWR pid_d.prev_int\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_21044_ net2075 net2074 net1731 VGND VGND VPWR VPWR _01060_ sky130_fd_sc_hd__a21oi_1
Xwire2028 net2029 VGND VGND VPWR VPWR net2028 sky130_fd_sc_hd__buf_1
Xwire2039 _02661_ VGND VGND VPWR VPWR net2039 sky130_fd_sc_hd__buf_1
Xwire1305 _06245_ VGND VGND VPWR VPWR net1305 sky130_fd_sc_hd__buf_1
Xwire1316 _05687_ VGND VGND VPWR VPWR net1316 sky130_fd_sc_hd__buf_1
Xwire1327 net1328 VGND VGND VPWR VPWR net1327 sky130_fd_sc_hd__buf_1
XFILLER_0_157_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25852_ clknet_leaf_23_clk _00725_ net8586 VGND VGND VPWR VPWR pid_q.mult0.b\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1338 net1339 VGND VGND VPWR VPWR net1338 sky130_fd_sc_hd__clkbuf_2
Xwire1349 net1351 VGND VGND VPWR VPWR net1349 sky130_fd_sc_hd__clkbuf_1
X_24803_ _04618_ net7961 _06533_ _04619_ VGND VGND VPWR VPWR _04627_ sky130_fd_sc_hd__a211o_1
XFILLER_0_158_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25783_ clknet_leaf_73_clk _00656_ net8476 VGND VGND VPWR VPWR matmul0.beta_pass\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22995_ net6447 net6445 net9110 _02865_ VGND VGND VPWR VPWR _00664_ sky130_fd_sc_hd__o2bb2a_1
Xclkbuf_leaf_66_clk clknet_4_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_96_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24734_ _04565_ _04566_ VGND VGND VPWR VPWR _04567_ sky130_fd_sc_hd__and2_1
X_21946_ net1714 _01953_ VGND VGND VPWR VPWR _01954_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6023 net6018 VGND VGND VPWR VPWR net6023 sky130_fd_sc_hd__buf_1
XFILLER_0_189_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24665_ pid_q.curr_error\[4\] net2382 net1372 VGND VGND VPWR VPWR _04515_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21877_ net2066 _01788_ VGND VGND VPWR VPWR _01886_ sky130_fd_sc_hd__or2_1
Xmax_length6045 net6046 VGND VGND VPWR VPWR net6045 sky130_fd_sc_hd__buf_1
XFILLER_0_139_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6056 net6051 VGND VGND VPWR VPWR net6056 sky130_fd_sc_hd__clkbuf_1
X_23616_ pid_q.prev_int\[2\] _03391_ _03482_ VGND VGND VPWR VPWR _03483_ sky130_fd_sc_hd__o21ai_2
Xwire8901 net8902 VGND VGND VPWR VPWR net8901 sky130_fd_sc_hd__buf_1
Xmax_length6078 net6079 VGND VGND VPWR VPWR net6078 sky130_fd_sc_hd__buf_1
X_20828_ _00840_ _00843_ VGND VGND VPWR VPWR _00844_ sky130_fd_sc_hd__xnor2_2
X_24596_ _04448_ _04451_ VGND VGND VPWR VPWR _04452_ sky130_fd_sc_hd__xor2_1
Xwire8912 net8913 VGND VGND VPWR VPWR net8912 sky130_fd_sc_hd__clkbuf_1
Xmax_length6089 net6090 VGND VGND VPWR VPWR net6089 sky130_fd_sc_hd__clkbuf_1
Xwire8923 net113 VGND VGND VPWR VPWR net8923 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8934 net8935 VGND VGND VPWR VPWR net8934 sky130_fd_sc_hd__clkbuf_1
Xwire8945 net101 VGND VGND VPWR VPWR net8945 sky130_fd_sc_hd__clkbuf_1
X_23547_ _03411_ _03414_ VGND VGND VPWR VPWR _03415_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_21_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire602 _01552_ VGND VGND VPWR VPWR net602 sky130_fd_sc_hd__clkbuf_1
X_20759_ _12526_ _12529_ VGND VGND VPWR VPWR _12530_ sky130_fd_sc_hd__xnor2_1
Xmax_length4654 net4655 VGND VGND VPWR VPWR net4654 sky130_fd_sc_hd__buf_1
X_13300_ _05501_ _05515_ _05572_ VGND VGND VPWR VPWR _05573_ sky130_fd_sc_hd__o21a_1
XFILLER_0_52_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire624 _05760_ VGND VGND VPWR VPWR net624 sky130_fd_sc_hd__clkbuf_1
X_14280_ net65 net2902 net2265 net7934 VGND VGND VPWR VPWR _00051_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire635 _04166_ VGND VGND VPWR VPWR net635 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4687 net4680 VGND VGND VPWR VPWR net4687 sky130_fd_sc_hd__buf_1
X_23478_ _03341_ _03346_ VGND VGND VPWR VPWR _03347_ sky130_fd_sc_hd__xnor2_2
Xwire646 net647 VGND VGND VPWR VPWR net646 sky130_fd_sc_hd__buf_1
Xwire657 _10702_ VGND VGND VPWR VPWR net657 sky130_fd_sc_hd__buf_1
Xwire668 _09273_ VGND VGND VPWR VPWR net668 sky130_fd_sc_hd__buf_1
X_13231_ _04960_ VGND VGND VPWR VPWR _05504_ sky130_fd_sc_hd__clkbuf_1
X_25217_ clknet_leaf_59_clk _00106_ net8688 VGND VGND VPWR VPWR svm0.vC\[5\] sky130_fd_sc_hd__dfrtp_1
Xwire679 net680 VGND VGND VPWR VPWR net679 sky130_fd_sc_hd__buf_1
X_22429_ _02351_ _02356_ _02430_ VGND VGND VPWR VPWR _02431_ sky130_fd_sc_hd__o21a_1
XFILLER_0_21_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25148_ clknet_leaf_41_clk _00037_ net8767 VGND VGND VPWR VPWR pid_q.target\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13162_ _05383_ _05385_ VGND VGND VPWR VPWR _05435_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13093_ net7688 net1973 net1970 VGND VGND VPWR VPWR _05366_ sky130_fd_sc_hd__and3_1
X_25079_ net4406 net5174 VGND VGND VPWR VPWR _04825_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17970_ net6909 net6946 net6845 _09818_ _09819_ VGND VGND VPWR VPWR _09821_ sky130_fd_sc_hd__a311o_1
Xwire3230 _10063_ VGND VGND VPWR VPWR net3230 sky130_fd_sc_hd__clkbuf_1
Xwire3241 _09792_ VGND VGND VPWR VPWR net3241 sky130_fd_sc_hd__clkbuf_2
X_16921_ cordic0.slte0.opA\[3\] VGND VGND VPWR VPWR _08885_ sky130_fd_sc_hd__inv_2
Xwire3252 _09662_ VGND VGND VPWR VPWR net3252 sky130_fd_sc_hd__clkbuf_1
Xwire3274 _09332_ VGND VGND VPWR VPWR net3274 sky130_fd_sc_hd__buf_1
Xwire2540 _10276_ VGND VGND VPWR VPWR net2540 sky130_fd_sc_hd__buf_1
XFILLER_0_102_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2551 _09857_ VGND VGND VPWR VPWR net2551 sky130_fd_sc_hd__clkbuf_2
X_19640_ _11413_ _11415_ VGND VGND VPWR VPWR _11477_ sky130_fd_sc_hd__or2_1
Xwire3296 net3297 VGND VGND VPWR VPWR net3296 sky130_fd_sc_hd__buf_1
X_16852_ net6457 net3668 VGND VGND VPWR VPWR _08817_ sky130_fd_sc_hd__and2_1
Xwire2562 _09647_ VGND VGND VPWR VPWR net2562 sky130_fd_sc_hd__buf_1
Xwire2584 net2585 VGND VGND VPWR VPWR net2584 sky130_fd_sc_hd__clkbuf_1
Xwire2595 _09052_ VGND VGND VPWR VPWR net2595 sky130_fd_sc_hd__buf_1
Xwire1850 _07811_ VGND VGND VPWR VPWR net1850 sky130_fd_sc_hd__buf_1
X_15803_ net2647 net3481 VGND VGND VPWR VPWR _07873_ sky130_fd_sc_hd__nor2_1
X_19571_ net6012 _11348_ VGND VGND VPWR VPWR _11408_ sky130_fd_sc_hd__nand2_1
Xwire1861 net1862 VGND VGND VPWR VPWR net1861 sky130_fd_sc_hd__buf_1
X_16783_ net4289 VGND VGND VPWR VPWR _08781_ sky130_fd_sc_hd__clkbuf_1
X_13995_ _06172_ net677 _06259_ VGND VGND VPWR VPWR _06260_ sky130_fd_sc_hd__o21ai_2
Xwire1872 net1873 VGND VGND VPWR VPWR net1872 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_189_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_57_clk clknet_4_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_16
Xwire1883 _07249_ VGND VGND VPWR VPWR net1883 sky130_fd_sc_hd__buf_1
Xwire1894 _07171_ VGND VGND VPWR VPWR net1894 sky130_fd_sc_hd__clkbuf_2
X_15734_ net2661 _07717_ VGND VGND VPWR VPWR _07805_ sky130_fd_sc_hd__nor2_1
X_18522_ net6818 net3929 VGND VGND VPWR VPWR _10371_ sky130_fd_sc_hd__nand2_1
X_12946_ net7940 net7889 net1350 _05217_ _05218_ VGND VGND VPWR VPWR _05219_ sky130_fd_sc_hd__a41o_1
XFILLER_0_158_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15665_ net574 _07642_ _07736_ _07637_ VGND VGND VPWR VPWR _07737_ sky130_fd_sc_hd__a211o_1
X_18453_ net6933 net3331 VGND VGND VPWR VPWR _10303_ sky130_fd_sc_hd__nor2_1
X_12877_ _05079_ _05148_ _05149_ _05146_ VGND VGND VPWR VPWR _05150_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_29_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17404_ net2574 _09308_ VGND VGND VPWR VPWR _09309_ sky130_fd_sc_hd__or2_1
X_14616_ _06539_ _06786_ VGND VGND VPWR VPWR _06788_ sky130_fd_sc_hd__nand2_1
X_18384_ net3241 _10233_ VGND VGND VPWR VPWR _10235_ sky130_fd_sc_hd__or2_1
X_15596_ net1109 _07623_ net1270 VGND VGND VPWR VPWR _07668_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17335_ _09210_ _09229_ _09242_ _09248_ VGND VGND VPWR VPWR _09249_ sky130_fd_sc_hd__a211oi_1
Xmax_length6590 net6586 VGND VGND VPWR VPWR net6590 sky130_fd_sc_hd__clkbuf_1
X_14547_ _06711_ VGND VGND VPWR VPWR _06725_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17266_ net2160 net284 net1798 svm0.tA\[2\] VGND VGND VPWR VPWR _00360_ sky130_fd_sc_hd__a22o_1
X_14478_ _06658_ _06657_ _06659_ VGND VGND VPWR VPWR _06664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19005_ net6352 net6342 VGND VGND VPWR VPWR _10842_ sky130_fd_sc_hd__and2b_1
X_16217_ _08276_ _08281_ VGND VGND VPWR VPWR _08282_ sky130_fd_sc_hd__xor2_1
XFILLER_0_183_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13429_ net7792 net1942 net2291 VGND VGND VPWR VPWR _05702_ sky130_fd_sc_hd__and3_1
XFILLER_0_140_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17197_ net617 VGND VGND VPWR VPWR _09147_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16148_ net1093 net1092 _08213_ VGND VGND VPWR VPWR _08214_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_12_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16079_ net1517 net1256 VGND VGND VPWR VPWR _08146_ sky130_fd_sc_hd__xor2_1
X_19907_ _11738_ VGND VGND VPWR VPWR _11739_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19838_ _11621_ _11671_ VGND VGND VPWR VPWR _11672_ sky130_fd_sc_hd__xnor2_1
Xinput1 angle_in[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
X_19769_ net2502 _11494_ _11603_ VGND VGND VPWR VPWR _11604_ sky130_fd_sc_hd__o21ai_2
Xclkbuf_leaf_48_clk clknet_4_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21800_ net5969 VGND VGND VPWR VPWR _01810_ sky130_fd_sc_hd__inv_2
XFILLER_0_190_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22780_ pid_d.kp\[2\] _02666_ net1680 VGND VGND VPWR VPWR _02698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21731_ _01654_ _01716_ _01708_ VGND VGND VPWR VPWR _01741_ sky130_fd_sc_hd__a21o_1
X_24450_ _04279_ _04307_ VGND VGND VPWR VPWR _04308_ sky130_fd_sc_hd__xnor2_1
X_21662_ net5783 net5484 VGND VGND VPWR VPWR _01673_ sky130_fd_sc_hd__nand2_2
XFILLER_0_136_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8208 net8209 VGND VGND VPWR VPWR net8208 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8219 net8220 VGND VGND VPWR VPWR net8219 sky130_fd_sc_hd__clkbuf_1
X_23401_ _03201_ _03202_ _03270_ VGND VGND VPWR VPWR _03271_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_136_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20613_ net6766 net4038 _09055_ net3849 VGND VGND VPWR VPWR _12394_ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24381_ _04152_ _04160_ _04239_ VGND VGND VPWR VPWR _04240_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_149_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21593_ net1725 _01499_ _01604_ VGND VGND VPWR VPWR _01605_ sky130_fd_sc_hd__a21o_1
Xwire7518 net7519 VGND VGND VPWR VPWR net7518 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7529 pid_q.state\[1\] VGND VGND VPWR VPWR net7529 sky130_fd_sc_hd__clkbuf_1
X_23332_ net5124 net4568 VGND VGND VPWR VPWR _03202_ sky130_fd_sc_hd__nand2_1
X_20544_ net2079 VGND VGND VPWR VPWR _12329_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23263_ _03126_ _03132_ VGND VGND VPWR VPWR _03133_ sky130_fd_sc_hd__xnor2_1
Xmax_length2537 _10770_ VGND VGND VPWR VPWR net2537 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20475_ net6890 net6853 net6840 net6824 net6521 net6488 VGND VGND VPWR VPWR _12264_
+ sky130_fd_sc_hd__mux4_1
X_25002_ net7472 _04757_ _04758_ net7498 net538 VGND VGND VPWR VPWR _04759_ sky130_fd_sc_hd__a32o_1
X_22214_ _02215_ _02218_ VGND VGND VPWR VPWR _02219_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_14_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23194_ _03035_ _03063_ VGND VGND VPWR VPWR _03064_ sky130_fd_sc_hd__xnor2_1
X_22145_ net2065 _01964_ _02150_ net5817 VGND VGND VPWR VPWR _02151_ sky130_fd_sc_hd__a2bb2o_1
X_22076_ net2067 _01973_ VGND VGND VPWR VPWR _02083_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1102 net1103 VGND VGND VPWR VPWR net1102 sky130_fd_sc_hd__clkbuf_1
X_25904_ clknet_leaf_65_clk _00777_ net8654 VGND VGND VPWR VPWR pid_q.out\[0\] sky130_fd_sc_hd__dfrtp_1
X_21027_ net5631 net5820 VGND VGND VPWR VPWR _01043_ sky130_fd_sc_hd__nand2_1
Xwire1113 net1114 VGND VGND VPWR VPWR net1113 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_195_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1124 net1125 VGND VGND VPWR VPWR net1124 sky130_fd_sc_hd__buf_1
Xwire1135 _05494_ VGND VGND VPWR VPWR net1135 sky130_fd_sc_hd__buf_1
Xwire1146 _05066_ VGND VGND VPWR VPWR net1146 sky130_fd_sc_hd__clkbuf_1
X_25835_ clknet_leaf_31_clk _00708_ net8696 VGND VGND VPWR VPWR pid_q.curr_error\[11\]
+ sky130_fd_sc_hd__dfrtp_2
Xwire1157 _04782_ VGND VGND VPWR VPWR net1157 sky130_fd_sc_hd__buf_1
XFILLER_0_16_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1168 _02147_ VGND VGND VPWR VPWR net1168 sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_39_clk clknet_4_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_16
Xwire1179 _01505_ VGND VGND VPWR VPWR net1179 sky130_fd_sc_hd__clkbuf_2
X_12800_ net1343 _04969_ VGND VGND VPWR VPWR _05073_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13780_ _05942_ _06046_ _06047_ VGND VGND VPWR VPWR _06048_ sky130_fd_sc_hd__a21oi_2
X_25766_ clknet_leaf_67_clk _00639_ net8646 VGND VGND VPWR VPWR pid_d.out\[7\] sky130_fd_sc_hd__dfrtp_1
X_22978_ net5243 net720 net6571 VGND VGND VPWR VPWR _02857_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24717_ _04550_ _04551_ net4232 VGND VGND VPWR VPWR _04552_ sky130_fd_sc_hd__a21o_1
X_12731_ _04989_ _05003_ VGND VGND VPWR VPWR _05004_ sky130_fd_sc_hd__xnor2_2
X_21929_ _01933_ _01936_ VGND VGND VPWR VPWR _01937_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_69_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25697_ clknet_leaf_120_clk _00570_ net8395 VGND VGND VPWR VPWR pid_d.mult0.b\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15450_ net1539 net1869 net1872 VGND VGND VPWR VPWR _07524_ sky130_fd_sc_hd__a21o_1
X_24648_ _04446_ _04451_ _04447_ VGND VGND VPWR VPWR _04503_ sky130_fd_sc_hd__o21a_1
X_12662_ _04922_ _04934_ VGND VGND VPWR VPWR _04935_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length5141 net5142 VGND VGND VPWR VPWR net5141 sky130_fd_sc_hd__buf_1
Xfanout8658 net8706 VGND VGND VPWR VPWR net8658 sky130_fd_sc_hd__clkbuf_1
X_14401_ net8151 net3635 VGND VGND VPWR VPWR _06604_ sky130_fd_sc_hd__and2_1
Xfanout8669 net8703 VGND VGND VPWR VPWR net8669 sky130_fd_sc_hd__buf_1
XFILLER_0_26_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15381_ _07327_ _07453_ _07454_ VGND VGND VPWR VPWR _07455_ sky130_fd_sc_hd__mux2_1
X_24579_ _04430_ _04433_ _04434_ VGND VGND VPWR VPWR _04435_ sky130_fd_sc_hd__and3_1
X_12593_ net4384 VGND VGND VPWR VPWR _04875_ sky130_fd_sc_hd__inv_2
Xwire8742 net8731 VGND VGND VPWR VPWR net8742 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_170_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8753 net8755 VGND VGND VPWR VPWR net8753 sky130_fd_sc_hd__buf_1
X_17120_ _09060_ _09062_ net6961 VGND VGND VPWR VPWR _09076_ sky130_fd_sc_hd__o21a_1
Xwire8764 net8765 VGND VGND VPWR VPWR net8764 sky130_fd_sc_hd__buf_1
Xmax_length4451 pid_q.out\[5\] VGND VGND VPWR VPWR net4451 sky130_fd_sc_hd__clkbuf_1
Xwire410 net411 VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14332_ net8253 net3642 VGND VGND VPWR VPWR _06551_ sky130_fd_sc_hd__and2_1
Xmax_length4462 pid_q.out\[3\] VGND VGND VPWR VPWR net4462 sky130_fd_sc_hd__buf_1
Xwire421 _10518_ VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire432 _07829_ VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__clkbuf_1
Xwire8797 net8798 VGND VGND VPWR VPWR net8797 sky130_fd_sc_hd__buf_1
Xwire443 net444 VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__clkbuf_1
Xwire454 _05334_ VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__clkbuf_1
X_17051_ _08971_ _09007_ _09008_ _09009_ _08955_ VGND VGND VPWR VPWR _09010_ sky130_fd_sc_hd__o221a_1
X_14263_ net56 net2931 net2278 net8986 VGND VGND VPWR VPWR _00036_ sky130_fd_sc_hd__a22o_1
Xwire465 net466 VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire476 net477 VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__buf_1
X_16002_ net3546 net2846 net2732 net1846 VGND VGND VPWR VPWR _08070_ sky130_fd_sc_hd__and4_1
Xwire487 _11742_ VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_80_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13214_ net7728 net2368 net2365 VGND VGND VPWR VPWR _05487_ sky130_fd_sc_hd__and3_1
Xwire498 net499 VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__clkbuf_1
X_14194_ _06403_ _06411_ _06415_ VGND VGND VPWR VPWR _06454_ sky130_fd_sc_hd__and3_1
X_13145_ net7877 net1949 _05338_ VGND VGND VPWR VPWR _05418_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13076_ _05290_ _05296_ VGND VGND VPWR VPWR _05349_ sky130_fd_sc_hd__nand2_1
X_17953_ net3239 net3238 _09797_ _09799_ VGND VGND VPWR VPWR _09804_ sky130_fd_sc_hd__a211oi_1
Xwire3060 _03108_ VGND VGND VPWR VPWR net3060 sky130_fd_sc_hd__buf_1
Xwire3071 _02680_ VGND VGND VPWR VPWR net3071 sky130_fd_sc_hd__clkbuf_1
X_16904_ cordic0.slte0.opA\[9\] _08866_ VGND VGND VPWR VPWR _08868_ sky130_fd_sc_hd__nand2_1
Xwire3082 net3086 VGND VGND VPWR VPWR net3082 sky130_fd_sc_hd__buf_1
XFILLER_0_174_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3093 _02546_ VGND VGND VPWR VPWR net3093 sky130_fd_sc_hd__dlymetal6s2s_1
X_17884_ net6873 VGND VGND VPWR VPWR _09735_ sky130_fd_sc_hd__inv_2
Xwire2381 _00006_ VGND VGND VPWR VPWR net2381 sky130_fd_sc_hd__buf_1
X_19623_ net3186 _10918_ VGND VGND VPWR VPWR _11460_ sky130_fd_sc_hd__or2_1
X_16835_ _08808_ VGND VGND VPWR VPWR _00315_ sky130_fd_sc_hd__clkbuf_1
Xwire2392 net2393 VGND VGND VPWR VPWR net2392 sky130_fd_sc_hd__buf_1
XFILLER_0_189_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1680 net1681 VGND VGND VPWR VPWR net1680 sky130_fd_sc_hd__clkbuf_2
Xwire1691 net1692 VGND VGND VPWR VPWR net1691 sky130_fd_sc_hd__clkbuf_1
X_19554_ net6252 net3190 VGND VGND VPWR VPWR _11391_ sky130_fd_sc_hd__nor2_1
X_13978_ net835 _06242_ VGND VGND VPWR VPWR _06243_ sky130_fd_sc_hd__xor2_1
X_16766_ _08772_ VGND VGND VPWR VPWR _00282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18505_ net6775 _10289_ _10351_ VGND VGND VPWR VPWR _10354_ sky130_fd_sc_hd__and3_1
X_12929_ _05102_ _05200_ _05201_ VGND VGND VPWR VPWR _05202_ sky130_fd_sc_hd__a21oi_2
X_15717_ _07786_ _07787_ VGND VGND VPWR VPWR _07788_ sky130_fd_sc_hd__xnor2_1
X_16697_ matmul0.alpha_pass\[11\] net423 net6550 VGND VGND VPWR VPWR _08727_ sky130_fd_sc_hd__mux2_1
X_19485_ net6267 _11318_ _11321_ VGND VGND VPWR VPWR _11322_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_38_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18436_ net7000 net7016 net3297 net6956 VGND VGND VPWR VPWR _10286_ sky130_fd_sc_hd__a22o_1
X_15648_ net2696 _07570_ VGND VGND VPWR VPWR _07720_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15579_ _07647_ _07650_ VGND VGND VPWR VPWR _07651_ sky130_fd_sc_hd__xnor2_1
X_18367_ net6863 net6876 VGND VGND VPWR VPWR _10218_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17318_ net6720 net7787 VGND VGND VPWR VPWR _09232_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18298_ _10075_ _10074_ VGND VGND VPWR VPWR _10149_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17249_ net2164 net192 net1799 net9132 VGND VGND VPWR VPWR _00347_ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20260_ net16 net2 _12065_ VGND VGND VPWR VPWR _12072_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20191_ cordic0.cos\[11\] net2122 net1784 VGND VGND VPWR VPWR _12017_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23950_ _03681_ _03683_ _03682_ VGND VGND VPWR VPWR _03814_ sky130_fd_sc_hd__o21a_1
XFILLER_0_138_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22901_ net338 _02793_ VGND VGND VPWR VPWR _02794_ sky130_fd_sc_hd__nor2_1
X_23881_ _03737_ _03745_ VGND VGND VPWR VPWR _03746_ sky130_fd_sc_hd__xnor2_2
X_25620_ clknet_leaf_116_clk _00493_ net8329 VGND VGND VPWR VPWR cordic0.slte0.opA\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_22832_ net5365 net3065 _02732_ net8897 VGND VGND VPWR VPWR _00634_ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25551_ clknet_leaf_69_clk net6555 net8452 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_22763_ pid_d.ki\[12\] _02686_ net2038 VGND VGND VPWR VPWR _02687_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24502_ net4516 net4537 net3054 net4793 _04358_ VGND VGND VPWR VPWR _04359_ sky130_fd_sc_hd__a32o_1
XFILLER_0_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21714_ _01626_ _01723_ _01722_ VGND VGND VPWR VPWR _01725_ sky130_fd_sc_hd__a21o_1
X_25482_ clknet_leaf_45_clk _00362_ net8789 VGND VGND VPWR VPWR svm0.tA\[4\] sky130_fd_sc_hd__dfrtp_1
X_22694_ _02637_ net5512 net2451 VGND VGND VPWR VPWR _02638_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8005 net8006 VGND VGND VPWR VPWR net8005 sky130_fd_sc_hd__clkbuf_1
X_24433_ net4896 net3745 VGND VGND VPWR VPWR _04291_ sky130_fd_sc_hd__nand2_1
X_21645_ _01570_ _01581_ _01655_ VGND VGND VPWR VPWR _01656_ sky130_fd_sc_hd__o21a_1
XFILLER_0_81_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8038 net8039 VGND VGND VPWR VPWR net8038 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7304 net7305 VGND VGND VPWR VPWR net7304 sky130_fd_sc_hd__clkbuf_1
Xwire8049 net8050 VGND VGND VPWR VPWR net8049 sky130_fd_sc_hd__buf_1
Xwire7315 matmul0.alpha_pass\[5\] VGND VGND VPWR VPWR net7315 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7326 net7327 VGND VGND VPWR VPWR net7326 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24364_ net4993 net4959 net4937 _04147_ VGND VGND VPWR VPWR _04223_ sky130_fd_sc_hd__a31o_1
XFILLER_0_133_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7337 net7338 VGND VGND VPWR VPWR net7337 sky130_fd_sc_hd__buf_1
X_21576_ _01586_ _01587_ VGND VGND VPWR VPWR _01588_ sky130_fd_sc_hd__xnor2_1
Xwire6603 net6597 VGND VGND VPWR VPWR net6603 sky130_fd_sc_hd__buf_1
Xwire7348 net7349 VGND VGND VPWR VPWR net7348 sky130_fd_sc_hd__clkbuf_1
Xwire6614 net6615 VGND VGND VPWR VPWR net6614 sky130_fd_sc_hd__buf_1
Xwire7359 net7360 VGND VGND VPWR VPWR net7359 sky130_fd_sc_hd__clkbuf_1
X_23315_ _02956_ _02959_ _03184_ VGND VGND VPWR VPWR _03185_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_145_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6625 matmul0.matmul_stage_inst.state\[2\] VGND VGND VPWR VPWR net6625 sky130_fd_sc_hd__buf_1
X_20527_ net6804 _08945_ _12312_ _08824_ VGND VGND VPWR VPWR _12313_ sky130_fd_sc_hd__a22o_1
Xwire6636 net6637 VGND VGND VPWR VPWR net6636 sky130_fd_sc_hd__buf_1
X_24295_ net3044 _04154_ VGND VGND VPWR VPWR _04155_ sky130_fd_sc_hd__xnor2_1
Xmax_length3079 _02604_ VGND VGND VPWR VPWR net3079 sky130_fd_sc_hd__buf_1
XFILLER_0_6_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5902 net5895 VGND VGND VPWR VPWR net5902 sky130_fd_sc_hd__clkbuf_1
Xwire6658 net6659 VGND VGND VPWR VPWR net6658 sky130_fd_sc_hd__buf_1
XFILLER_0_43_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5913 net5914 VGND VGND VPWR VPWR net5913 sky130_fd_sc_hd__clkbuf_1
Xwire6669 net6670 VGND VGND VPWR VPWR net6669 sky130_fd_sc_hd__buf_1
XFILLER_0_160_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5924 net5917 VGND VGND VPWR VPWR net5924 sky130_fd_sc_hd__buf_1
X_23246_ _03020_ _03022_ _03115_ VGND VGND VPWR VPWR _03116_ sky130_fd_sc_hd__a21o_1
XFILLER_0_133_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5935 net5931 VGND VGND VPWR VPWR net5935 sky130_fd_sc_hd__clkbuf_1
X_20458_ net8044 cordic0.slte0.opA\[15\] VGND VGND VPWR VPWR _12250_ sky130_fd_sc_hd__nand2_1
Xwire5946 net5947 VGND VGND VPWR VPWR net5946 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length1644 _04529_ VGND VGND VPWR VPWR net1644 sky130_fd_sc_hd__buf_1
Xwire5957 net5953 VGND VGND VPWR VPWR net5957 sky130_fd_sc_hd__clkbuf_1
Xwire5968 pid_d.curr_error\[6\] VGND VGND VPWR VPWR net5968 sky130_fd_sc_hd__clkbuf_2
Xwire5979 pid_d.curr_int\[6\] VGND VGND VPWR VPWR net5979 sky130_fd_sc_hd__buf_1
X_23177_ _03044_ _03045_ _03026_ VGND VGND VPWR VPWR _03047_ sky130_fd_sc_hd__a21oi_1
X_20389_ net865 _12187_ VGND VGND VPWR VPWR _12188_ sky130_fd_sc_hd__xnor2_1
X_22128_ _02128_ _02133_ VGND VGND VPWR VPWR _02134_ sky130_fd_sc_hd__xnor2_1
X_14950_ net3582 net3580 net4143 net4140 VGND VGND VPWR VPWR _07024_ sky130_fd_sc_hd__o22a_1
X_22059_ _02064_ _02065_ VGND VGND VPWR VPWR _02066_ sky130_fd_sc_hd__and2_1
X_13901_ net839 _06110_ _06166_ VGND VGND VPWR VPWR _06167_ sky130_fd_sc_hd__o21a_1
X_14881_ _06958_ VGND VGND VPWR VPWR _00211_ sky130_fd_sc_hd__clkbuf_1
X_13832_ net7744 net1580 VGND VGND VPWR VPWR _06099_ sky130_fd_sc_hd__and2_1
X_16620_ _08660_ VGND VGND VPWR VPWR _00248_ sky130_fd_sc_hd__clkbuf_1
X_25818_ clknet_leaf_37_clk _00691_ net8744 VGND VGND VPWR VPWR pid_q.prev_error\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16551_ _08555_ _08556_ _08609_ VGND VGND VPWR VPWR _08610_ sky130_fd_sc_hd__o21a_1
X_13763_ _06027_ _06029_ _06030_ VGND VGND VPWR VPWR _06031_ sky130_fd_sc_hd__and3_1
X_25749_ clknet_leaf_10_clk _00622_ net8590 VGND VGND VPWR VPWR pid_d.kp\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12714_ net7911 net1981 net2359 VGND VGND VPWR VPWR _04987_ sky130_fd_sc_hd__and3_1
X_15502_ net3407 net3404 VGND VGND VPWR VPWR _07575_ sky130_fd_sc_hd__xnor2_1
X_19270_ _11099_ _11102_ VGND VGND VPWR VPWR _11107_ sky130_fd_sc_hd__nand2_1
X_16482_ _08499_ _08541_ VGND VGND VPWR VPWR _08543_ sky130_fd_sc_hd__nand2_1
XFILLER_0_168_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13694_ net7637 net1149 VGND VGND VPWR VPWR _05963_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15433_ net4172 net4166 net4199 _06977_ VGND VGND VPWR VPWR _07507_ sky130_fd_sc_hd__o22a_1
X_18221_ _10057_ _10071_ VGND VGND VPWR VPWR _10072_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_194_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12645_ net5295 _04892_ net3694 net2990 svm0.vC\[2\] VGND VGND VPWR VPWR _04918_
+ sky130_fd_sc_hd__a32oi_1
XFILLER_0_150_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8488 net8494 VGND VGND VPWR VPWR net8488 sky130_fd_sc_hd__buf_1
Xwire8550 net8537 VGND VGND VPWR VPWR net8550 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18152_ _09998_ net3234 _10002_ VGND VGND VPWR VPWR _10003_ sky130_fd_sc_hd__a21oi_1
X_15364_ net3596 net3590 VGND VGND VPWR VPWR _07438_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8499 net8501 VGND VGND VPWR VPWR net8499 sky130_fd_sc_hd__buf_1
XFILLER_0_109_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12576_ net9148 _04863_ net6597 VGND VGND VPWR VPWR _00012_ sky130_fd_sc_hd__a21o_1
Xwire8572 net8569 VGND VGND VPWR VPWR net8572 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_109_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8583 net8584 VGND VGND VPWR VPWR net8583 sky130_fd_sc_hd__buf_1
XFILLER_0_182_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire240 net241 VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__clkbuf_1
Xwire8594 net8595 VGND VGND VPWR VPWR net8594 sky130_fd_sc_hd__buf_1
X_14315_ matmul0.state\[1\] net6597 cordic_done net6432 VGND VGND VPWR VPWR _06537_
+ sky130_fd_sc_hd__a31o_1
X_17103_ net1476 _09059_ VGND VGND VPWR VPWR _09060_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7860 net7861 VGND VGND VPWR VPWR net7860 sky130_fd_sc_hd__clkbuf_1
X_18083_ net6984 net7066 VGND VGND VPWR VPWR _09934_ sky130_fd_sc_hd__nand2_1
Xwire7871 net7872 VGND VGND VPWR VPWR net7871 sky130_fd_sc_hd__clkbuf_1
X_15295_ net6616 matmul0.matmul_stage_inst.b\[12\] matmul0.matmul_stage_inst.a\[12\]
+ net6589 VGND VGND VPWR VPWR _07369_ sky130_fd_sc_hd__a22o_1
Xwire251 net252 VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__clkbuf_1
Xwire262 _04624_ VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__clkbuf_1
Xwire273 _02390_ VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__clkbuf_1
Xwire7882 net7883 VGND VGND VPWR VPWR net7882 sky130_fd_sc_hd__buf_1
Xwire284 net285 VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__buf_1
Xwire7893 net7894 VGND VGND VPWR VPWR net7893 sky130_fd_sc_hd__dlymetal6s2s_1
X_17034_ _08980_ VGND VGND VPWR VPWR _08994_ sky130_fd_sc_hd__inv_2
Xwire295 net296 VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__clkbuf_1
X_14246_ _06500_ VGND VGND VPWR VPWR _06501_ sky130_fd_sc_hd__buf_1
XFILLER_0_159_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14177_ _06395_ _06421_ VGND VGND VPWR VPWR _06437_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13128_ _05400_ VGND VGND VPWR VPWR _05401_ sky130_fd_sc_hd__clkbuf_2
X_18985_ net6320 net6289 VGND VGND VPWR VPWR _10822_ sky130_fd_sc_hd__nor2b_1
XFILLER_0_187_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13059_ _05330_ _05331_ _05318_ VGND VGND VPWR VPWR _05332_ sky130_fd_sc_hd__mux2_1
X_17936_ net2561 net2559 VGND VGND VPWR VPWR _09787_ sky130_fd_sc_hd__nor2_1
XFILLER_0_178_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17867_ net3258 net3266 net7031 VGND VGND VPWR VPWR _09718_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19606_ net1418 _11403_ _11442_ VGND VGND VPWR VPWR _11443_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16818_ _08799_ VGND VGND VPWR VPWR _00307_ sky130_fd_sc_hd__clkbuf_1
X_17798_ _09648_ VGND VGND VPWR VPWR _09649_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_132_Left_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19537_ _11346_ net3155 _11347_ VGND VGND VPWR VPWR _11374_ sky130_fd_sc_hd__o21a_1
XFILLER_0_177_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16749_ _08763_ VGND VGND VPWR VPWR _00274_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19468_ _11000_ _11006_ _11001_ VGND VGND VPWR VPWR _11305_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_173_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18419_ _10217_ net1210 _10268_ VGND VGND VPWR VPWR _10269_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19399_ _11168_ _11184_ VGND VGND VPWR VPWR _11236_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21430_ net5426 net5894 VGND VGND VPWR VPWR _01443_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21361_ net5865 net5457 VGND VGND VPWR VPWR _01375_ sky130_fd_sc_hd__nand2_1
Xwire5209 matmul0.beta_pass\[12\] VGND VGND VPWR VPWR net5209 sky130_fd_sc_hd__clkbuf_1
X_23100_ net5015 net4718 VGND VGND VPWR VPWR _02970_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20312_ cordic0.slte0.opA\[2\] net2281 _12115_ VGND VGND VPWR VPWR _12117_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_141_Left_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput70 periodTop[14] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_1
X_24080_ _03942_ VGND VGND VPWR VPWR _03943_ sky130_fd_sc_hd__inv_2
Xinput81 pid_d_addr[0] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21292_ net3811 _12515_ _12516_ VGND VGND VPWR VPWR _01307_ sky130_fd_sc_hd__a21o_1
Xwire4508 net4511 VGND VGND VPWR VPWR net4508 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput92 pid_d_addr[5] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_1
Xwire4519 net4521 VGND VGND VPWR VPWR net4519 sky130_fd_sc_hd__buf_1
X_23031_ net4948 net4753 VGND VGND VPWR VPWR _02901_ sky130_fd_sc_hd__nand2_1
X_20243_ net14 _12058_ VGND VGND VPWR VPWR _12059_ sky130_fd_sc_hd__xor2_1
Xwire3807 _01049_ VGND VGND VPWR VPWR net3807 sky130_fd_sc_hd__buf_1
Xwire3818 net3819 VGND VGND VPWR VPWR net3818 sky130_fd_sc_hd__buf_1
X_20174_ net6059 net2580 net6024 VGND VGND VPWR VPWR _12000_ sky130_fd_sc_hd__and3_1
X_24982_ pid_q.kp\[10\] _04722_ net1634 VGND VGND VPWR VPWR _04746_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23933_ _03688_ _03691_ _03796_ VGND VGND VPWR VPWR _03797_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_157_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23864_ _03728_ VGND VGND VPWR VPWR _03729_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_150_Left_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25603_ clknet_leaf_109_clk _00476_ net8345 VGND VGND VPWR VPWR cordic0.slte0.opB\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_22815_ _02717_ net5986 pid_d.out\[0\] VGND VGND VPWR VPWR _02718_ sky130_fd_sc_hd__mux2_1
X_23795_ pid_q.curr_error\[3\] VGND VGND VPWR VPWR _03661_ sky130_fd_sc_hd__inv_2
XFILLER_0_149_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25534_ clknet_leaf_32_clk _00414_ net8692 VGND VGND VPWR VPWR pid_q.prev_int\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_22746_ _02675_ VGND VGND VPWR VPWR _00605_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_183_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25465_ clknet_leaf_53_clk _00345_ net8807 VGND VGND VPWR VPWR svm0.tB\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_176_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22677_ _02626_ VGND VGND VPWR VPWR _00585_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout7039 cordic0.vec\[1\]\[5\] VGND VGND VPWR VPWR net7039 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_165_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24416_ net4791 _04273_ VGND VGND VPWR VPWR _04274_ sky130_fd_sc_hd__xnor2_1
Xwire7101 net7102 VGND VGND VPWR VPWR net7101 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7112 net7110 VGND VGND VPWR VPWR net7112 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout6316 net6322 VGND VGND VPWR VPWR net6316 sky130_fd_sc_hd__clkbuf_1
X_21628_ _01638_ _01639_ VGND VGND VPWR VPWR _01640_ sky130_fd_sc_hd__nand2_1
Xwire7123 net7124 VGND VGND VPWR VPWR net7123 sky130_fd_sc_hd__buf_1
X_25396_ clknet_leaf_76_clk _00279_ net8460 VGND VGND VPWR VPWR matmul0.b\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_164_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6400 net6401 VGND VGND VPWR VPWR net6400 sky130_fd_sc_hd__clkbuf_1
Xwire7145 net7146 VGND VGND VPWR VPWR net7145 sky130_fd_sc_hd__buf_1
XFILLER_0_90_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6411 net6412 VGND VGND VPWR VPWR net6411 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24347_ _04131_ _04133_ _04205_ VGND VGND VPWR VPWR _04206_ sky130_fd_sc_hd__a21bo_1
Xwire7156 net7157 VGND VGND VPWR VPWR net7156 sky130_fd_sc_hd__buf_1
X_21559_ net5806 net5471 VGND VGND VPWR VPWR _01571_ sky130_fd_sc_hd__nand2_1
Xwire7167 matmul0.cos\[12\] VGND VGND VPWR VPWR net7167 sky130_fd_sc_hd__buf_1
Xwire6422 cordic0.sin\[10\] VGND VGND VPWR VPWR net6422 sky130_fd_sc_hd__clkbuf_1
Xwire7178 net7179 VGND VGND VPWR VPWR net7178 sky130_fd_sc_hd__clkbuf_1
Xwire6433 net6434 VGND VGND VPWR VPWR net6433 sky130_fd_sc_hd__clkbuf_1
X_14100_ _06358_ _06362_ VGND VGND VPWR VPWR _06363_ sky130_fd_sc_hd__xnor2_1
Xfanout4903 pid_q.mult0.b\[10\] VGND VGND VPWR VPWR net4903 sky130_fd_sc_hd__buf_1
Xwire7189 matmul0.b\[2\] VGND VGND VPWR VPWR net7189 sky130_fd_sc_hd__clkbuf_1
Xwire5710 net5711 VGND VGND VPWR VPWR net5710 sky130_fd_sc_hd__buf_1
Xwire5721 net5723 VGND VGND VPWR VPWR net5721 sky130_fd_sc_hd__buf_1
X_15080_ _07149_ net3483 net2768 net3486 VGND VGND VPWR VPWR _07154_ sky130_fd_sc_hd__o22a_1
X_24278_ _04081_ _04083_ net3040 VGND VGND VPWR VPWR _04138_ sky130_fd_sc_hd__a21o_1
XFILLER_0_133_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6466 net6463 VGND VGND VPWR VPWR net6466 sky130_fd_sc_hd__buf_1
Xwire5732 net5733 VGND VGND VPWR VPWR net5732 sky130_fd_sc_hd__clkbuf_1
Xwire6477 net6478 VGND VGND VPWR VPWR net6477 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire5743 net5739 VGND VGND VPWR VPWR net5743 sky130_fd_sc_hd__buf_1
X_14031_ _06293_ _06294_ VGND VGND VPWR VPWR _06295_ sky130_fd_sc_hd__xnor2_2
Xwire5754 net5755 VGND VGND VPWR VPWR net5754 sky130_fd_sc_hd__buf_1
Xwire6499 net6500 VGND VGND VPWR VPWR net6499 sky130_fd_sc_hd__buf_1
X_23229_ _02996_ _02997_ VGND VGND VPWR VPWR _03099_ sky130_fd_sc_hd__xnor2_1
Xwire5776 net5774 VGND VGND VPWR VPWR net5776 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire5787 net5788 VGND VGND VPWR VPWR net5787 sky130_fd_sc_hd__clkbuf_1
X_18770_ _10516_ _10604_ _10614_ VGND VGND VPWR VPWR _10615_ sky130_fd_sc_hd__a21oi_1
X_15982_ net1525 net1523 VGND VGND VPWR VPWR _08050_ sky130_fd_sc_hd__and2_1
X_17721_ net9185 net1456 net1789 net5175 VGND VGND VPWR VPWR _00426_ sky130_fd_sc_hd__a22o_1
X_14933_ net1902 net2252 VGND VGND VPWR VPWR _07007_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17652_ _09528_ _09529_ _09530_ _09531_ VGND VGND VPWR VPWR _09532_ sky130_fd_sc_hd__a22o_1
X_14864_ _06949_ VGND VGND VPWR VPWR _00203_ sky130_fd_sc_hd__clkbuf_1
X_16603_ _08651_ VGND VGND VPWR VPWR _00240_ sky130_fd_sc_hd__clkbuf_1
X_13815_ _06080_ _06082_ VGND VGND VPWR VPWR _06083_ sky130_fd_sc_hd__nand2_1
X_17583_ net3278 svm0.tC\[11\] svm0.tC\[10\] _09393_ VGND VGND VPWR VPWR _09465_ sky130_fd_sc_hd__a31o_1
XFILLER_0_159_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14795_ net7441 net3614 VGND VGND VPWR VPWR _06914_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19322_ net3888 net2510 VGND VGND VPWR VPWR _11159_ sky130_fd_sc_hd__xnor2_2
X_13746_ _06012_ _06013_ net404 VGND VGND VPWR VPWR _06014_ sky130_fd_sc_hd__mux2_1
X_16534_ _08593_ VGND VGND VPWR VPWR _00229_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19253_ net1753 _11089_ VGND VGND VPWR VPWR _11090_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13677_ net2300 net2296 net7789 VGND VGND VPWR VPWR _05946_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_128_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16465_ net2623 net2622 net2213 VGND VGND VPWR VPWR _08526_ sky130_fd_sc_hd__or3_1
Xmax_cap4277 _04896_ VGND VGND VPWR VPWR net4277 sky130_fd_sc_hd__buf_1
XFILLER_0_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18204_ _10036_ _10054_ VGND VGND VPWR VPWR _10055_ sky130_fd_sc_hd__xnor2_1
X_12628_ _04900_ VGND VGND VPWR VPWR _04901_ sky130_fd_sc_hd__dlymetal6s2s_1
X_15416_ net2755 net3441 net2696 net2795 VGND VGND VPWR VPWR _07490_ sky130_fd_sc_hd__o211a_1
X_19184_ _11018_ _11019_ _11020_ VGND VGND VPWR VPWR _11021_ sky130_fd_sc_hd__and3b_1
X_16396_ net2204 _08388_ _08457_ net2791 VGND VGND VPWR VPWR _08458_ sky130_fd_sc_hd__o22a_1
XFILLER_0_171_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18135_ _09971_ _09899_ VGND VGND VPWR VPWR _09986_ sky130_fd_sc_hd__nor2_1
X_15347_ net2835 net2702 VGND VGND VPWR VPWR _07421_ sky130_fd_sc_hd__nor2_1
Xfanout6850 cordic0.vec\[1\]\[13\] VGND VGND VPWR VPWR net6850 sky130_fd_sc_hd__clkbuf_2
Xwire8391 net8392 VGND VGND VPWR VPWR net8391 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout6861 net6866 VGND VGND VPWR VPWR net6861 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout6872 net6886 VGND VGND VPWR VPWR net6872 sky130_fd_sc_hd__buf_2
XFILLER_0_79_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7690 net7684 VGND VGND VPWR VPWR net7690 sky130_fd_sc_hd__buf_1
Xfanout6883 net6888 VGND VGND VPWR VPWR net6883 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18066_ _09916_ VGND VGND VPWR VPWR _09917_ sky130_fd_sc_hd__inv_2
Xhold106 cordic0.sin\[0\] VGND VGND VPWR VPWR net9059 sky130_fd_sc_hd__dlygate4sd3_1
X_15278_ net6546 net6594 matmul0.matmul_stage_inst.e\[12\] VGND VGND VPWR VPWR _07352_
+ sky130_fd_sc_hd__o21a_1
Xhold117 svm0.vC\[1\] VGND VGND VPWR VPWR net9070 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold128 matmul0.matmul_stage_inst.b\[1\] VGND VGND VPWR VPWR net9081 sky130_fd_sc_hd__dlygate4sd3_1
X_14229_ net1304 _06484_ _06486_ net1119 VGND VGND VPWR VPWR _06487_ sky130_fd_sc_hd__a22o_1
X_17017_ net7086 _08959_ _08961_ _08960_ VGND VGND VPWR VPWR _08978_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold139 matmul0.matmul_stage_inst.b\[12\] VGND VGND VPWR VPWR net9092 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_107_Right_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18968_ _10800_ net3906 _10802_ net3905 _10804_ VGND VGND VPWR VPWR _10805_ sky130_fd_sc_hd__a221o_1
X_17919_ _09629_ _09767_ _09768_ VGND VGND VPWR VPWR _09770_ sky130_fd_sc_hd__nand3_1
X_18899_ _10738_ _10739_ VGND VGND VPWR VPWR _10740_ sky130_fd_sc_hd__xor2_1
X_20930_ net5575 net5869 VGND VGND VPWR VPWR _00946_ sky130_fd_sc_hd__nand2_1
XFILLER_0_179_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20861_ net1052 _00876_ VGND VGND VPWR VPWR _00877_ sky130_fd_sc_hd__xnor2_2
X_22600_ net2042 _02574_ _02575_ net2459 pid_d.curr_error\[8\] VGND VGND VPWR VPWR
+ _00559_ sky130_fd_sc_hd__a32o_1
XFILLER_0_113_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23580_ _03446_ _03447_ VGND VGND VPWR VPWR _03448_ sky130_fd_sc_hd__and2b_1
X_20792_ _12561_ _12562_ VGND VGND VPWR VPWR _12563_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22531_ net5970 net2380 net2046 VGND VGND VPWR VPWR _02528_ sky130_fd_sc_hd__and3_1
XFILLER_0_187_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25250_ clknet_leaf_87_clk _00133_ net8442 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.a\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22462_ _02461_ _02462_ VGND VGND VPWR VPWR _02463_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24201_ net4520 net4928 VGND VGND VPWR VPWR _04062_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21413_ net4320 net555 VGND VGND VPWR VPWR _01427_ sky130_fd_sc_hd__nand2_1
XFILLER_0_162_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25181_ clknet_leaf_70_clk _00070_ net8452 VGND VGND VPWR VPWR matmul0.a_in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_22393_ net4382 _02336_ net272 net4316 _02395_ VGND VGND VPWR VPWR _02396_ sky130_fd_sc_hd__a221o_1
XFILLER_0_161_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5006 net5007 VGND VGND VPWR VPWR net5006 sky130_fd_sc_hd__clkbuf_1
X_24132_ _03983_ _03993_ VGND VGND VPWR VPWR _03994_ sky130_fd_sc_hd__xnor2_2
Xwire5017 net5018 VGND VGND VPWR VPWR net5017 sky130_fd_sc_hd__buf_1
X_21344_ _01347_ _01357_ VGND VGND VPWR VPWR _01358_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5028 net5029 VGND VGND VPWR VPWR net5028 sky130_fd_sc_hd__buf_1
Xwire5039 net5040 VGND VGND VPWR VPWR net5039 sky130_fd_sc_hd__buf_1
XFILLER_0_163_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4305 net4306 VGND VGND VPWR VPWR net4305 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4316 net4317 VGND VGND VPWR VPWR net4316 sky130_fd_sc_hd__buf_1
X_24063_ net4816 net3042 _03924_ VGND VGND VPWR VPWR _03926_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4327 net4324 VGND VGND VPWR VPWR net4327 sky130_fd_sc_hd__buf_1
X_21275_ net5637 net5674 VGND VGND VPWR VPWR _01290_ sky130_fd_sc_hd__nand2_1
Xwire4338 net4339 VGND VGND VPWR VPWR net4338 sky130_fd_sc_hd__buf_1
Xwire4349 net4350 VGND VGND VPWR VPWR net4349 sky130_fd_sc_hd__clkbuf_1
Xwire3604 net3605 VGND VGND VPWR VPWR net3604 sky130_fd_sc_hd__clkbuf_2
X_23014_ _02881_ _02882_ _02883_ VGND VGND VPWR VPWR _02884_ sky130_fd_sc_hd__o21a_1
Xwire3615 _06862_ VGND VGND VPWR VPWR net3615 sky130_fd_sc_hd__buf_1
X_20226_ _12045_ cordic0.slte0.opB\[5\] net2936 VGND VGND VPWR VPWR _12046_ sky130_fd_sc_hd__mux2_1
Xwire3626 _06818_ VGND VGND VPWR VPWR net3626 sky130_fd_sc_hd__clkbuf_1
Xwire3637 _06575_ VGND VGND VPWR VPWR net3637 sky130_fd_sc_hd__buf_1
Xwire2903 net2904 VGND VGND VPWR VPWR net2903 sky130_fd_sc_hd__buf_1
Xwire3648 _06524_ VGND VGND VPWR VPWR net3648 sky130_fd_sc_hd__buf_1
Xwire3659 net3660 VGND VGND VPWR VPWR net3659 sky130_fd_sc_hd__clkbuf_1
Xwire2925 net2926 VGND VGND VPWR VPWR net2925 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2936 net2937 VGND VGND VPWR VPWR net2936 sky130_fd_sc_hd__clkbuf_2
X_20157_ _11910_ _11930_ VGND VGND VPWR VPWR _11984_ sky130_fd_sc_hd__and2_1
Xwire2947 net2949 VGND VGND VPWR VPWR net2947 sky130_fd_sc_hd__buf_1
Xwire2958 net2960 VGND VGND VPWR VPWR net2958 sky130_fd_sc_hd__buf_1
Xwire2969 net2970 VGND VGND VPWR VPWR net2969 sky130_fd_sc_hd__clkbuf_1
X_24965_ _04737_ VGND VGND VPWR VPWR _00762_ sky130_fd_sc_hd__clkbuf_1
X_20088_ _11914_ _11915_ _11916_ VGND VGND VPWR VPWR _11917_ sky130_fd_sc_hd__a21o_1
X_23916_ _03731_ _03732_ net1162 VGND VGND VPWR VPWR _03780_ sky130_fd_sc_hd__a21bo_1
X_24896_ _04688_ net4525 net2399 VGND VGND VPWR VPWR _04689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length8355 net8356 VGND VGND VPWR VPWR net8355 sky130_fd_sc_hd__buf_1
XFILLER_0_196_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23847_ net4704 net4811 VGND VGND VPWR VPWR _03712_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13600_ _05784_ net533 VGND VGND VPWR VPWR _05870_ sky130_fd_sc_hd__nand2_1
XFILLER_0_196_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14580_ _04860_ _06755_ VGND VGND VPWR VPWR _06756_ sky130_fd_sc_hd__nand2_1
X_23778_ net4708 net4729 _03372_ VGND VGND VPWR VPWR _03644_ sky130_fd_sc_hd__and3_1
X_13531_ net912 net997 net998 VGND VGND VPWR VPWR _05802_ sky130_fd_sc_hd__a21o_1
X_25517_ clknet_leaf_41_clk _00397_ net8784 VGND VGND VPWR VPWR svm0.counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_22729_ net3718 net104 VGND VGND VPWR VPWR _02664_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16250_ net2210 _08313_ VGND VGND VPWR VPWR _08314_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13462_ _05731_ _05734_ VGND VGND VPWR VPWR _05735_ sky130_fd_sc_hd__xnor2_1
X_25448_ clknet_leaf_113_clk _00331_ net8340 VGND VGND VPWR VPWR cordic0.vec\[1\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_165_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6113 net6118 VGND VGND VPWR VPWR net6113 sky130_fd_sc_hd__buf_1
XFILLER_0_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15201_ _07274_ VGND VGND VPWR VPWR _07275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout6146 cordic0.vec\[0\]\[10\] VGND VGND VPWR VPWR net6146 sky130_fd_sc_hd__buf_1
X_16181_ _08186_ _08206_ VGND VGND VPWR VPWR _08246_ sky130_fd_sc_hd__and2_1
X_25379_ clknet_leaf_64_clk _00262_ net8663 VGND VGND VPWR VPWR matmul0.alpha_pass\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13393_ net684 _05664_ _05665_ VGND VGND VPWR VPWR _05666_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout5423 net5448 VGND VGND VPWR VPWR net5423 sky130_fd_sc_hd__clkbuf_1
Xwire6230 net6232 VGND VGND VPWR VPWR net6230 sky130_fd_sc_hd__buf_1
X_15132_ net2759 net2749 VGND VGND VPWR VPWR _07206_ sky130_fd_sc_hd__nor2_1
Xwire6241 net6242 VGND VGND VPWR VPWR net6241 sky130_fd_sc_hd__buf_1
Xwire6252 net6250 VGND VGND VPWR VPWR net6252 sky130_fd_sc_hd__clkbuf_2
Xwire6274 net6269 VGND VGND VPWR VPWR net6274 sky130_fd_sc_hd__buf_1
Xfanout5478 net5489 VGND VGND VPWR VPWR net5478 sky130_fd_sc_hd__clkbuf_1
Xwire6285 cordic0.vec\[0\]\[4\] VGND VGND VPWR VPWR net6285 sky130_fd_sc_hd__buf_1
Xfanout4744 pid_q.mult0.a\[2\] VGND VGND VPWR VPWR net4744 sky130_fd_sc_hd__buf_1
XFILLER_0_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19940_ _11744_ _11771_ VGND VGND VPWR VPWR _11772_ sky130_fd_sc_hd__xnor2_1
X_15063_ matmul0.matmul_stage_inst.e\[11\] _07135_ _07136_ net7382 VGND VGND VPWR
+ VPWR _07137_ sky130_fd_sc_hd__a22o_1
Xwire5551 net5548 VGND VGND VPWR VPWR net5551 sky130_fd_sc_hd__buf_1
XFILLER_0_121_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6296 net6295 VGND VGND VPWR VPWR net6296 sky130_fd_sc_hd__buf_1
Xwire5562 net5556 VGND VGND VPWR VPWR net5562 sky130_fd_sc_hd__buf_1
Xwire5573 net5574 VGND VGND VPWR VPWR net5573 sky130_fd_sc_hd__clkbuf_1
X_14014_ _06260_ VGND VGND VPWR VPWR _06278_ sky130_fd_sc_hd__inv_2
Xwire5584 net5585 VGND VGND VPWR VPWR net5584 sky130_fd_sc_hd__buf_1
Xwire4850 net4851 VGND VGND VPWR VPWR net4850 sky130_fd_sc_hd__buf_1
Xwire4861 pid_q.mult0.b\[12\] VGND VGND VPWR VPWR net4861 sky130_fd_sc_hd__buf_1
XFILLER_0_121_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19871_ _11698_ _11703_ VGND VGND VPWR VPWR _11704_ sky130_fd_sc_hd__xnor2_1
Xwire4872 net4871 VGND VGND VPWR VPWR net4872 sky130_fd_sc_hd__buf_1
Xwire4883 net4884 VGND VGND VPWR VPWR net4883 sky130_fd_sc_hd__buf_1
X_18822_ _10661_ _10663_ VGND VGND VPWR VPWR _10665_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18753_ _10597_ net2127 VGND VGND VPWR VPWR _10598_ sky130_fd_sc_hd__nor2_1
X_15965_ _07970_ net1522 _07967_ VGND VGND VPWR VPWR _08033_ sky130_fd_sc_hd__o21ba_1
X_17704_ net1455 VGND VGND VPWR VPWR _09580_ sky130_fd_sc_hd__clkbuf_1
X_14916_ _06988_ _06989_ _06981_ _06986_ VGND VGND VPWR VPWR _06990_ sky130_fd_sc_hd__a22o_1
X_18684_ net6896 net6877 VGND VGND VPWR VPWR _10530_ sky130_fd_sc_hd__nand2_1
X_15896_ net3515 net3465 VGND VGND VPWR VPWR _07965_ sky130_fd_sc_hd__nor2_1
X_17635_ svm0.tB\[15\] _09472_ net4030 VGND VGND VPWR VPWR _09516_ sky130_fd_sc_hd__a21o_1
X_14847_ matmul0.a\[12\] matmul0.matmul_stage_inst.e\[12\] net3607 VGND VGND VPWR
+ VPWR _06941_ sky130_fd_sc_hd__mux2_1
X_17566_ net6739 svm0.tC\[0\] VGND VGND VPWR VPWR _09448_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14778_ matmul0.sin\[12\] _06902_ VGND VGND VPWR VPWR _06903_ sky130_fd_sc_hd__xnor2_1
X_19305_ net6312 net6352 net6338 VGND VGND VPWR VPWR _11142_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_86_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16517_ net2208 _08575_ VGND VGND VPWR VPWR _08577_ sky130_fd_sc_hd__nor2_1
X_13729_ _05993_ _05994_ _05997_ _05931_ VGND VGND VPWR VPWR _05998_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_2_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17497_ net6705 net2579 VGND VGND VPWR VPWR _09386_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19236_ net6321 _11072_ net3206 VGND VGND VPWR VPWR _11073_ sky130_fd_sc_hd__a21oi_1
X_16448_ _08507_ _08508_ net2245 VGND VGND VPWR VPWR _08509_ sky130_fd_sc_hd__a21o_1
XFILLER_0_116_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19167_ _10947_ _10948_ VGND VGND VPWR VPWR _11004_ sky130_fd_sc_hd__nand2_1
XFILLER_0_171_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16379_ net2841 net2682 net1250 VGND VGND VPWR VPWR _08441_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_182_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18118_ _09967_ _09961_ _09964_ VGND VGND VPWR VPWR _09969_ sky130_fd_sc_hd__nand3_1
XFILLER_0_14_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19098_ _10934_ net1757 VGND VGND VPWR VPWR _10935_ sky130_fd_sc_hd__or2b_1
XFILLER_0_83_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18049_ _09887_ _09895_ VGND VGND VPWR VPWR _09900_ sky130_fd_sc_hd__xor2_2
XFILLER_0_2_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21060_ _01029_ _01065_ _01075_ VGND VGND VPWR VPWR _01076_ sky130_fd_sc_hd__o21ai_1
X_20011_ net567 _11716_ _11739_ _11823_ _11836_ VGND VGND VPWR VPWR _11841_ sky130_fd_sc_hd__a2111o_1
Xwire1509 net1510 VGND VGND VPWR VPWR net1509 sky130_fd_sc_hd__buf_1
X_24750_ net8002 _04572_ VGND VGND VPWR VPWR _04581_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21962_ _01845_ _01856_ net1719 VGND VGND VPWR VPWR _01970_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_69_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23701_ _03475_ _03476_ _03567_ VGND VGND VPWR VPWR _03568_ sky130_fd_sc_hd__a21o_1
X_20913_ _12536_ _00928_ VGND VGND VPWR VPWR _00929_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24681_ net5167 net3021 net1646 VGND VGND VPWR VPWR _04523_ sky130_fd_sc_hd__and3_1
X_21893_ _01894_ _01899_ _01901_ VGND VGND VPWR VPWR _01902_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23632_ _03497_ _03498_ VGND VGND VPWR VPWR _03499_ sky130_fd_sc_hd__xor2_1
X_20844_ _00838_ _00859_ VGND VGND VPWR VPWR _00860_ sky130_fd_sc_hd__xnor2_2
Xmax_length5526 net5527 VGND VGND VPWR VPWR net5526 sky130_fd_sc_hd__clkbuf_1
X_23563_ _03350_ _03352_ _03351_ VGND VGND VPWR VPWR _03431_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20775_ _12542_ _12545_ VGND VGND VPWR VPWR _12546_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_193_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25302_ clknet_leaf_70_clk _00185_ net8459 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.e\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_22514_ _02457_ net517 VGND VGND VPWR VPWR _02515_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23494_ _03354_ _03362_ VGND VGND VPWR VPWR _03363_ sky130_fd_sc_hd__xnor2_2
Xmax_length4847 net4848 VGND VGND VPWR VPWR net4847 sky130_fd_sc_hd__clkbuf_1
Xwire806 _01411_ VGND VGND VPWR VPWR net806 sky130_fd_sc_hd__clkbuf_2
Xwire817 _10019_ VGND VGND VPWR VPWR net817 sky130_fd_sc_hd__clkbuf_1
X_25233_ clknet_leaf_23_clk _00016_ net8587 VGND VGND VPWR VPWR pid_q.state\[0\] sky130_fd_sc_hd__dfstp_1
Xwire828 _07860_ VGND VGND VPWR VPWR net828 sky130_fd_sc_hd__clkbuf_1
Xwire839 _06109_ VGND VGND VPWR VPWR net839 sky130_fd_sc_hd__buf_1
XFILLER_0_161_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22445_ net944 _02446_ VGND VGND VPWR VPWR _02447_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_88_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25164_ clknet_leaf_54_clk _00053_ net8730 VGND VGND VPWR VPWR svm0.periodTop\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22376_ _02377_ _02378_ VGND VGND VPWR VPWR _02379_ sky130_fd_sc_hd__and2b_1
XFILLER_0_5_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24115_ _03885_ _03888_ _03872_ VGND VGND VPWR VPWR _03977_ sky130_fd_sc_hd__o21ba_1
Xwire4102 net4103 VGND VGND VPWR VPWR net4102 sky130_fd_sc_hd__clkbuf_1
X_21327_ _01339_ _01340_ VGND VGND VPWR VPWR _01341_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_4_4__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_4_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_25095_ net4401 net5172 _04837_ _04838_ VGND VGND VPWR VPWR _04839_ sky130_fd_sc_hd__o211ai_2
Xwire4113 _07126_ VGND VGND VPWR VPWR net4113 sky130_fd_sc_hd__clkbuf_1
Xwire4124 net4125 VGND VGND VPWR VPWR net4124 sky130_fd_sc_hd__buf_1
XFILLER_0_13_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4135 net4136 VGND VGND VPWR VPWR net4135 sky130_fd_sc_hd__clkbuf_1
Xwire3401 net3402 VGND VGND VPWR VPWR net3401 sky130_fd_sc_hd__clkbuf_1
X_24046_ _03897_ _03908_ VGND VGND VPWR VPWR _03909_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4146 net4147 VGND VGND VPWR VPWR net4146 sky130_fd_sc_hd__buf_1
Xwire4157 net4158 VGND VGND VPWR VPWR net4157 sky130_fd_sc_hd__buf_1
Xwire3412 _07528_ VGND VGND VPWR VPWR net3412 sky130_fd_sc_hd__buf_1
X_21258_ _00825_ _00830_ _00823_ VGND VGND VPWR VPWR _01273_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3423 _07507_ VGND VGND VPWR VPWR net3423 sky130_fd_sc_hd__buf_1
Xwire4168 _07003_ VGND VGND VPWR VPWR net4168 sky130_fd_sc_hd__clkbuf_1
Xwire4179 net4180 VGND VGND VPWR VPWR net4179 sky130_fd_sc_hd__buf_1
Xwire3434 net3437 VGND VGND VPWR VPWR net3434 sky130_fd_sc_hd__buf_1
XFILLER_0_25_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3445 net3446 VGND VGND VPWR VPWR net3445 sky130_fd_sc_hd__clkbuf_1
Xwire2700 net2701 VGND VGND VPWR VPWR net2700 sky130_fd_sc_hd__clkbuf_2
Xwire3456 net3457 VGND VGND VPWR VPWR net3456 sky130_fd_sc_hd__buf_1
Xwire2711 net2713 VGND VGND VPWR VPWR net2711 sky130_fd_sc_hd__clkbuf_1
X_20209_ cordic0.cos\[13\] net2123 net1784 VGND VGND VPWR VPWR _12033_ sky130_fd_sc_hd__and3_1
Xwire2722 net2723 VGND VGND VPWR VPWR net2722 sky130_fd_sc_hd__buf_1
X_21189_ _01157_ _01161_ _01148_ VGND VGND VPWR VPWR _01205_ sky130_fd_sc_hd__or3b_1
Xwire2733 net2734 VGND VGND VPWR VPWR net2733 sky130_fd_sc_hd__buf_1
Xwire3478 net3479 VGND VGND VPWR VPWR net3478 sky130_fd_sc_hd__buf_1
Xwire3489 net3490 VGND VGND VPWR VPWR net3489 sky130_fd_sc_hd__buf_1
Xwire2744 net2745 VGND VGND VPWR VPWR net2744 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2755 net2756 VGND VGND VPWR VPWR net2755 sky130_fd_sc_hd__buf_1
Xwire2766 net2767 VGND VGND VPWR VPWR net2766 sky130_fd_sc_hd__buf_1
Xwire2788 _07138_ VGND VGND VPWR VPWR net2788 sky130_fd_sc_hd__buf_1
XFILLER_0_95_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2799 net2800 VGND VGND VPWR VPWR net2799 sky130_fd_sc_hd__buf_1
X_12962_ net1002 _05234_ VGND VGND VPWR VPWR _05235_ sky130_fd_sc_hd__nand2_1
X_15750_ _07712_ _07732_ _07820_ VGND VGND VPWR VPWR _07821_ sky130_fd_sc_hd__a21o_1
X_24948_ net8870 net133 VGND VGND VPWR VPWR _04726_ sky130_fd_sc_hd__and2b_1
XFILLER_0_99_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14701_ net7151 _06845_ VGND VGND VPWR VPWR _06846_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_169_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12893_ _05159_ _05164_ _05165_ VGND VGND VPWR VPWR _05166_ sky130_fd_sc_hd__and3_1
X_15681_ net3498 net3413 VGND VGND VPWR VPWR _07752_ sky130_fd_sc_hd__nor2_2
X_24879_ _04677_ VGND VGND VPWR VPWR _00736_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_185_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17420_ net611 _09321_ _09319_ VGND VGND VPWR VPWR _09322_ sky130_fd_sc_hd__a21oi_1
Xmax_length7451 net7452 VGND VGND VPWR VPWR net7451 sky130_fd_sc_hd__clkbuf_1
X_14632_ _06798_ VGND VGND VPWR VPWR _00122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17351_ net4031 net7607 _09214_ net7630 _09264_ VGND VGND VPWR VPWR _09265_ sky130_fd_sc_hd__a221o_1
X_14563_ net7257 _06738_ _06739_ VGND VGND VPWR VPWR _06740_ sky130_fd_sc_hd__a21o_1
XFILLER_0_184_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16302_ _08245_ _08365_ _08360_ VGND VGND VPWR VPWR _08366_ sky130_fd_sc_hd__o21bai_1
X_13514_ net7786 net1586 VGND VGND VPWR VPWR _05785_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17282_ net4035 net6738 svm0.counter\[3\] net6736 VGND VGND VPWR VPWR _09197_ sky130_fd_sc_hd__or4_1
X_14494_ net9047 net831 net1292 _06677_ VGND VGND VPWR VPWR _00105_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19021_ _10855_ _10857_ VGND VGND VPWR VPWR _10858_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13445_ _05715_ _05716_ _05601_ _05717_ _05595_ VGND VGND VPWR VPWR _05718_ sky130_fd_sc_hd__o32a_1
X_16233_ net1088 net1511 _08214_ VGND VGND VPWR VPWR _08298_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_67_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13376_ _05645_ _05646_ VGND VGND VPWR VPWR _05649_ sky130_fd_sc_hd__nor2_1
X_16164_ _08226_ _08229_ VGND VGND VPWR VPWR _08230_ sky130_fd_sc_hd__xor2_1
XFILLER_0_2_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6060 net6062 VGND VGND VPWR VPWR net6060 sky130_fd_sc_hd__buf_1
Xwire6071 net6072 VGND VGND VPWR VPWR net6071 sky130_fd_sc_hd__buf_1
X_15115_ net4160 net4156 VGND VGND VPWR VPWR _07189_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6082 net6080 VGND VGND VPWR VPWR net6082 sky130_fd_sc_hd__clkbuf_1
X_16095_ matmul0.matmul_stage_inst.mult1\[7\] net354 net2679 VGND VGND VPWR VPWR _08162_
+ sky130_fd_sc_hd__mux2_1
Xwire6093 net6094 VGND VGND VPWR VPWR net6093 sky130_fd_sc_hd__buf_1
XFILLER_0_181_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_192_Right_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5370 net5371 VGND VGND VPWR VPWR net5370 sky130_fd_sc_hd__buf_1
XFILLER_0_103_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19923_ net6027 net3125 VGND VGND VPWR VPWR _11755_ sky130_fd_sc_hd__xnor2_2
X_15046_ _07116_ _07117_ _07119_ VGND VGND VPWR VPWR _07120_ sky130_fd_sc_hd__o21a_1
XFILLER_0_167_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5392 net5397 VGND VGND VPWR VPWR net5392 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19854_ net6110 net6127 net6212 VGND VGND VPWR VPWR _11687_ sky130_fd_sc_hd__nand3b_1
Xwire4691 pid_q.mult0.a\[5\] VGND VGND VPWR VPWR net4691 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18805_ _10629_ _10648_ VGND VGND VPWR VPWR _10649_ sky130_fd_sc_hd__xnor2_2
Xwire3990 net3991 VGND VGND VPWR VPWR net3990 sky130_fd_sc_hd__buf_1
X_19785_ _11613_ _11614_ _11615_ _11618_ _11488_ VGND VGND VPWR VPWR _11619_ sky130_fd_sc_hd__a32o_1
X_16997_ net2173 _08958_ VGND VGND VPWR VPWR _08959_ sky130_fd_sc_hd__xnor2_1
X_18736_ net3985 _10580_ net6855 VGND VGND VPWR VPWR _10581_ sky130_fd_sc_hd__mux2_1
X_15948_ net1527 net1262 _08015_ VGND VGND VPWR VPWR _08016_ sky130_fd_sc_hd__o21ai_2
X_18667_ _10503_ _10504_ _10502_ VGND VGND VPWR VPWR _10513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15879_ _07946_ _07947_ VGND VGND VPWR VPWR _07948_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17618_ _09495_ _09496_ _09497_ _09498_ VGND VGND VPWR VPWR _09499_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18598_ net3930 net3281 VGND VGND VPWR VPWR _10446_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17549_ svm0.tC\[6\] net6722 VGND VGND VPWR VPWR _09431_ sky130_fd_sc_hd__and2b_1
XFILLER_0_73_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20560_ _12337_ _12344_ VGND VGND VPWR VPWR _12345_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19219_ net6271 _10822_ VGND VGND VPWR VPWR _11056_ sky130_fd_sc_hd__xnor2_2
X_20491_ net6758 net2492 net3345 VGND VGND VPWR VPWR _12279_ sky130_fd_sc_hd__mux2_1
X_22230_ net1389 _02145_ _02234_ VGND VGND VPWR VPWR _02235_ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22161_ _02119_ _02166_ VGND VGND VPWR VPWR _02167_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21112_ net5644 net5833 VGND VGND VPWR VPWR _01128_ sky130_fd_sc_hd__nand2_1
X_22092_ _02022_ _02098_ VGND VGND VPWR VPWR _02099_ sky130_fd_sc_hd__xnor2_1
Xwire2007 net2008 VGND VGND VPWR VPWR net2007 sky130_fd_sc_hd__buf_1
X_25920_ clknet_leaf_96_clk _00793_ net8400 VGND VGND VPWR VPWR pid_d.prev_int\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_21043_ net2075 net2074 net1731 net2480 _01058_ VGND VGND VPWR VPWR _01059_ sky130_fd_sc_hd__a311o_1
Xwire2018 _04280_ VGND VGND VPWR VPWR net2018 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2029 _02870_ VGND VGND VPWR VPWR net2029 sky130_fd_sc_hd__buf_1
Xwire1306 net1307 VGND VGND VPWR VPWR net1306 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1317 net1318 VGND VGND VPWR VPWR net1317 sky130_fd_sc_hd__buf_1
X_25851_ clknet_leaf_20_clk _00724_ net8616 VGND VGND VPWR VPWR pid_q.mult0.b\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1328 net1329 VGND VGND VPWR VPWR net1328 sky130_fd_sc_hd__buf_1
Xwire1339 net1340 VGND VGND VPWR VPWR net1339 sky130_fd_sc_hd__buf_1
X_24802_ net7961 _04620_ _06533_ _04618_ VGND VGND VPWR VPWR _04626_ sky130_fd_sc_hd__a211o_1
Xclkbuf_4_12__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_4_12__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_22994_ net2885 _06513_ VGND VGND VPWR VPWR _02865_ sky130_fd_sc_hd__nor2_1
X_25782_ clknet_leaf_82_clk _00655_ net8500 VGND VGND VPWR VPWR matmul0.beta_pass\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24733_ net8012 _04557_ VGND VGND VPWR VPWR _04566_ sky130_fd_sc_hd__or2_1
X_21945_ _01941_ _01952_ VGND VGND VPWR VPWR _01953_ sky130_fd_sc_hd__xor2_1
XFILLER_0_9_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6002 net5999 VGND VGND VPWR VPWR net6002 sky130_fd_sc_hd__buf_1
XFILLER_0_173_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24664_ net9175 net1377 _04514_ VGND VGND VPWR VPWR _00684_ sky130_fd_sc_hd__a21o_1
X_21876_ _01878_ _01884_ VGND VGND VPWR VPWR _01885_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_194_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout8807 net8812 VGND VGND VPWR VPWR net8807 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_179_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23615_ pid_q.prev_int\[2\] _03391_ net5180 VGND VGND VPWR VPWR _03482_ sky130_fd_sc_hd__a21o_1
Xmax_length6057 net6051 VGND VGND VPWR VPWR net6057 sky130_fd_sc_hd__clkbuf_2
X_20827_ _00841_ _00842_ VGND VGND VPWR VPWR _00843_ sky130_fd_sc_hd__xnor2_1
X_24595_ net328 _04449_ _04450_ VGND VGND VPWR VPWR _04451_ sky130_fd_sc_hd__o21ai_2
Xwire8902 net8903 VGND VGND VPWR VPWR net8902 sky130_fd_sc_hd__buf_1
XFILLER_0_194_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8913 net8914 VGND VGND VPWR VPWR net8913 sky130_fd_sc_hd__clkbuf_1
Xwire8924 net8925 VGND VGND VPWR VPWR net8924 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8935 net103 VGND VGND VPWR VPWR net8935 sky130_fd_sc_hd__clkbuf_1
Xmax_length4622 pid_q.mult0.a\[8\] VGND VGND VPWR VPWR net4622 sky130_fd_sc_hd__clkbuf_1
X_23546_ _03412_ _03413_ VGND VGND VPWR VPWR _03414_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_147_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20758_ _12527_ _12528_ VGND VGND VPWR VPWR _12529_ sky130_fd_sc_hd__xnor2_1
Xwire8946 net8947 VGND VGND VPWR VPWR net8946 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire603 _12186_ VGND VGND VPWR VPWR net603 sky130_fd_sc_hd__clkbuf_1
Xwire614 _09276_ VGND VGND VPWR VPWR net614 sky130_fd_sc_hd__buf_1
Xwire625 net626 VGND VGND VPWR VPWR net625 sky130_fd_sc_hd__buf_1
Xmax_length3921 _10597_ VGND VGND VPWR VPWR net3921 sky130_fd_sc_hd__clkbuf_1
X_23477_ net2424 _03345_ VGND VGND VPWR VPWR _03346_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_162_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire636 net637 VGND VGND VPWR VPWR net636 sky130_fd_sc_hd__clkbuf_1
X_20689_ _12451_ _12452_ VGND VGND VPWR VPWR _12464_ sky130_fd_sc_hd__or2_1
Xwire647 net648 VGND VGND VPWR VPWR net647 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13230_ _05456_ _05461_ _05502_ VGND VGND VPWR VPWR _05503_ sky130_fd_sc_hd__o21a_1
X_25216_ clknet_leaf_59_clk _00105_ net8732 VGND VGND VPWR VPWR svm0.vC\[4\] sky130_fd_sc_hd__dfrtp_1
Xwire658 _10692_ VGND VGND VPWR VPWR net658 sky130_fd_sc_hd__buf_1
Xwire669 _09270_ VGND VGND VPWR VPWR net669 sky130_fd_sc_hd__buf_1
X_22428_ _02351_ _02356_ _02347_ VGND VGND VPWR VPWR _02430_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25147_ clknet_leaf_41_clk _00036_ net8767 VGND VGND VPWR VPWR pid_q.target\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13161_ _05383_ _05385_ _05384_ VGND VGND VPWR VPWR _05434_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22359_ _02284_ _02286_ _02361_ VGND VGND VPWR VPWR _02362_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13092_ _05362_ _05363_ _05361_ VGND VGND VPWR VPWR _05365_ sky130_fd_sc_hd__a21o_1
X_25078_ _04822_ _04817_ _04823_ VGND VGND VPWR VPWR _04824_ sky130_fd_sc_hd__a21oi_2
Xwire3220 _10789_ VGND VGND VPWR VPWR net3220 sky130_fd_sc_hd__clkbuf_1
X_24029_ _03817_ _03822_ _03891_ VGND VGND VPWR VPWR _03892_ sky130_fd_sc_hd__o21ai_2
X_16920_ cordic0.slte0.opA\[4\] VGND VGND VPWR VPWR _08884_ sky130_fd_sc_hd__inv_2
Xwire3231 net3232 VGND VGND VPWR VPWR net3231 sky130_fd_sc_hd__clkbuf_2
Xwire3242 net3243 VGND VGND VPWR VPWR net3242 sky130_fd_sc_hd__buf_1
XFILLER_0_137_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3264 _09615_ VGND VGND VPWR VPWR net3264 sky130_fd_sc_hd__buf_1
Xwire3275 _09332_ VGND VGND VPWR VPWR net3275 sky130_fd_sc_hd__buf_1
Xwire2530 _10799_ VGND VGND VPWR VPWR net2530 sky130_fd_sc_hd__clkbuf_2
Xwire2541 net2542 VGND VGND VPWR VPWR net2541 sky130_fd_sc_hd__clkbuf_2
X_16851_ _08816_ VGND VGND VPWR VPWR _00323_ sky130_fd_sc_hd__clkbuf_1
Xwire2552 _09794_ VGND VGND VPWR VPWR net2552 sky130_fd_sc_hd__buf_1
Xwire3297 net3299 VGND VGND VPWR VPWR net3297 sky130_fd_sc_hd__buf_1
Xwire2563 _09631_ VGND VGND VPWR VPWR net2563 sky130_fd_sc_hd__clkbuf_2
Xwire2574 net2575 VGND VGND VPWR VPWR net2574 sky130_fd_sc_hd__buf_1
XFILLER_0_102_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2585 _09164_ VGND VGND VPWR VPWR net2585 sky130_fd_sc_hd__clkbuf_1
X_15802_ net2732 net2788 VGND VGND VPWR VPWR _07872_ sky130_fd_sc_hd__nand2_1
Xwire1840 _08396_ VGND VGND VPWR VPWR net1840 sky130_fd_sc_hd__buf_1
X_19570_ _11332_ _11338_ _11406_ VGND VGND VPWR VPWR _11407_ sky130_fd_sc_hd__o21ai_1
Xwire1851 _07676_ VGND VGND VPWR VPWR net1851 sky130_fd_sc_hd__buf_1
Xwire2596 net2598 VGND VGND VPWR VPWR net2596 sky130_fd_sc_hd__buf_1
X_16782_ _08780_ VGND VGND VPWR VPWR _00290_ sky130_fd_sc_hd__clkbuf_1
X_13994_ _06172_ net677 _06208_ VGND VGND VPWR VPWR _06259_ sky130_fd_sc_hd__a21o_1
Xwire1862 net1863 VGND VGND VPWR VPWR net1862 sky130_fd_sc_hd__clkbuf_1
Xwire1873 net1874 VGND VGND VPWR VPWR net1873 sky130_fd_sc_hd__clkbuf_1
Xwire1884 net1885 VGND VGND VPWR VPWR net1884 sky130_fd_sc_hd__buf_1
X_18521_ net6818 net6793 _10369_ net6860 VGND VGND VPWR VPWR _10370_ sky130_fd_sc_hd__a211o_1
XFILLER_0_1_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15733_ net1269 net1268 _07803_ VGND VGND VPWR VPWR _07804_ sky130_fd_sc_hd__o21a_1
Xwire1895 _07103_ VGND VGND VPWR VPWR net1895 sky130_fd_sc_hd__buf_1
X_12945_ net7916 net7883 _05216_ _05217_ VGND VGND VPWR VPWR _05218_ sky130_fd_sc_hd__and4_1
XFILLER_0_133_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18452_ net3961 net7045 VGND VGND VPWR VPWR _10302_ sky130_fd_sc_hd__nor2_1
X_15664_ _07645_ _07735_ VGND VGND VPWR VPWR _07736_ sky130_fd_sc_hd__xnor2_1
X_12876_ _05079_ _05083_ _05032_ VGND VGND VPWR VPWR _05149_ sky130_fd_sc_hd__and3b_1
X_17403_ svm0.delta\[8\] net1461 VGND VGND VPWR VPWR _09308_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14615_ net6432 _06786_ cordic_done VGND VGND VPWR VPWR _06787_ sky130_fd_sc_hd__a21o_1
X_18383_ net3241 _10233_ _09909_ VGND VGND VPWR VPWR _10234_ sky130_fd_sc_hd__a21o_1
X_15595_ net1108 _07666_ VGND VGND VPWR VPWR _07667_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_83_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17334_ net4017 _09246_ _09247_ VGND VGND VPWR VPWR _09248_ sky130_fd_sc_hd__o21ba_1
X_14546_ _06653_ _06721_ _06724_ _06651_ net8964 VGND VGND VPWR VPWR _00110_ sky130_fd_sc_hd__a32o_1
XFILLER_0_55_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17265_ net2160 net287 net1798 net9108 VGND VGND VPWR VPWR _00359_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14477_ net7340 net5296 VGND VGND VPWR VPWR _06663_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_183_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19004_ _10836_ net3211 _10838_ _10840_ VGND VGND VPWR VPWR _10841_ sky130_fd_sc_hd__a22o_1
X_16216_ _08279_ _08280_ VGND VGND VPWR VPWR _08281_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_181_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13428_ net7770 net2307 net1952 VGND VGND VPWR VPWR _05701_ sky130_fd_sc_hd__and3_1
X_17196_ _09142_ _09145_ VGND VGND VPWR VPWR _09146_ sky130_fd_sc_hd__xor2_2
Xfanout5061 net5073 VGND VGND VPWR VPWR net5061 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13359_ _05629_ net842 VGND VGND VPWR VPWR _05632_ sky130_fd_sc_hd__xor2_1
X_16147_ net1093 net1092 _08127_ VGND VGND VPWR VPWR _08213_ sky130_fd_sc_hd__o21a_1
XFILLER_0_178_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5072 pid_q.mult0.b\[3\] VGND VGND VPWR VPWR net5072 sky130_fd_sc_hd__buf_1
Xfanout5083 net5104 VGND VGND VPWR VPWR net5083 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16078_ net2224 _08026_ _08028_ _08143_ _08144_ VGND VGND VPWR VPWR _08145_ sky130_fd_sc_hd__a311o_1
XFILLER_0_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19906_ _11661_ net708 _11737_ VGND VGND VPWR VPWR _11738_ sky130_fd_sc_hd__a21oi_1
X_15029_ _07097_ _07098_ _07102_ VGND VGND VPWR VPWR _07103_ sky130_fd_sc_hd__a21o_1
X_19837_ _11661_ _11670_ VGND VGND VPWR VPWR _11671_ sky130_fd_sc_hd__xor2_1
XFILLER_0_194_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput2 angle_in[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_1
X_19768_ _11602_ _11493_ net3135 VGND VGND VPWR VPWR _11603_ sky130_fd_sc_hd__a21o_1
XFILLER_0_190_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18719_ _10561_ net764 VGND VGND VPWR VPWR _10565_ sky130_fd_sc_hd__nand2_1
X_19699_ net3131 net3138 VGND VGND VPWR VPWR _11535_ sky130_fd_sc_hd__nor2_1
X_21730_ _01738_ _01739_ VGND VGND VPWR VPWR _01740_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21661_ _01660_ _01671_ VGND VGND VPWR VPWR _01672_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_143_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8209 net32 VGND VGND VPWR VPWR net8209 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23400_ _03201_ _03202_ _03203_ VGND VGND VPWR VPWR _03270_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20612_ _12362_ _12380_ _12392_ VGND VGND VPWR VPWR _12393_ sky130_fd_sc_hd__nor3_1
X_24380_ _04152_ _04160_ _04123_ VGND VGND VPWR VPWR _04239_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21592_ net1725 _01499_ _01495_ VGND VGND VPWR VPWR _01604_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_163_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire7508 net7509 VGND VGND VPWR VPWR net7508 sky130_fd_sc_hd__clkbuf_1
Xwire7519 net7520 VGND VGND VPWR VPWR net7519 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23331_ net5108 net4576 VGND VGND VPWR VPWR _03201_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20543_ net1822 net2082 net2084 net2079 VGND VGND VPWR VPWR _12328_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_28_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6818 net6815 VGND VGND VPWR VPWR net6818 sky130_fd_sc_hd__buf_1
XFILLER_0_7_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23262_ _03131_ _03123_ VGND VGND VPWR VPWR _03132_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20474_ net4054 _12262_ _12263_ net9216 VGND VGND VPWR VPWR _00500_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25001_ net4474 net5183 _04756_ VGND VGND VPWR VPWR _04758_ sky130_fd_sc_hd__nand3_1
X_22213_ _02216_ _02217_ VGND VGND VPWR VPWR _02218_ sky130_fd_sc_hd__xor2_1
XFILLER_0_131_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_18_Left_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23193_ _03037_ _03042_ VGND VGND VPWR VPWR _03063_ sky130_fd_sc_hd__xor2_1
XFILLER_0_131_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length1848 net1849 VGND VGND VPWR VPWR net1848 sky130_fd_sc_hd__buf_1
X_22144_ net5841 net5858 net2067 VGND VGND VPWR VPWR _02150_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22075_ _01975_ _01976_ _01973_ VGND VGND VPWR VPWR _02082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25903_ clknet_leaf_40_clk _00776_ net8769 VGND VGND VPWR VPWR pid_q.kp\[15\] sky130_fd_sc_hd__dfrtp_1
X_21026_ _01036_ _01041_ VGND VGND VPWR VPWR _01042_ sky130_fd_sc_hd__or2_1
Xwire1103 _07744_ VGND VGND VPWR VPWR net1103 sky130_fd_sc_hd__clkbuf_1
Xwire1114 net1115 VGND VGND VPWR VPWR net1114 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1125 _06218_ VGND VGND VPWR VPWR net1125 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1136 _05439_ VGND VGND VPWR VPWR net1136 sky130_fd_sc_hd__buf_1
XFILLER_0_57_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25834_ clknet_leaf_37_clk _00707_ net8745 VGND VGND VPWR VPWR pid_q.curr_error\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1147 _05045_ VGND VGND VPWR VPWR net1147 sky130_fd_sc_hd__buf_1
Xwire1158 _04548_ VGND VGND VPWR VPWR net1158 sky130_fd_sc_hd__clkbuf_1
Xwire1169 _02061_ VGND VGND VPWR VPWR net1169 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_27_Left_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22977_ _02856_ VGND VGND VPWR VPWR _00655_ sky130_fd_sc_hd__clkbuf_1
X_25765_ clknet_leaf_67_clk _00638_ net8453 VGND VGND VPWR VPWR pid_d.out\[6\] sky130_fd_sc_hd__dfrtp_1
X_24716_ net8022 _04546_ VGND VGND VPWR VPWR _04551_ sky130_fd_sc_hd__or2_1
X_12730_ _04984_ _04992_ VGND VGND VPWR VPWR _05003_ sky130_fd_sc_hd__xor2_1
X_21928_ _01934_ _01935_ VGND VGND VPWR VPWR _01936_ sky130_fd_sc_hd__xnor2_1
X_25696_ clknet_leaf_3_clk _00569_ net8575 VGND VGND VPWR VPWR pid_d.mult0.b\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout8615 net8634 VGND VGND VPWR VPWR net8615 sky130_fd_sc_hd__buf_1
X_12661_ _04927_ _04933_ VGND VGND VPWR VPWR _04934_ sky130_fd_sc_hd__xnor2_1
X_24647_ pid_q.prev_error\[15\] pid_q.curr_error\[15\] VGND VGND VPWR VPWR _04502_
+ sky130_fd_sc_hd__xnor2_1
X_21859_ _01867_ VGND VGND VPWR VPWR _01868_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14400_ net3647 VGND VGND VPWR VPWR _06603_ sky130_fd_sc_hd__buf_1
XFILLER_0_33_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout7914 net7918 VGND VGND VPWR VPWR net7914 sky130_fd_sc_hd__buf_1
Xwire8721 net8717 VGND VGND VPWR VPWR net8721 sky130_fd_sc_hd__dlymetal6s2s_1
X_12592_ net3016 VGND VGND VPWR VPWR _00006_ sky130_fd_sc_hd__clkbuf_1
X_15380_ _07310_ _07312_ VGND VGND VPWR VPWR _07454_ sky130_fd_sc_hd__nand2_1
Xmax_length5164 net5165 VGND VGND VPWR VPWR net5164 sky130_fd_sc_hd__clkbuf_1
X_24578_ _04347_ _04350_ net4919 VGND VGND VPWR VPWR _04434_ sky130_fd_sc_hd__a21o_1
Xwire8732 net8738 VGND VGND VPWR VPWR net8732 sky130_fd_sc_hd__buf_1
XFILLER_0_136_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length4430 pid_q.out\[9\] VGND VGND VPWR VPWR net4430 sky130_fd_sc_hd__buf_1
XFILLER_0_37_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8754 net8755 VGND VGND VPWR VPWR net8754 sky130_fd_sc_hd__buf_1
XFILLER_0_80_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire400 net401 VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__clkbuf_1
X_14331_ _06550_ VGND VGND VPWR VPWR _00069_ sky130_fd_sc_hd__clkbuf_1
X_23529_ net4795 _03396_ VGND VGND VPWR VPWR _03397_ sky130_fd_sc_hd__xnor2_1
Xwire8765 net8763 VGND VGND VPWR VPWR net8765 sky130_fd_sc_hd__buf_1
Xmax_length5197 matmul0.beta_pass\[14\] VGND VGND VPWR VPWR net5197 sky130_fd_sc_hd__buf_1
Xwire8776 net8777 VGND VGND VPWR VPWR net8776 sky130_fd_sc_hd__buf_1
XFILLER_0_52_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8787 net8788 VGND VGND VPWR VPWR net8787 sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_length4474 pid_q.out\[0\] VGND VGND VPWR VPWR net4474 sky130_fd_sc_hd__clkbuf_2
Xwire433 net434 VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__clkbuf_1
Xwire8798 net8800 VGND VGND VPWR VPWR net8798 sky130_fd_sc_hd__buf_1
Xwire444 net445 VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__clkbuf_1
X_14262_ net49 net2931 net2278 net9010 VGND VGND VPWR VPWR _00035_ sky130_fd_sc_hd__a22o_1
X_17050_ _08927_ _08929_ _08969_ VGND VGND VPWR VPWR _09009_ sky130_fd_sc_hd__mux2_1
Xwire455 net456 VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_36_Left_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire466 _03660_ VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire477 _01635_ VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__clkbuf_1
X_13213_ _05471_ _05477_ _05478_ _05485_ _05475_ VGND VGND VPWR VPWR _05486_ sky130_fd_sc_hd__o32ai_4
Xwire488 _11619_ VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__clkbuf_1
X_16001_ net3459 net2803 _07900_ net2224 net2829 VGND VGND VPWR VPWR _08069_ sky130_fd_sc_hd__o32a_1
Xmax_length3795 _01405_ VGND VGND VPWR VPWR net3795 sky130_fd_sc_hd__clkbuf_1
Xwire499 net500 VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__clkbuf_1
X_14193_ _06403_ VGND VGND VPWR VPWR _06453_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13144_ net7877 net1949 _05338_ net1947 net7909 VGND VGND VPWR VPWR _05417_ sky130_fd_sc_hd__a32o_1
XFILLER_0_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13075_ _05346_ net4255 VGND VGND VPWR VPWR _05348_ sky130_fd_sc_hd__and2_1
X_17952_ _09797_ _09799_ net3239 net3238 VGND VGND VPWR VPWR _09803_ sky130_fd_sc_hd__o211a_1
Xwire3050 net3051 VGND VGND VPWR VPWR net3050 sky130_fd_sc_hd__clkbuf_1
Xwire3061 net3062 VGND VGND VPWR VPWR net3061 sky130_fd_sc_hd__buf_1
X_16903_ cordic0.slte0.opA\[9\] _08866_ net6404 VGND VGND VPWR VPWR _08867_ sky130_fd_sc_hd__o21bai_1
Xwire3072 net3073 VGND VGND VPWR VPWR net3072 sky130_fd_sc_hd__buf_1
X_17883_ net1214 _09733_ VGND VGND VPWR VPWR _09734_ sky130_fd_sc_hd__xor2_1
Xwire3083 net3084 VGND VGND VPWR VPWR net3083 sky130_fd_sc_hd__buf_1
Xwire3094 net3095 VGND VGND VPWR VPWR net3094 sky130_fd_sc_hd__clkbuf_2
Xwire2360 net2361 VGND VGND VPWR VPWR net2360 sky130_fd_sc_hd__buf_1
X_19622_ net3186 _10918_ _11401_ VGND VGND VPWR VPWR _11459_ sky130_fd_sc_hd__a21o_1
Xwire2371 net2372 VGND VGND VPWR VPWR net2371 sky130_fd_sc_hd__clkbuf_1
X_16834_ net6425 matmul0.sin\[5\] net3366 VGND VGND VPWR VPWR _08808_ sky130_fd_sc_hd__mux2_1
Xwire2382 _00011_ VGND VGND VPWR VPWR net2382 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_45_Left_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_189_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2393 _04850_ VGND VGND VPWR VPWR net2393 sky130_fd_sc_hd__clkbuf_2
Xwire1670 net1671 VGND VGND VPWR VPWR net1670 sky130_fd_sc_hd__clkbuf_2
X_19553_ _11380_ _11389_ VGND VGND VPWR VPWR _11390_ sky130_fd_sc_hd__xnor2_1
Xwire1681 net1682 VGND VGND VPWR VPWR net1681 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_87_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16765_ matmul0.a_in\[2\] matmul0.a\[2\] net3378 VGND VGND VPWR VPWR _08772_ sky130_fd_sc_hd__mux2_1
X_13977_ _06191_ _06196_ _06241_ VGND VGND VPWR VPWR _06242_ sky130_fd_sc_hd__o21ai_2
Xwire1692 net1693 VGND VGND VPWR VPWR net1692 sky130_fd_sc_hd__clkbuf_1
X_18504_ net2540 _10290_ _10351_ VGND VGND VPWR VPWR _10353_ sky130_fd_sc_hd__or3b_1
X_15716_ net3574 net3570 net4095 net4094 VGND VGND VPWR VPWR _07787_ sky130_fd_sc_hd__o22a_1
XFILLER_0_158_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12928_ net1006 net1005 _05119_ _05120_ VGND VGND VPWR VPWR _05201_ sky130_fd_sc_hd__o211a_1
X_19484_ net6359 _11264_ _11319_ _11320_ net6267 VGND VGND VPWR VPWR _11321_ sky130_fd_sc_hd__o2111a_1
X_16696_ _08724_ _08725_ VGND VGND VPWR VPWR _08726_ sky130_fd_sc_hd__xnor2_1
X_18435_ net6897 net6921 VGND VGND VPWR VPWR _10285_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15647_ _07570_ net3405 net2666 net2776 net2781 VGND VGND VPWR VPWR _07719_ sky130_fd_sc_hd__a221o_1
X_12859_ net2310 net1955 VGND VGND VPWR VPWR _05132_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18366_ _10206_ _10216_ VGND VGND VPWR VPWR _10217_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_111_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15578_ _07648_ _07649_ VGND VGND VPWR VPWR _07650_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17317_ net7806 _09208_ VGND VGND VPWR VPWR _09231_ sky130_fd_sc_hd__nand2_1
X_14529_ net7279 VGND VGND VPWR VPWR _06708_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_54_Left_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18297_ net815 _10147_ VGND VGND VPWR VPWR _10148_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17248_ net2164 net257 net1799 net9140 VGND VGND VPWR VPWR _00346_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17179_ net1475 _09130_ net3323 VGND VGND VPWR VPWR _09131_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20190_ net243 _12015_ VGND VGND VPWR VPWR _12016_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_179_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_63_Left_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22900_ net4370 net3761 VGND VGND VPWR VPWR _02793_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23880_ _03743_ _03744_ VGND VGND VPWR VPWR _03745_ sky130_fd_sc_hd__xor2_1
X_22831_ net4354 net553 _02731_ net4335 net2463 VGND VGND VPWR VPWR _02732_ sky130_fd_sc_hd__a221o_1
XFILLER_0_195_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22762_ net4303 net8946 VGND VGND VPWR VPWR _02686_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25550_ clknet_leaf_66_clk _00012_ net8647 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_155_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24501_ net4555 VGND VGND VPWR VPWR _04358_ sky130_fd_sc_hd__inv_2
X_21713_ _01626_ _01722_ _01723_ VGND VGND VPWR VPWR _01724_ sky130_fd_sc_hd__and3_1
X_25481_ clknet_leaf_45_clk _00361_ net8789 VGND VGND VPWR VPWR svm0.tA\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22693_ pid_d.ki\[8\] net2445 net3000 pid_d.kp\[8\] VGND VGND VPWR VPWR _02637_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8006 pid_q.target\[6\] VGND VGND VPWR VPWR net8006 sky130_fd_sc_hd__clkbuf_1
Xwire8017 net8018 VGND VGND VPWR VPWR net8017 sky130_fd_sc_hd__clkbuf_2
X_24432_ net4872 VGND VGND VPWR VPWR _04290_ sky130_fd_sc_hd__inv_2
X_21644_ _01570_ _01581_ net1722 VGND VGND VPWR VPWR _01655_ sky130_fd_sc_hd__a21bo_1
Xwire8028 net8029 VGND VGND VPWR VPWR net8028 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_136_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8039 net8040 VGND VGND VPWR VPWR net8039 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24363_ net2020 net1653 net2409 VGND VGND VPWR VPWR _04222_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3003 net3004 VGND VGND VPWR VPWR net3003 sky130_fd_sc_hd__buf_1
XFILLER_0_170_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21575_ net5851 net5423 VGND VGND VPWR VPWR _01587_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7327 matmul0.alpha_pass\[4\] VGND VGND VPWR VPWR net7327 sky130_fd_sc_hd__clkbuf_1
Xwire7338 net7339 VGND VGND VPWR VPWR net7338 sky130_fd_sc_hd__clkbuf_1
Xwire6604 net6605 VGND VGND VPWR VPWR net6604 sky130_fd_sc_hd__clkbuf_1
Xwire7349 net7350 VGND VGND VPWR VPWR net7349 sky130_fd_sc_hd__clkbuf_1
X_23314_ _02956_ _02959_ _02953_ VGND VGND VPWR VPWR _03184_ sky130_fd_sc_hd__o21ba_1
Xmax_length3047 net3048 VGND VGND VPWR VPWR net3047 sky130_fd_sc_hd__clkbuf_1
Xfanout5819 net5827 VGND VGND VPWR VPWR net5819 sky130_fd_sc_hd__buf_1
X_20526_ net6823 net6767 net6502 VGND VGND VPWR VPWR _12312_ sky130_fd_sc_hd__mux2_1
Xwire6615 net6613 VGND VGND VPWR VPWR net6615 sky130_fd_sc_hd__buf_1
X_24294_ net4580 net4590 net3053 VGND VGND VPWR VPWR _04154_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6637 net6632 VGND VGND VPWR VPWR net6637 sky130_fd_sc_hd__clkbuf_1
Xwire6648 matmul0.matmul_stage_inst.state\[1\] VGND VGND VPWR VPWR net6648 sky130_fd_sc_hd__buf_1
Xwire6659 net6656 VGND VGND VPWR VPWR net6659 sky130_fd_sc_hd__buf_1
XFILLER_0_132_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2346 net2347 VGND VGND VPWR VPWR net2346 sky130_fd_sc_hd__buf_1
XFILLER_0_105_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5914 net5915 VGND VGND VPWR VPWR net5914 sky130_fd_sc_hd__buf_1
X_23245_ _03020_ _03022_ _03021_ VGND VGND VPWR VPWR _03115_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5925 net5926 VGND VGND VPWR VPWR net5925 sky130_fd_sc_hd__clkbuf_1
X_20457_ net3667 net967 net2607 VGND VGND VPWR VPWR _12249_ sky130_fd_sc_hd__o21a_1
XFILLER_0_63_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length1634 net1635 VGND VGND VPWR VPWR net1634 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5947 net5941 VGND VGND VPWR VPWR net5947 sky130_fd_sc_hd__clkbuf_1
Xmax_length1645 net1646 VGND VGND VPWR VPWR net1645 sky130_fd_sc_hd__buf_1
Xwire5969 pid_d.curr_error\[5\] VGND VGND VPWR VPWR net5969 sky130_fd_sc_hd__buf_1
X_23176_ _03026_ _03044_ _03045_ VGND VGND VPWR VPWR _03046_ sky130_fd_sc_hd__and3_1
XFILLER_0_113_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20388_ _12182_ net603 VGND VGND VPWR VPWR _12187_ sky130_fd_sc_hd__and2_1
X_22127_ _02129_ _02132_ VGND VGND VPWR VPWR _02133_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_24_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22058_ net1710 _02060_ _02061_ VGND VGND VPWR VPWR _02065_ sky130_fd_sc_hd__or3_1
XFILLER_0_27_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13900_ net839 _06110_ _06105_ VGND VGND VPWR VPWR _06166_ sky130_fd_sc_hd__a21bo_1
X_21009_ net1185 _01024_ VGND VGND VPWR VPWR _01025_ sky130_fd_sc_hd__nand2_1
X_14880_ matmul0.b\[12\] matmul0.matmul_stage_inst.f\[12\] net3604 VGND VGND VPWR
+ VPWR _06958_ sky130_fd_sc_hd__mux2_1
X_13831_ _06036_ _06037_ _06097_ VGND VGND VPWR VPWR _06098_ sky130_fd_sc_hd__a21o_1
X_25817_ clknet_leaf_37_clk _00690_ net8746 VGND VGND VPWR VPWR pid_q.prev_error\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16550_ _08555_ _08556_ _08557_ VGND VGND VPWR VPWR _08609_ sky130_fd_sc_hd__a21o_1
X_13762_ net7789 net2948 net1940 _06028_ net3676 VGND VGND VPWR VPWR _06030_ sky130_fd_sc_hd__a311o_1
X_25748_ clknet_leaf_9_clk _00621_ net8601 VGND VGND VPWR VPWR pid_d.kp\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15501_ net4111 net4108 net4079 net4077 VGND VGND VPWR VPWR _07574_ sky130_fd_sc_hd__o22a_1
XFILLER_0_168_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12713_ net7882 net2356 net1978 VGND VGND VPWR VPWR _04986_ sky130_fd_sc_hd__and3_1
XFILLER_0_195_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16481_ _08499_ _08541_ VGND VGND VPWR VPWR _08542_ sky130_fd_sc_hd__nor2_1
Xfanout8401 net8408 VGND VGND VPWR VPWR net8401 sky130_fd_sc_hd__buf_1
X_13693_ net7621 net1605 VGND VGND VPWR VPWR _05962_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25679_ clknet_leaf_1_clk _00552_ net8405 VGND VGND VPWR VPWR pid_d.curr_error\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout8423 net8521 VGND VGND VPWR VPWR net8423 sky130_fd_sc_hd__buf_1
X_18220_ _10062_ _10070_ VGND VGND VPWR VPWR _10071_ sky130_fd_sc_hd__xor2_1
Xfanout7700 net7708 VGND VGND VPWR VPWR net7700 sky130_fd_sc_hd__clkbuf_1
X_15432_ net3450 net2690 VGND VGND VPWR VPWR _07506_ sky130_fd_sc_hd__nor2_1
Xfanout8445 net8480 VGND VGND VPWR VPWR net8445 sky130_fd_sc_hd__buf_1
Xfanout7711 svm0.periodTop\[10\] VGND VGND VPWR VPWR net7711 sky130_fd_sc_hd__clkbuf_1
X_12644_ net7341 net3030 net3695 VGND VGND VPWR VPWR _04917_ sky130_fd_sc_hd__nand3_1
XFILLER_0_150_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout7722 net7730 VGND VGND VPWR VPWR net7722 sky130_fd_sc_hd__buf_1
XFILLER_0_109_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18151_ _09998_ net3234 _09956_ VGND VGND VPWR VPWR _10002_ sky130_fd_sc_hd__o21ba_1
Xwire8540 net8541 VGND VGND VPWR VPWR net8540 sky130_fd_sc_hd__buf_1
Xfanout7755 net7774 VGND VGND VPWR VPWR net7755 sky130_fd_sc_hd__clkbuf_1
X_15363_ _07426_ _07436_ VGND VGND VPWR VPWR _07437_ sky130_fd_sc_hd__xnor2_1
X_12575_ matmul0.matmul_stage_inst.start VGND VGND VPWR VPWR _04863_ sky130_fd_sc_hd__inv_2
Xwire8562 net8561 VGND VGND VPWR VPWR net8562 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_124_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout7777 net7797 VGND VGND VPWR VPWR net7777 sky130_fd_sc_hd__buf_1
X_17102_ net1505 _09058_ VGND VGND VPWR VPWR _09059_ sky130_fd_sc_hd__or2_1
Xwire230 net231 VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__clkbuf_1
X_14314_ net6443 _06535_ VGND VGND VPWR VPWR _06536_ sky130_fd_sc_hd__nor2_1
Xwire241 net242 VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__buf_1
Xwire8595 net8596 VGND VGND VPWR VPWR net8595 sky130_fd_sc_hd__clkbuf_1
Xwire7850 net7844 VGND VGND VPWR VPWR net7850 sky130_fd_sc_hd__buf_1
XFILLER_0_29_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18082_ net3257 net3264 _09849_ VGND VGND VPWR VPWR _09933_ sky130_fd_sc_hd__mux2_1
Xwire7861 net7868 VGND VGND VPWR VPWR net7861 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15294_ net3602 VGND VGND VPWR VPWR _07368_ sky130_fd_sc_hd__buf_1
Xwire252 net253 VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__clkbuf_1
Xwire7872 svm0.periodTop\[3\] VGND VGND VPWR VPWR net7872 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire263 _04402_ VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__buf_1
XFILLER_0_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7883 net7880 VGND VGND VPWR VPWR net7883 sky130_fd_sc_hd__buf_1
XFILLER_0_180_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7894 net7898 VGND VGND VPWR VPWR net7894 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17033_ net1077 VGND VGND VPWR VPWR _08993_ sky130_fd_sc_hd__buf_1
Xwire274 _11958_ VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__buf_1
Xwire285 net286 VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__buf_1
X_14245_ _06499_ net7535 VGND VGND VPWR VPWR _06500_ sky130_fd_sc_hd__nand2_1
Xwire296 net297 VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14176_ _06395_ _06421_ _06424_ _06435_ VGND VGND VPWR VPWR _06436_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13127_ _05398_ _05399_ VGND VGND VPWR VPWR _05400_ sky130_fd_sc_hd__or2_1
X_18984_ _10820_ VGND VGND VPWR VPWR _10821_ sky130_fd_sc_hd__buf_1
XFILLER_0_178_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13058_ _05204_ net790 _05208_ VGND VGND VPWR VPWR _05331_ sky130_fd_sc_hd__or3_1
X_17935_ _09780_ _09784_ _09785_ VGND VGND VPWR VPWR _09786_ sky130_fd_sc_hd__o21ba_1
X_17866_ _09622_ _09623_ _08966_ VGND VGND VPWR VPWR _09717_ sky130_fd_sc_hd__mux2_1
Xwire2190 net2191 VGND VGND VPWR VPWR net2190 sky130_fd_sc_hd__buf_1
X_19605_ net1418 _11403_ net1417 VGND VGND VPWR VPWR _11442_ sky130_fd_sc_hd__a21bo_1
X_16817_ net9210 matmul0.cos\[11\] net3368 VGND VGND VPWR VPWR _08799_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17797_ net7095 VGND VGND VPWR VPWR _09648_ sky130_fd_sc_hd__inv_2
XFILLER_0_177_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19536_ net1060 _11342_ _11372_ VGND VGND VPWR VPWR _11373_ sky130_fd_sc_hd__o21a_1
X_16748_ net7564 matmul0.b\[10\] net3380 VGND VGND VPWR VPWR _08763_ sky130_fd_sc_hd__mux2_1
X_19467_ net1064 _11019_ _11020_ _11018_ VGND VGND VPWR VPWR _11304_ sky130_fd_sc_hd__a31o_1
XFILLER_0_158_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16679_ _08710_ _08706_ matmul0.matmul_stage_inst.mult2\[8\] VGND VGND VPWR VPWR
+ _08711_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_146_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18418_ _10217_ net1210 _10245_ VGND VGND VPWR VPWR _10268_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_115_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19398_ _11234_ _11196_ _11198_ _11199_ VGND VGND VPWR VPWR _11235_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18349_ _10147_ _10074_ _10075_ VGND VGND VPWR VPWR _10200_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_12_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21360_ net5811 net5495 VGND VGND VPWR VPWR _01374_ sky130_fd_sc_hd__nand2_1
XFILLER_0_185_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20311_ net1491 _12115_ net3317 VGND VGND VPWR VPWR _12116_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput60 currT_in[5] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_1
X_21291_ _00819_ _00820_ _01305_ VGND VGND VPWR VPWR _01306_ sky130_fd_sc_hd__a21oi_2
Xinput71 periodTop[15] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput82 pid_d_addr[10] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_1
Xwire4509 net4510 VGND VGND VPWR VPWR net4509 sky130_fd_sc_hd__buf_1
XFILLER_0_40_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput93 pid_d_addr[6] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_1
X_23030_ net4968 net4740 VGND VGND VPWR VPWR _02900_ sky130_fd_sc_hd__nand2_1
XFILLER_0_142_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20242_ net12 net13 _12050_ net8122 VGND VGND VPWR VPWR _12058_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3808 net3809 VGND VGND VPWR VPWR net3808 sky130_fd_sc_hd__clkbuf_1
Xwire3819 net3820 VGND VGND VPWR VPWR net3819 sky130_fd_sc_hd__clkbuf_1
X_20173_ _11348_ _11588_ net3128 net6067 net6088 VGND VGND VPWR VPWR _11999_ sky130_fd_sc_hd__o221a_1
X_24981_ _04745_ VGND VGND VPWR VPWR _00770_ sky130_fd_sc_hd__clkbuf_1
X_23932_ _03688_ _03691_ _03685_ VGND VGND VPWR VPWR _03796_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23863_ _03724_ _03726_ VGND VGND VPWR VPWR _03728_ sky130_fd_sc_hd__and2_1
XFILLER_0_169_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length7803 net7804 VGND VGND VPWR VPWR net7803 sky130_fd_sc_hd__buf_1
XFILLER_0_54_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25602_ clknet_leaf_106_clk _00475_ net8355 VGND VGND VPWR VPWR cordic0.slte0.opB\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_22814_ net5986 net3759 VGND VGND VPWR VPWR _02717_ sky130_fd_sc_hd__nand2_1
X_23794_ _03586_ _03659_ VGND VGND VPWR VPWR _03660_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_168_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25533_ clknet_leaf_35_clk _00413_ net8765 VGND VGND VPWR VPWR svm0.ready sky130_fd_sc_hd__dfstp_1
XFILLER_0_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22745_ pid_d.ki\[6\] _02674_ net1689 VGND VGND VPWR VPWR _02675_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25464_ clknet_leaf_53_clk _00344_ net8807 VGND VGND VPWR VPWR svm0.tB\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_149_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22676_ _02625_ net5620 net2448 VGND VGND VPWR VPWR _02626_ sky130_fd_sc_hd__mux2_1
Xfanout7018 net7024 VGND VGND VPWR VPWR net7018 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24415_ net4537 net4555 net3054 VGND VGND VPWR VPWR _04273_ sky130_fd_sc_hd__and3_1
Xwire7102 cordic0.vec\[1\]\[3\] VGND VGND VPWR VPWR net7102 sky130_fd_sc_hd__buf_1
X_21627_ pid_d.prev_error\[4\] pid_d.curr_error\[4\] VGND VGND VPWR VPWR _01639_ sky130_fd_sc_hd__xnor2_1
Xwire7113 net7110 VGND VGND VPWR VPWR net7113 sky130_fd_sc_hd__buf_1
Xfanout6306 cordic0.vec\[0\]\[3\] VGND VGND VPWR VPWR net6306 sky130_fd_sc_hd__buf_1
X_25395_ clknet_leaf_74_clk _00278_ net8498 VGND VGND VPWR VPWR matmul0.b\[14\] sky130_fd_sc_hd__dfrtp_1
Xwire7124 net7122 VGND VGND VPWR VPWR net7124 sky130_fd_sc_hd__buf_2
XFILLER_0_8_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6401 cordic0.slte0.opB\[12\] VGND VGND VPWR VPWR net6401 sky130_fd_sc_hd__clkbuf_1
Xwire7146 net7143 VGND VGND VPWR VPWR net7146 sky130_fd_sc_hd__buf_1
X_24346_ _04131_ _04133_ _04132_ VGND VGND VPWR VPWR _04205_ sky130_fd_sc_hd__o21ai_1
X_21558_ _01454_ _01459_ _01569_ VGND VGND VPWR VPWR _01570_ sky130_fd_sc_hd__o21a_1
Xwire6412 cordic0.slte0.opB\[7\] VGND VGND VPWR VPWR net6412 sky130_fd_sc_hd__buf_1
Xwire7168 matmul0.cos\[11\] VGND VGND VPWR VPWR net7168 sky130_fd_sc_hd__buf_1
Xwire6423 cordic0.sin\[8\] VGND VGND VPWR VPWR net6423 sky130_fd_sc_hd__clkbuf_1
Xwire6434 net6435 VGND VGND VPWR VPWR net6434 sky130_fd_sc_hd__clkbuf_1
Xwire7179 matmul0.cos\[5\] VGND VGND VPWR VPWR net7179 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5700 pid_d.mult0.b\[13\] VGND VGND VPWR VPWR net5700 sky130_fd_sc_hd__clkbuf_1
Xwire6445 net6446 VGND VGND VPWR VPWR net6445 sky130_fd_sc_hd__buf_1
X_20509_ net6917 net6890 net6904 net6871 net6491 net6521 VGND VGND VPWR VPWR _12296_
+ sky130_fd_sc_hd__mux4_1
X_24277_ _04128_ _04136_ VGND VGND VPWR VPWR _04137_ sky130_fd_sc_hd__xnor2_2
Xwire5711 net5706 VGND VGND VPWR VPWR net5711 sky130_fd_sc_hd__buf_1
Xwire6456 net6455 VGND VGND VPWR VPWR net6456 sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_length2154 net2155 VGND VGND VPWR VPWR net2154 sky130_fd_sc_hd__clkbuf_1
Xwire5722 net5723 VGND VGND VPWR VPWR net5722 sky130_fd_sc_hd__clkbuf_1
X_21489_ net1180 _01501_ VGND VGND VPWR VPWR _01502_ sky130_fd_sc_hd__xor2_1
Xwire5733 net5734 VGND VGND VPWR VPWR net5733 sky130_fd_sc_hd__clkbuf_1
X_14030_ net7604 net1332 VGND VGND VPWR VPWR _06294_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23228_ net5143 net4631 VGND VGND VPWR VPWR _03098_ sky130_fd_sc_hd__nand2_1
Xwire6489 net6490 VGND VGND VPWR VPWR net6489 sky130_fd_sc_hd__clkbuf_2
Xwire5755 net5756 VGND VGND VPWR VPWR net5755 sky130_fd_sc_hd__clkbuf_1
Xwire5788 net5789 VGND VGND VPWR VPWR net5788 sky130_fd_sc_hd__buf_1
XFILLER_0_28_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5799 net5801 VGND VGND VPWR VPWR net5799 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_28_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23159_ net5013 net4776 VGND VGND VPWR VPWR _03029_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15981_ net1520 _08048_ VGND VGND VPWR VPWR _08049_ sky130_fd_sc_hd__xnor2_2
X_17720_ net9201 net1456 net1789 net5177 VGND VGND VPWR VPWR _00425_ sky130_fd_sc_hd__a22o_1
X_14932_ _06996_ _07005_ VGND VGND VPWR VPWR _07006_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17651_ net6704 svm0.tA\[11\] VGND VGND VPWR VPWR _09531_ sky130_fd_sc_hd__nand2_1
X_14863_ net7186 matmul0.matmul_stage_inst.f\[4\] _06939_ VGND VGND VPWR VPWR _06949_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16602_ matmul0.matmul_stage_inst.mult2\[8\] net311 net2618 VGND VGND VPWR VPWR _08651_
+ sky130_fd_sc_hd__mux2_1
X_13814_ _06081_ VGND VGND VPWR VPWR _06082_ sky130_fd_sc_hd__inv_2
X_17582_ _09449_ _09463_ _09444_ VGND VGND VPWR VPWR _09464_ sky130_fd_sc_hd__a21oi_1
X_14794_ net9052 net3006 _06913_ VGND VGND VPWR VPWR _00169_ sky130_fd_sc_hd__o21a_1
XFILLER_0_85_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19321_ net6312 net3203 _10823_ _11140_ _11147_ VGND VGND VPWR VPWR _11158_ sky130_fd_sc_hd__a221o_1
X_16533_ matmul0.matmul_stage_inst.mult1\[14\] net167 net3474 VGND VGND VPWR VPWR
+ _08593_ sky130_fd_sc_hd__mux2_1
X_13745_ _05872_ net451 VGND VGND VPWR VPWR _06013_ sky130_fd_sc_hd__nor2_1
XFILLER_0_168_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_196_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19252_ _11028_ _11088_ VGND VGND VPWR VPWR _11089_ sky130_fd_sc_hd__xnor2_1
X_16464_ _08449_ _08451_ VGND VGND VPWR VPWR _08525_ sky130_fd_sc_hd__nor2_1
XFILLER_0_195_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13676_ _05943_ _05944_ VGND VGND VPWR VPWR _05945_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18203_ _10038_ _10053_ VGND VGND VPWR VPWR _10054_ sky130_fd_sc_hd__xnor2_1
X_15415_ _07488_ VGND VGND VPWR VPWR _07489_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12627_ _04895_ net2367 VGND VGND VPWR VPWR _04900_ sky130_fd_sc_hd__and2_1
X_19183_ net3187 _11017_ _10935_ VGND VGND VPWR VPWR _11020_ sky130_fd_sc_hd__or3_1
X_16395_ net3402 net2642 VGND VGND VPWR VPWR _08457_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8370 net8371 VGND VGND VPWR VPWR net8370 sky130_fd_sc_hd__clkbuf_1
X_18134_ _09977_ net1778 _09984_ net962 VGND VGND VPWR VPWR _09985_ sky130_fd_sc_hd__a211o_1
X_15346_ net3528 net2801 VGND VGND VPWR VPWR _07420_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8392 net8393 VGND VGND VPWR VPWR net8392 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7680 net7681 VGND VGND VPWR VPWR net7680 sky130_fd_sc_hd__dlymetal6s2s_1
X_18065_ net7007 _09915_ VGND VGND VPWR VPWR _09916_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_80_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout6895 net6902 VGND VGND VPWR VPWR net6895 sky130_fd_sc_hd__buf_1
X_15277_ net6622 net6639 net7381 VGND VGND VPWR VPWR _07351_ sky130_fd_sc_hd__o21a_1
Xhold107 pid_q.target\[7\] VGND VGND VPWR VPWR net9060 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold118 matmul0.matmul_stage_inst.c\[1\] VGND VGND VPWR VPWR net9071 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17016_ net1804 _08976_ VGND VGND VPWR VPWR _08977_ sky130_fd_sc_hd__xnor2_2
Xhold129 matmul0.matmul_stage_inst.b\[10\] VGND VGND VPWR VPWR net9082 sky130_fd_sc_hd__dlygate4sd3_1
X_14228_ _06446_ _06470_ _06485_ VGND VGND VPWR VPWR _06486_ sky130_fd_sc_hd__a21o_1
Xwire6990 net6991 VGND VGND VPWR VPWR net6990 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_145_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14159_ _06402_ _06419_ VGND VGND VPWR VPWR _06420_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18967_ net6232 net6249 VGND VGND VPWR VPWR _10804_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17918_ _09767_ _09768_ _09629_ VGND VGND VPWR VPWR _09769_ sky130_fd_sc_hd__a21o_1
X_18898_ _10718_ _10719_ _10713_ VGND VGND VPWR VPWR _10739_ sky130_fd_sc_hd__mux2_1
X_17849_ _09688_ _09699_ VGND VGND VPWR VPWR _09700_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_179_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20860_ _00860_ _00875_ VGND VGND VPWR VPWR _00876_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_178_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19519_ _11294_ _11354_ VGND VGND VPWR VPWR _11356_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20791_ net5637 net5702 VGND VGND VPWR VPWR _12562_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22530_ net9135 net1699 _02527_ VGND VGND VPWR VPWR _00537_ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22461_ pid_d.prev_error\[15\] net5964 VGND VGND VPWR VPWR _02462_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24200_ net4553 net4867 VGND VGND VPWR VPWR _04061_ sky130_fd_sc_hd__nand2_1
X_21412_ _01342_ _01425_ VGND VGND VPWR VPWR _01426_ sky130_fd_sc_hd__xor2_1
XFILLER_0_173_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25180_ clknet_leaf_68_clk _00069_ net8452 VGND VGND VPWR VPWR matmul0.a_in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_22392_ _02393_ _02394_ net4364 VGND VGND VPWR VPWR _02395_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24131_ _03991_ _03992_ VGND VGND VPWR VPWR _03993_ sky130_fd_sc_hd__or2b_1
Xwire5007 net4999 VGND VGND VPWR VPWR net5007 sky130_fd_sc_hd__clkbuf_1
X_21343_ _01351_ _01353_ _01356_ VGND VGND VPWR VPWR _01357_ sky130_fd_sc_hd__and3_1
Xwire5018 net5020 VGND VGND VPWR VPWR net5018 sky130_fd_sc_hd__clkbuf_1
Xwire5029 net5030 VGND VGND VPWR VPWR net5029 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24062_ net4790 _03924_ VGND VGND VPWR VPWR _03925_ sky130_fd_sc_hd__xnor2_1
Xwire4306 net4307 VGND VGND VPWR VPWR net4306 sky130_fd_sc_hd__clkbuf_1
X_21274_ net3842 _00856_ VGND VGND VPWR VPWR _01289_ sky130_fd_sc_hd__nor2_1
Xwire4328 net4329 VGND VGND VPWR VPWR net4328 sky130_fd_sc_hd__buf_1
Xwire4339 net4334 VGND VGND VPWR VPWR net4339 sky130_fd_sc_hd__clkbuf_1
X_23013_ net5141 net4595 VGND VGND VPWR VPWR _02883_ sky130_fd_sc_hd__nand2_1
X_20225_ net10 _12044_ VGND VGND VPWR VPWR _12045_ sky130_fd_sc_hd__xnor2_1
Xwire3616 _06862_ VGND VGND VPWR VPWR net3616 sky130_fd_sc_hd__buf_1
Xwire3627 net3628 VGND VGND VPWR VPWR net3627 sky130_fd_sc_hd__buf_1
Xwire3638 net3639 VGND VGND VPWR VPWR net3638 sky130_fd_sc_hd__clkbuf_1
Xwire2904 net2905 VGND VGND VPWR VPWR net2904 sky130_fd_sc_hd__clkbuf_1
Xwire3649 net3650 VGND VGND VPWR VPWR net3649 sky130_fd_sc_hd__buf_1
Xwire2915 net2916 VGND VGND VPWR VPWR net2915 sky130_fd_sc_hd__buf_1
X_20156_ _11979_ _11982_ _11934_ VGND VGND VPWR VPWR _11983_ sky130_fd_sc_hd__mux2_1
Xwire2926 net2927 VGND VGND VPWR VPWR net2926 sky130_fd_sc_hd__clkbuf_1
Xwire2937 net2938 VGND VGND VPWR VPWR net2937 sky130_fd_sc_hd__clkbuf_2
Xwire2948 net2949 VGND VGND VPWR VPWR net2948 sky130_fd_sc_hd__buf_1
Xwire2959 net2960 VGND VGND VPWR VPWR net2959 sky130_fd_sc_hd__buf_1
X_24964_ pid_q.kp\[1\] _04704_ _04735_ VGND VGND VPWR VPWR _04737_ sky130_fd_sc_hd__mux2_1
X_20087_ _11844_ _11873_ VGND VGND VPWR VPWR _11916_ sky130_fd_sc_hd__nor2_1
X_23915_ _03748_ _03755_ VGND VGND VPWR VPWR _03779_ sky130_fd_sc_hd__or2_1
X_24895_ pid_q.ki\[13\] net3711 net3701 pid_q.kp\[13\] VGND VGND VPWR VPWR _04688_
+ sky130_fd_sc_hd__a22o_1
Xmax_length8345 net8346 VGND VGND VPWR VPWR net8345 sky130_fd_sc_hd__buf_1
Xmax_length8356 net8353 VGND VGND VPWR VPWR net8356 sky130_fd_sc_hd__clkbuf_2
X_23846_ _03709_ _03710_ VGND VGND VPWR VPWR _03711_ sky130_fd_sc_hd__xor2_2
XFILLER_0_196_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23777_ net1666 _03507_ _03642_ VGND VGND VPWR VPWR _03643_ sky130_fd_sc_hd__a21o_1
X_20989_ net2482 _00878_ VGND VGND VPWR VPWR _01005_ sky130_fd_sc_hd__xor2_1
XFILLER_0_178_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length7688 net7689 VGND VGND VPWR VPWR net7688 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25516_ clknet_leaf_44_clk _00396_ net8785 VGND VGND VPWR VPWR svm0.counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13530_ net912 net997 VGND VGND VPWR VPWR _05801_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22728_ _02663_ VGND VGND VPWR VPWR _00599_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13461_ _05732_ _05733_ VGND VGND VPWR VPWR _05734_ sky130_fd_sc_hd__xor2_1
X_25447_ clknet_leaf_114_clk _00330_ net8334 VGND VGND VPWR VPWR cordic0.vec\[1\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22659_ net5712 net3085 net294 net8888 VGND VGND VPWR VPWR _00579_ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_173_Right_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15200_ _07095_ net3508 VGND VGND VPWR VPWR _07274_ sky130_fd_sc_hd__or2_1
XFILLER_0_180_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16180_ net672 _08222_ _08244_ VGND VGND VPWR VPWR _08245_ sky130_fd_sc_hd__o21ai_2
X_13392_ net684 _05664_ _05307_ VGND VGND VPWR VPWR _05665_ sky130_fd_sc_hd__a21o_1
X_25378_ clknet_leaf_63_clk _00261_ net8667 VGND VGND VPWR VPWR matmul0.alpha_pass\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout5413 net5419 VGND VGND VPWR VPWR net5413 sky130_fd_sc_hd__clkbuf_1
Xfanout6169 net6193 VGND VGND VPWR VPWR net6169 sky130_fd_sc_hd__clkbuf_2
Xwire6231 net6232 VGND VGND VPWR VPWR net6231 sky130_fd_sc_hd__clkbuf_1
X_15131_ net3465 VGND VGND VPWR VPWR _07205_ sky130_fd_sc_hd__clkbuf_1
Xfanout4701 pid_q.mult0.a\[4\] VGND VGND VPWR VPWR net4701 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24329_ _04187_ _04174_ net3736 VGND VGND VPWR VPWR _04188_ sky130_fd_sc_hd__o21a_1
XFILLER_0_90_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout4734 net4745 VGND VGND VPWR VPWR net4734 sky130_fd_sc_hd__buf_1
Xwire5530 net5531 VGND VGND VPWR VPWR net5530 sky130_fd_sc_hd__clkbuf_1
X_15062_ net6618 net6639 VGND VGND VPWR VPWR _07136_ sky130_fd_sc_hd__or2_1
Xwire5552 net5553 VGND VGND VPWR VPWR net5552 sky130_fd_sc_hd__buf_1
X_14013_ net282 net319 VGND VGND VPWR VPWR _06277_ sky130_fd_sc_hd__nand2_1
Xwire5574 net5568 VGND VGND VPWR VPWR net5574 sky130_fd_sc_hd__buf_1
Xwire4851 net4852 VGND VGND VPWR VPWR net4851 sky130_fd_sc_hd__buf_1
XFILLER_0_102_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19870_ net3292 _11699_ _11701_ net6043 _11702_ VGND VGND VPWR VPWR _11703_ sky130_fd_sc_hd__o221a_1
XFILLER_0_102_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4873 net4871 VGND VGND VPWR VPWR net4873 sky130_fd_sc_hd__buf_1
Xwire4884 net4879 VGND VGND VPWR VPWR net4884 sky130_fd_sc_hd__clkbuf_1
X_18821_ _10661_ _10663_ VGND VGND VPWR VPWR _10664_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18752_ net6779 net6795 VGND VGND VPWR VPWR _10597_ sky130_fd_sc_hd__nand2_1
X_15964_ _08023_ _08031_ VGND VGND VPWR VPWR _08032_ sky130_fd_sc_hd__xnor2_1
X_17703_ _09578_ VGND VGND VPWR VPWR _09579_ sky130_fd_sc_hd__clkbuf_1
X_14915_ net4198 net4197 VGND VGND VPWR VPWR _06989_ sky130_fd_sc_hd__or2_1
X_18683_ net3988 _10524_ _10527_ _10528_ VGND VGND VPWR VPWR _10529_ sky130_fd_sc_hd__o211a_1
X_15895_ net3530 net3481 VGND VGND VPWR VPWR _07964_ sky130_fd_sc_hd__nor2_1
X_17634_ net4004 net6747 net1458 _09493_ _09514_ VGND VGND VPWR VPWR _09515_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14846_ _06940_ VGND VGND VPWR VPWR _00194_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_187_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17565_ net6739 svm0.tC\[0\] VGND VGND VPWR VPWR _09447_ sky130_fd_sc_hd__and2_1
X_14777_ net3616 _06855_ VGND VGND VPWR VPWR _06902_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19304_ net6312 net3888 net6342 VGND VGND VPWR VPWR _11141_ sky130_fd_sc_hd__a21o_1
X_16516_ net2623 net2208 _08575_ VGND VGND VPWR VPWR _08576_ sky130_fd_sc_hd__and3_1
X_13728_ _05919_ _05996_ VGND VGND VPWR VPWR _05997_ sky130_fd_sc_hd__and2b_1
XFILLER_0_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17496_ net3275 _09384_ net6660 VGND VGND VPWR VPWR _09385_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_156_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19235_ net6336 net6225 VGND VGND VPWR VPWR _11072_ sky130_fd_sc_hd__or2b_1
XFILLER_0_73_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16447_ net2621 net2639 _08389_ VGND VGND VPWR VPWR _08508_ sky130_fd_sc_hd__or3_1
X_13659_ _05806_ _05833_ _05928_ VGND VGND VPWR VPWR _05929_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_112_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_140_Right_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19166_ net3189 _10945_ VGND VGND VPWR VPWR _11003_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16378_ _08438_ _08439_ net1252 VGND VGND VPWR VPWR _08440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18117_ _09961_ _09964_ _09967_ VGND VGND VPWR VPWR _09968_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15329_ _07366_ _07367_ _07402_ VGND VGND VPWR VPWR _07403_ sky130_fd_sc_hd__o21ai_1
X_19097_ _10925_ _10926_ net1756 _10910_ _10933_ VGND VGND VPWR VPWR _10934_ sky130_fd_sc_hd__a41oi_2
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18048_ _09884_ _09897_ _09898_ VGND VGND VPWR VPWR _09899_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5991 net5997 VGND VGND VPWR VPWR net5991 sky130_fd_sc_hd__clkbuf_1
X_20010_ net350 _11839_ net3126 VGND VGND VPWR VPWR _11840_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19999_ net351 _11782_ VGND VGND VPWR VPWR _11830_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21961_ _01959_ _01968_ VGND VGND VPWR VPWR _01969_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_179_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23700_ pid_q.curr_error\[2\] VGND VGND VPWR VPWR _03567_ sky130_fd_sc_hd__inv_2
X_20912_ _00810_ _00816_ VGND VGND VPWR VPWR _00928_ sky130_fd_sc_hd__xnor2_1
X_24680_ net9184 net1647 _04522_ VGND VGND VPWR VPWR _00692_ sky130_fd_sc_hd__a21o_1
X_21892_ _01896_ _01900_ _01744_ VGND VGND VPWR VPWR _01901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23631_ net4728 net4822 VGND VGND VPWR VPWR _03498_ sky130_fd_sc_hd__nand2_1
X_20843_ net1735 net1393 VGND VGND VPWR VPWR _00859_ sky130_fd_sc_hd__xor2_1
XFILLER_0_7_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23562_ _03426_ _03429_ VGND VGND VPWR VPWR _03430_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_159_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20774_ _12543_ _12544_ VGND VGND VPWR VPWR _12545_ sky130_fd_sc_hd__xnor2_1
Xmax_length4804 net4805 VGND VGND VPWR VPWR net4804 sky130_fd_sc_hd__buf_1
XFILLER_0_71_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25301_ clknet_leaf_70_clk _00184_ net8447 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.e\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22513_ _02455_ net517 VGND VGND VPWR VPWR _02514_ sky130_fd_sc_hd__and2_1
XFILLER_0_190_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23493_ net2420 _03361_ VGND VGND VPWR VPWR _03362_ sky130_fd_sc_hd__xnor2_1
Xmax_length4848 net4841 VGND VGND VPWR VPWR net4848 sky130_fd_sc_hd__buf_1
Xwire807 _01215_ VGND VGND VPWR VPWR net807 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_174_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire818 _09996_ VGND VGND VPWR VPWR net818 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22444_ net5377 _02445_ VGND VGND VPWR VPWR _02446_ sky130_fd_sc_hd__nand2_1
X_25232_ clknet_leaf_65_clk _00121_ net8655 VGND VGND VPWR VPWR pid_d.iterate_enable
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire829 _07330_ VGND VGND VPWR VPWR net829 sky130_fd_sc_hd__buf_1
XFILLER_0_73_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22375_ _02371_ _02376_ VGND VGND VPWR VPWR _02378_ sky130_fd_sc_hd__or2_1
X_25163_ clknet_leaf_54_clk _00052_ net8730 VGND VGND VPWR VPWR svm0.periodTop\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24114_ net2025 _03975_ VGND VGND VPWR VPWR _03976_ sky130_fd_sc_hd__xnor2_2
X_21326_ net5983 pid_d.prev_int\[2\] VGND VGND VPWR VPWR _01340_ sky130_fd_sc_hd__xnor2_1
X_25094_ net4401 net5172 _04824_ net5174 VGND VGND VPWR VPWR _04838_ sky130_fd_sc_hd__a211o_1
Xwire4103 net4104 VGND VGND VPWR VPWR net4103 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4125 _07037_ VGND VGND VPWR VPWR net4125 sky130_fd_sc_hd__buf_1
Xwire4136 net4137 VGND VGND VPWR VPWR net4136 sky130_fd_sc_hd__buf_1
X_24045_ _03906_ _03907_ VGND VGND VPWR VPWR _03908_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4147 _07020_ VGND VGND VPWR VPWR net4147 sky130_fd_sc_hd__clkbuf_1
Xwire3402 net3403 VGND VGND VPWR VPWR net3402 sky130_fd_sc_hd__dlymetal6s2s_1
X_21257_ _00844_ _00848_ _01271_ VGND VGND VPWR VPWR _01272_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4158 net4159 VGND VGND VPWR VPWR net4158 sky130_fd_sc_hd__buf_1
Xwire3413 net3414 VGND VGND VPWR VPWR net3413 sky130_fd_sc_hd__buf_1
Xwire3424 _07486_ VGND VGND VPWR VPWR net3424 sky130_fd_sc_hd__buf_1
Xwire4169 net4170 VGND VGND VPWR VPWR net4169 sky130_fd_sc_hd__buf_1
X_20208_ _12029_ net3126 net179 VGND VGND VPWR VPWR _12032_ sky130_fd_sc_hd__mux2_1
Xwire3435 net3436 VGND VGND VPWR VPWR net3435 sky130_fd_sc_hd__buf_1
Xwire2701 net2702 VGND VGND VPWR VPWR net2701 sky130_fd_sc_hd__buf_1
Xwire3446 _07245_ VGND VGND VPWR VPWR net3446 sky130_fd_sc_hd__buf_1
X_21188_ _01157_ _01161_ _01203_ VGND VGND VPWR VPWR _01204_ sky130_fd_sc_hd__o21a_1
Xwire3457 _07192_ VGND VGND VPWR VPWR net3457 sky130_fd_sc_hd__clkbuf_1
Xwire2723 net2724 VGND VGND VPWR VPWR net2723 sky130_fd_sc_hd__buf_1
Xwire3468 net3469 VGND VGND VPWR VPWR net3468 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2734 net2735 VGND VGND VPWR VPWR net2734 sky130_fd_sc_hd__buf_1
Xwire3479 net3480 VGND VGND VPWR VPWR net3479 sky130_fd_sc_hd__clkbuf_1
X_20139_ net8972 net2124 net1445 _11966_ VGND VGND VPWR VPWR _00462_ sky130_fd_sc_hd__a31o_1
Xwire2745 net2746 VGND VGND VPWR VPWR net2745 sky130_fd_sc_hd__clkbuf_1
Xwire2756 net2757 VGND VGND VPWR VPWR net2756 sky130_fd_sc_hd__buf_1
Xwire2767 net2768 VGND VGND VPWR VPWR net2767 sky130_fd_sc_hd__clkbuf_1
Xwire2778 _07142_ VGND VGND VPWR VPWR net2778 sky130_fd_sc_hd__buf_1
X_24947_ _04725_ VGND VGND VPWR VPWR _00756_ sky130_fd_sc_hd__clkbuf_1
X_12961_ _05224_ net1003 _05214_ net1593 _05233_ VGND VGND VPWR VPWR _05234_ sky130_fd_sc_hd__a41o_1
XFILLER_0_35_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14700_ net7152 _06842_ net7459 VGND VGND VPWR VPWR _06845_ sky130_fd_sc_hd__o21ai_1
X_15680_ net2674 _07687_ _07750_ net2728 VGND VGND VPWR VPWR _07751_ sky130_fd_sc_hd__a2bb2o_1
X_24878_ _04676_ net4630 net1996 VGND VGND VPWR VPWR _04677_ sky130_fd_sc_hd__mux2_1
X_12892_ _05162_ _05163_ _05160_ _05161_ VGND VGND VPWR VPWR _05165_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_169_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14631_ net7551 net7461 _04877_ VGND VGND VPWR VPWR _06798_ sky130_fd_sc_hd__mux2_1
X_23829_ net5066 net4483 VGND VGND VPWR VPWR _03694_ sky130_fd_sc_hd__nand2_2
XFILLER_0_135_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17350_ net7630 _09214_ _09205_ VGND VGND VPWR VPWR _09264_ sky130_fd_sc_hd__o21a_1
X_14562_ net7257 net5223 VGND VGND VPWR VPWR _06739_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16301_ _08361_ _08364_ VGND VGND VPWR VPWR _08365_ sky130_fd_sc_hd__or2_1
X_13513_ _05694_ net728 _05693_ VGND VGND VPWR VPWR _05784_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17281_ net6741 VGND VGND VPWR VPWR _09196_ sky130_fd_sc_hd__inv_2
X_14493_ _06673_ _06676_ VGND VGND VPWR VPWR _06677_ sky130_fd_sc_hd__xnor2_1
X_19020_ net6248 _10856_ VGND VGND VPWR VPWR _10857_ sky130_fd_sc_hd__xnor2_1
X_16232_ _08247_ _08296_ VGND VGND VPWR VPWR _08297_ sky130_fd_sc_hd__xnor2_4
X_13444_ _05596_ _05597_ _05599_ _05600_ VGND VGND VPWR VPWR _05717_ sky130_fd_sc_hd__and4_1
XFILLER_0_152_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16163_ _08147_ _08227_ _08228_ VGND VGND VPWR VPWR _08229_ sky130_fd_sc_hd__o21ai_2
X_13375_ _05645_ _05646_ _05647_ VGND VGND VPWR VPWR _05648_ sky130_fd_sc_hd__and3_1
Xfanout5243 matmul0.beta_pass\[8\] VGND VGND VPWR VPWR net5243 sky130_fd_sc_hd__buf_1
Xwire6050 net6047 VGND VGND VPWR VPWR net6050 sky130_fd_sc_hd__buf_1
Xwire6061 net6062 VGND VGND VPWR VPWR net6061 sky130_fd_sc_hd__buf_1
X_15114_ _07186_ _07187_ VGND VGND VPWR VPWR _07188_ sky130_fd_sc_hd__xnor2_1
Xwire6072 net6068 VGND VGND VPWR VPWR net6072 sky130_fd_sc_hd__buf_1
XFILLER_0_11_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16094_ net385 net493 VGND VGND VPWR VPWR _08161_ sky130_fd_sc_hd__xnor2_1
Xwire6094 net6095 VGND VGND VPWR VPWR net6094 sky130_fd_sc_hd__buf_1
XFILLER_0_142_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19922_ net6072 _10996_ VGND VGND VPWR VPWR _11754_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15045_ net2850 _07118_ _07116_ _07117_ VGND VGND VPWR VPWR _07119_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5393 net5394 VGND VGND VPWR VPWR net5393 sky130_fd_sc_hd__buf_1
XFILLER_0_76_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4670 net4671 VGND VGND VPWR VPWR net4670 sky130_fd_sc_hd__clkbuf_1
Xwire4681 net4682 VGND VGND VPWR VPWR net4681 sky130_fd_sc_hd__buf_1
X_19853_ net6049 net3856 VGND VGND VPWR VPWR _11686_ sky130_fd_sc_hd__xnor2_4
X_18804_ _10589_ _10647_ VGND VGND VPWR VPWR _10648_ sky130_fd_sc_hd__xor2_1
Xwire3980 net3984 VGND VGND VPWR VPWR net3980 sky130_fd_sc_hd__clkbuf_1
X_16996_ _08952_ net1806 VGND VGND VPWR VPWR _08958_ sky130_fd_sc_hd__nand2_1
X_19784_ _11616_ _11617_ VGND VGND VPWR VPWR _11618_ sky130_fd_sc_hd__nand2_1
XFILLER_0_183_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15947_ net1527 net1262 _07988_ VGND VGND VPWR VPWR _08015_ sky130_fd_sc_hd__a21bo_1
X_18735_ net6955 net6878 VGND VGND VPWR VPWR _10580_ sky130_fd_sc_hd__or2_1
XFILLER_0_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18666_ net9075 net2287 net1450 _10512_ VGND VGND VPWR VPWR _00443_ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15878_ net1845 net1842 VGND VGND VPWR VPWR _07947_ sky130_fd_sc_hd__and2_1
XFILLER_0_188_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17617_ net6739 svm0.tB\[0\] VGND VGND VPWR VPWR _09498_ sky130_fd_sc_hd__or2_1
X_14829_ _06931_ VGND VGND VPWR VPWR _00186_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18597_ net6860 net3285 net2129 VGND VGND VPWR VPWR _10445_ sky130_fd_sc_hd__a21o_1
XFILLER_0_188_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17548_ net6722 svm0.tC\[6\] VGND VGND VPWR VPWR _09430_ sky130_fd_sc_hd__and2b_1
XFILLER_0_86_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17479_ net6718 _09369_ _09370_ _09368_ VGND VGND VPWR VPWR _00397_ sky130_fd_sc_hd__a22o_1
XFILLER_0_184_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19218_ net6340 net3882 _11051_ net3874 _10846_ VGND VGND VPWR VPWR _11055_ sky130_fd_sc_hd__o221a_1
XFILLER_0_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20490_ net3848 _12275_ net3847 _12277_ net3334 net3333 VGND VGND VPWR VPWR _12278_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_26_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19149_ net3895 _10985_ VGND VGND VPWR VPWR _10986_ sky130_fd_sc_hd__nor2_2
XFILLER_0_15_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22160_ net859 _02165_ VGND VGND VPWR VPWR _02166_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_124_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21111_ net5630 net5870 VGND VGND VPWR VPWR _01127_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22091_ _02096_ _02097_ VGND VGND VPWR VPWR _02098_ sky130_fd_sc_hd__nor2_1
X_21042_ _01001_ _01057_ VGND VGND VPWR VPWR _01058_ sky130_fd_sc_hd__xnor2_2
Xwire2008 _04641_ VGND VGND VPWR VPWR net2008 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2019 _04217_ VGND VGND VPWR VPWR net2019 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1307 _05873_ VGND VGND VPWR VPWR net1307 sky130_fd_sc_hd__dlymetal6s2s_1
X_25850_ clknet_leaf_20_clk _00723_ net8745 VGND VGND VPWR VPWR pid_q.mult0.b\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1318 net1319 VGND VGND VPWR VPWR net1318 sky130_fd_sc_hd__buf_1
Xwire1329 _05556_ VGND VGND VPWR VPWR net1329 sky130_fd_sc_hd__clkbuf_1
X_24801_ net8983 net1644 _04542_ _04625_ VGND VGND VPWR VPWR _00710_ sky130_fd_sc_hd__a22o_1
X_25781_ clknet_leaf_58_clk _00654_ net8713 VGND VGND VPWR VPWR matmul0.beta_pass\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_22993_ _02864_ VGND VGND VPWR VPWR _00663_ sky130_fd_sc_hd__clkbuf_1
X_24732_ _04563_ _04564_ net4232 VGND VGND VPWR VPWR _04565_ sky130_fd_sc_hd__a21o_1
X_21944_ _01946_ _01951_ VGND VGND VPWR VPWR _01952_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_179_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24663_ pid_q.curr_error\[3\] net2382 net1372 VGND VGND VPWR VPWR _04514_ sky130_fd_sc_hd__and3_1
X_21875_ _01879_ _01882_ _01883_ VGND VGND VPWR VPWR _01884_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_16_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout8808 net8834 VGND VGND VPWR VPWR net8808 sky130_fd_sc_hd__buf_1
X_23614_ net8996 net3062 net2028 _03481_ VGND VGND VPWR VPWR _00667_ sky130_fd_sc_hd__a22o_1
X_20826_ net5761 net5577 VGND VGND VPWR VPWR _00842_ sky130_fd_sc_hd__nand2_1
X_24594_ pid_q.prev_error\[13\] net5166 VGND VGND VPWR VPWR _04450_ sky130_fd_sc_hd__nand2_1
Xwire8903 net8899 VGND VGND VPWR VPWR net8903 sky130_fd_sc_hd__buf_1
XFILLER_0_119_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8914 net8916 VGND VGND VPWR VPWR net8914 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length4612 net4613 VGND VGND VPWR VPWR net4612 sky130_fd_sc_hd__clkbuf_1
X_23545_ net4575 net5024 VGND VGND VPWR VPWR _03413_ sky130_fd_sc_hd__nand2_1
XFILLER_0_181_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8925 net8926 VGND VGND VPWR VPWR net8925 sky130_fd_sc_hd__clkbuf_1
Xmax_length5357 pid_d.out\[8\] VGND VGND VPWR VPWR net5357 sky130_fd_sc_hd__buf_1
Xwire8936 net8937 VGND VGND VPWR VPWR net8936 sky130_fd_sc_hd__clkbuf_1
X_20757_ net5954 net5454 VGND VGND VPWR VPWR _12528_ sky130_fd_sc_hd__nand2_1
Xwire8947 net8948 VGND VGND VPWR VPWR net8947 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4645 pid_q.mult0.a\[7\] VGND VGND VPWR VPWR net4645 sky130_fd_sc_hd__clkbuf_1
Xmax_length3900 net3901 VGND VGND VPWR VPWR net3900 sky130_fd_sc_hd__clkbuf_1
Xwire604 _11548_ VGND VGND VPWR VPWR net604 sky130_fd_sc_hd__buf_2
Xwire615 net616 VGND VGND VPWR VPWR net615 sky130_fd_sc_hd__buf_1
XFILLER_0_80_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23476_ _03272_ _03273_ _03344_ VGND VGND VPWR VPWR _03345_ sky130_fd_sc_hd__a21oi_2
Xwire626 net627 VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__clkbuf_1
X_20688_ net6762 _12295_ _09096_ VGND VGND VPWR VPWR _12463_ sky130_fd_sc_hd__mux2_2
XFILLER_0_52_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire637 net638 VGND VGND VPWR VPWR net637 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire648 net649 VGND VGND VPWR VPWR net648 sky130_fd_sc_hd__clkbuf_1
X_25215_ clknet_leaf_61_clk _00104_ net8688 VGND VGND VPWR VPWR svm0.vC\[3\] sky130_fd_sc_hd__dfrtp_1
Xmax_length3955 _09798_ VGND VGND VPWR VPWR net3955 sky130_fd_sc_hd__buf_1
XFILLER_0_190_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22427_ _02419_ _02428_ VGND VGND VPWR VPWR _02429_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_134_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire659 net660 VGND VGND VPWR VPWR net659 sky130_fd_sc_hd__buf_1
XFILLER_0_122_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length268 net269 VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25146_ clknet_leaf_41_clk _00035_ net8767 VGND VGND VPWR VPWR pid_q.target\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13160_ _05372_ net1138 _05370_ VGND VGND VPWR VPWR _05433_ sky130_fd_sc_hd__a21oi_1
X_22358_ _02284_ _02286_ _02285_ VGND VGND VPWR VPWR _02361_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13091_ _05361_ _05362_ _05363_ VGND VGND VPWR VPWR _05364_ sky130_fd_sc_hd__nand3_1
X_21309_ _01321_ _01323_ VGND VGND VPWR VPWR _01324_ sky130_fd_sc_hd__xor2_1
X_22289_ net5691 net5435 VGND VGND VPWR VPWR _02293_ sky130_fd_sc_hd__nand2_1
X_25077_ _04822_ _04817_ net4418 VGND VGND VPWR VPWR _04823_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_130_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3210 _10829_ VGND VGND VPWR VPWR net3210 sky130_fd_sc_hd__buf_1
XFILLER_0_130_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3221 net3222 VGND VGND VPWR VPWR net3221 sky130_fd_sc_hd__buf_1
X_24028_ _03817_ _03822_ _03806_ VGND VGND VPWR VPWR _03891_ sky130_fd_sc_hd__a21o_1
Xwire3243 net3244 VGND VGND VPWR VPWR net3243 sky130_fd_sc_hd__clkbuf_1
Xhold290 pid_d.curr_int\[6\] VGND VGND VPWR VPWR net9243 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3254 _09649_ VGND VGND VPWR VPWR net3254 sky130_fd_sc_hd__buf_1
Xwire2520 _10992_ VGND VGND VPWR VPWR net2520 sky130_fd_sc_hd__buf_1
Xwire3265 net3266 VGND VGND VPWR VPWR net3265 sky130_fd_sc_hd__clkbuf_2
Xwire3276 net3277 VGND VGND VPWR VPWR net3276 sky130_fd_sc_hd__buf_1
Xwire2531 net2532 VGND VGND VPWR VPWR net2531 sky130_fd_sc_hd__clkbuf_2
X_16850_ cordic0.sin\[13\] matmul0.sin\[13\] net4287 VGND VGND VPWR VPWR _08816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2542 _10228_ VGND VGND VPWR VPWR net2542 sky130_fd_sc_hd__clkbuf_1
Xwire3287 net3288 VGND VGND VPWR VPWR net3287 sky130_fd_sc_hd__buf_1
Xwire2553 _09743_ VGND VGND VPWR VPWR net2553 sky130_fd_sc_hd__buf_1
Xwire3298 net3299 VGND VGND VPWR VPWR net3298 sky130_fd_sc_hd__buf_1
Xwire2564 _09601_ VGND VGND VPWR VPWR net2564 sky130_fd_sc_hd__buf_1
X_15801_ _07778_ _07779_ _07870_ VGND VGND VPWR VPWR _07871_ sky130_fd_sc_hd__o21a_1
Xwire2575 _09278_ VGND VGND VPWR VPWR net2575 sky130_fd_sc_hd__buf_1
Xwire1830 net1831 VGND VGND VPWR VPWR net1830 sky130_fd_sc_hd__clkbuf_1
Xwire1841 _08253_ VGND VGND VPWR VPWR net1841 sky130_fd_sc_hd__clkbuf_1
X_16781_ net7595 matmul0.a\[10\] net3379 VGND VGND VPWR VPWR _08780_ sky130_fd_sc_hd__mux2_1
X_13993_ _06248_ _06257_ VGND VGND VPWR VPWR _06258_ sky130_fd_sc_hd__xnor2_1
Xwire2597 net2598 VGND VGND VPWR VPWR net2597 sky130_fd_sc_hd__buf_1
Xwire1852 _07653_ VGND VGND VPWR VPWR net1852 sky130_fd_sc_hd__buf_1
XFILLER_0_189_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1863 _07533_ VGND VGND VPWR VPWR net1863 sky130_fd_sc_hd__clkbuf_1
Xwire1874 _07376_ VGND VGND VPWR VPWR net1874 sky130_fd_sc_hd__clkbuf_1
X_18520_ net6817 net3929 VGND VGND VPWR VPWR _10369_ sky130_fd_sc_hd__nor2_1
X_15732_ net1269 net1268 net1108 VGND VGND VPWR VPWR _07803_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_88_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12944_ net2338 net1968 VGND VGND VPWR VPWR _05217_ sky130_fd_sc_hd__and2_1
Xwire1885 _07225_ VGND VGND VPWR VPWR net1885 sky130_fd_sc_hd__clkbuf_1
Xwire1896 net1897 VGND VGND VPWR VPWR net1896 sky130_fd_sc_hd__buf_1
XFILLER_0_153_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18451_ net3941 _10300_ net6970 VGND VGND VPWR VPWR _10301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15663_ net778 _07734_ VGND VGND VPWR VPWR _07735_ sky130_fd_sc_hd__xor2_1
X_12875_ _05083_ _05032_ VGND VGND VPWR VPWR _05148_ sky130_fd_sc_hd__nand2_1
X_17402_ svm0.delta\[9\] VGND VGND VPWR VPWR _09307_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14614_ net6453 _06784_ _06785_ VGND VGND VPWR VPWR _06786_ sky130_fd_sc_hd__and3_1
X_18382_ net7045 net7111 VGND VGND VPWR VPWR _10233_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15594_ net1269 net1268 VGND VGND VPWR VPWR _07666_ sky130_fd_sc_hd__xor2_1
XFILLER_0_29_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6570 net6571 VGND VGND VPWR VPWR net6570 sky130_fd_sc_hd__buf_1
X_17333_ net4017 _09207_ _09244_ _09245_ VGND VGND VPWR VPWR _09247_ sky130_fd_sc_hd__and4_1
XFILLER_0_7_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14545_ net1624 _06722_ _06723_ _06712_ VGND VGND VPWR VPWR _06724_ sky130_fd_sc_hd__a31o_1
XFILLER_0_172_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6592 net6594 VGND VGND VPWR VPWR net6592 sky130_fd_sc_hd__buf_1
XFILLER_0_83_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17264_ net2160 net323 net1798 net9089 VGND VGND VPWR VPWR _00358_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14476_ net9070 net831 net1292 _06662_ VGND VGND VPWR VPWR _00102_ sky130_fd_sc_hd__a22o_1
X_19003_ net3209 _10839_ VGND VGND VPWR VPWR _10840_ sky130_fd_sc_hd__nand2_1
X_16215_ net2691 net2659 VGND VGND VPWR VPWR _08280_ sky130_fd_sc_hd__nor2_1
X_13427_ net7815 net1586 VGND VGND VPWR VPWR _05700_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17195_ net3343 _09096_ _09144_ net5988 VGND VGND VPWR VPWR _09145_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16146_ _08131_ _08136_ _08211_ VGND VGND VPWR VPWR _08212_ sky130_fd_sc_hd__a21oi_1
X_13358_ net1330 _05536_ _05630_ VGND VGND VPWR VPWR _05631_ sky130_fd_sc_hd__o21a_1
Xfanout4361 net4368 VGND VGND VPWR VPWR net4361 sky130_fd_sc_hd__clkbuf_1
X_16077_ _08026_ _08028_ net2846 net2224 VGND VGND VPWR VPWR _08144_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_80_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13289_ _05558_ _05561_ VGND VGND VPWR VPWR _05562_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout4383 net4386 VGND VGND VPWR VPWR net4383 sky130_fd_sc_hd__buf_1
Xwire5190 net5191 VGND VGND VPWR VPWR net5190 sky130_fd_sc_hd__buf_1
X_19905_ _11712_ _11714_ VGND VGND VPWR VPWR _11737_ sky130_fd_sc_hd__and2_1
X_15028_ _07097_ _07098_ net2809 _07101_ VGND VGND VPWR VPWR _07102_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19836_ _11667_ net708 VGND VGND VPWR VPWR _11670_ sky130_fd_sc_hd__xnor2_1
X_19767_ net2504 VGND VGND VPWR VPWR _11602_ sky130_fd_sc_hd__inv_2
Xinput3 angle_in[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
X_16979_ net3349 _08941_ VGND VGND VPWR VPWR _08942_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18718_ _10561_ net764 VGND VGND VPWR VPWR _10564_ sky130_fd_sc_hd__or2_1
X_19698_ _11443_ _11470_ _11533_ VGND VGND VPWR VPWR _11534_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_78_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18649_ net2589 net2129 _10445_ net6831 VGND VGND VPWR VPWR _10496_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21660_ _01665_ _01670_ VGND VGND VPWR VPWR _01671_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20611_ net6217 _12369_ VGND VGND VPWR VPWR _12392_ sky130_fd_sc_hd__xnor2_1
X_21591_ net1178 _01602_ VGND VGND VPWR VPWR _01603_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7509 net7507 VGND VGND VPWR VPWR net7509 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23330_ net1675 _03199_ VGND VGND VPWR VPWR _03200_ sky130_fd_sc_hd__xnor2_2
X_20542_ net6326 _12326_ VGND VGND VPWR VPWR _12327_ sky130_fd_sc_hd__or2b_1
XFILLER_0_105_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length2506 _11446_ VGND VGND VPWR VPWR net2506 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_15_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23261_ _03121_ _03122_ VGND VGND VPWR VPWR _03131_ sky130_fd_sc_hd__nand2_1
X_20473_ net2178 _12258_ net3353 VGND VGND VPWR VPWR _12263_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25000_ net4474 net5183 _04756_ VGND VGND VPWR VPWR _04757_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22212_ net5707 net5430 VGND VGND VPWR VPWR _02217_ sky130_fd_sc_hd__nand2_1
X_23192_ _03053_ _03056_ _03061_ VGND VGND VPWR VPWR _03062_ sky130_fd_sc_hd__a21oi_1
X_22143_ _02038_ _02049_ _02148_ VGND VGND VPWR VPWR _02149_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22074_ _02070_ _02080_ VGND VGND VPWR VPWR _02081_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_168_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25902_ clknet_leaf_17_clk _00775_ net8632 VGND VGND VPWR VPWR pid_q.kp\[14\] sky130_fd_sc_hd__dfrtp_1
X_21025_ _01037_ _01038_ _01040_ VGND VGND VPWR VPWR _01041_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_96_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1104 net1105 VGND VGND VPWR VPWR net1104 sky130_fd_sc_hd__buf_1
Xwire1115 _07523_ VGND VGND VPWR VPWR net1115 sky130_fd_sc_hd__clkbuf_1
Xwire1126 net1127 VGND VGND VPWR VPWR net1126 sky130_fd_sc_hd__clkbuf_2
X_25833_ clknet_leaf_37_clk _00706_ net8746 VGND VGND VPWR VPWR pid_q.curr_error\[9\]
+ sky130_fd_sc_hd__dfrtp_2
Xwire1137 _05438_ VGND VGND VPWR VPWR net1137 sky130_fd_sc_hd__buf_1
Xwire1148 net1149 VGND VGND VPWR VPWR net1148 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1159 _04077_ VGND VGND VPWR VPWR net1159 sky130_fd_sc_hd__buf_1
XFILLER_0_57_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25764_ clknet_leaf_67_clk _00637_ net8456 VGND VGND VPWR VPWR pid_d.out\[5\] sky130_fd_sc_hd__dfrtp_1
X_22976_ matmul0.beta_pass\[7\] net823 net6569 VGND VGND VPWR VPWR _02856_ sky130_fd_sc_hd__mux2_1
X_24715_ net8022 _04546_ net5290 VGND VGND VPWR VPWR _04550_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21927_ net5750 net5463 VGND VGND VPWR VPWR _01935_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25695_ clknet_leaf_0_clk _00568_ net8406 VGND VGND VPWR VPWR pid_d.mult0.b\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout8605 net8821 VGND VGND VPWR VPWR net8605 sky130_fd_sc_hd__clkbuf_2
X_24646_ net509 _04500_ VGND VGND VPWR VPWR _04501_ sky130_fd_sc_hd__xor2_1
X_12660_ net7760 net2340 _04932_ VGND VGND VPWR VPWR _04933_ sky130_fd_sc_hd__and3_1
XFILLER_0_171_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21858_ _01866_ net5857 _01783_ VGND VGND VPWR VPWR _01867_ sky130_fd_sc_hd__a21bo_1
Xfanout8627 net8629 VGND VGND VPWR VPWR net8627 sky130_fd_sc_hd__buf_1
XFILLER_0_139_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8700 net8696 VGND VGND VPWR VPWR net8700 sky130_fd_sc_hd__buf_1
XFILLER_0_136_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout8649 net8653 VGND VGND VPWR VPWR net8649 sky130_fd_sc_hd__buf_1
XFILLER_0_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20809_ _12504_ _12505_ _00824_ VGND VGND VPWR VPWR _00825_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_154_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24577_ _04290_ net4506 _04431_ _04432_ net4491 VGND VGND VPWR VPWR _04433_ sky130_fd_sc_hd__o311a_1
X_12591_ net3709 VGND VGND VPWR VPWR _04874_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_116_clk clknet_4_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_116_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_167_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21789_ _01796_ net2063 VGND VGND VPWR VPWR _01799_ sky130_fd_sc_hd__xnor2_2
Xwire8733 net8734 VGND VGND VPWR VPWR net8733 sky130_fd_sc_hd__buf_1
Xwire8744 net8745 VGND VGND VPWR VPWR net8744 sky130_fd_sc_hd__buf_1
X_14330_ _06549_ matmul0.a_in\[2\] net902 VGND VGND VPWR VPWR _06550_ sky130_fd_sc_hd__mux2_1
X_23528_ _03394_ _03395_ VGND VGND VPWR VPWR _03396_ sky130_fd_sc_hd__xnor2_1
Xwire8755 net8751 VGND VGND VPWR VPWR net8755 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire401 net402 VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire412 net413 VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__clkbuf_1
Xwire8777 net8773 VGND VGND VPWR VPWR net8777 sky130_fd_sc_hd__clkbuf_2
Xmax_length3730 _04531_ VGND VGND VPWR VPWR net3730 sky130_fd_sc_hd__buf_1
Xwire423 _08726_ VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__buf_1
XFILLER_0_53_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8788 net8789 VGND VGND VPWR VPWR net8788 sky130_fd_sc_hd__buf_1
Xwire434 net435 VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__clkbuf_1
X_14261_ net2923 VGND VGND VPWR VPWR _06515_ sky130_fd_sc_hd__buf_1
Xmax_length4486 net4482 VGND VGND VPWR VPWR net4486 sky130_fd_sc_hd__buf_1
XFILLER_0_18_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire445 net446 VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__clkbuf_1
X_23459_ _03265_ _03266_ _03327_ VGND VGND VPWR VPWR _03328_ sky130_fd_sc_hd__a21bo_1
Xwire456 _04611_ VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire467 net468 VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__buf_1
XFILLER_0_135_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16000_ _07979_ net1094 _08067_ VGND VGND VPWR VPWR _08068_ sky130_fd_sc_hd__a21o_1
X_13212_ _05483_ _05484_ net682 VGND VGND VPWR VPWR _05485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire478 _01532_ VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__buf_1
XFILLER_0_151_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire489 _10341_ VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__clkbuf_1
X_14192_ _06451_ _06416_ _06415_ VGND VGND VPWR VPWR _06452_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_20_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25129_ clknet_leaf_52_clk _00018_ net8805 VGND VGND VPWR VPWR svm0.tC\[1\] sky130_fd_sc_hd__dfrtp_1
X_13143_ _05412_ _05415_ VGND VGND VPWR VPWR _05416_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13074_ net6664 net6673 net6677 svm0.vC\[12\] VGND VGND VPWR VPWR _05347_ sky130_fd_sc_hd__nand4b_1
X_17951_ _09800_ net3993 net4044 VGND VGND VPWR VPWR _09802_ sky130_fd_sc_hd__o21ai_1
Xwire3040 net3041 VGND VGND VPWR VPWR net3040 sky130_fd_sc_hd__clkbuf_2
Xwire3051 _03373_ VGND VGND VPWR VPWR net3051 sky130_fd_sc_hd__clkbuf_1
Xwire3062 net3063 VGND VGND VPWR VPWR net3062 sky130_fd_sc_hd__buf_1
X_16902_ cordic0.slte0.opA\[8\] net6407 VGND VGND VPWR VPWR _08866_ sky130_fd_sc_hd__or2b_1
X_17882_ _09728_ _09732_ VGND VGND VPWR VPWR _09733_ sky130_fd_sc_hd__xnor2_1
Xwire3073 net3074 VGND VGND VPWR VPWR net3073 sky130_fd_sc_hd__clkbuf_1
Xwire3095 net3096 VGND VGND VPWR VPWR net3095 sky130_fd_sc_hd__buf_1
Xwire2361 net2362 VGND VGND VPWR VPWR net2361 sky130_fd_sc_hd__buf_1
X_19621_ _11450_ _11457_ VGND VGND VPWR VPWR _11458_ sky130_fd_sc_hd__xnor2_2
Xwire2372 net2373 VGND VGND VPWR VPWR net2372 sky130_fd_sc_hd__clkbuf_1
X_16833_ _08807_ VGND VGND VPWR VPWR _00314_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2394 net2395 VGND VGND VPWR VPWR net2394 sky130_fd_sc_hd__buf_1
XFILLER_0_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1660 _03693_ VGND VGND VPWR VPWR net1660 sky130_fd_sc_hd__buf_1
Xwire1671 net1672 VGND VGND VPWR VPWR net1671 sky130_fd_sc_hd__clkbuf_1
X_19552_ _11387_ _11388_ VGND VGND VPWR VPWR _11389_ sky130_fd_sc_hd__nand2_1
X_16764_ _08771_ VGND VGND VPWR VPWR _00281_ sky130_fd_sc_hd__clkbuf_1
X_13976_ _06191_ _06196_ _06189_ VGND VGND VPWR VPWR _06241_ sky130_fd_sc_hd__a21bo_1
Xwire1682 net1683 VGND VGND VPWR VPWR net1682 sky130_fd_sc_hd__clkbuf_1
Xwire1693 net1694 VGND VGND VPWR VPWR net1693 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_189_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15715_ net3585 net3578 net4087 net4086 VGND VGND VPWR VPWR _07786_ sky130_fd_sc_hd__o22a_1
X_18503_ _10347_ _10348_ _10351_ _10289_ VGND VGND VPWR VPWR _10352_ sky130_fd_sc_hd__a211o_1
X_12927_ _05119_ _05120_ net1006 net1005 VGND VGND VPWR VPWR _05200_ sky130_fd_sc_hd__a211o_1
X_19483_ net3196 _11264_ _10851_ VGND VGND VPWR VPWR _11320_ sky130_fd_sc_hd__mux2_1
X_16695_ matmul0.matmul_stage_inst.mult2\[11\] matmul0.matmul_stage_inst.mult1\[11\]
+ VGND VGND VPWR VPWR _08725_ sky130_fd_sc_hd__xor2_1
XFILLER_0_38_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15646_ net2661 _07717_ VGND VGND VPWR VPWR _07718_ sky130_fd_sc_hd__xnor2_1
X_18434_ net6836 net6859 _10282_ _10283_ VGND VGND VPWR VPWR _10284_ sky130_fd_sc_hd__o211a_1
X_12858_ net2305 VGND VGND VPWR VPWR _05131_ sky130_fd_sc_hd__clkbuf_1
Xmax_length7090 net7091 VGND VGND VPWR VPWR net7090 sky130_fd_sc_hd__buf_1
XFILLER_0_146_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18365_ net6825 net6798 _10210_ _10215_ VGND VGND VPWR VPWR _10216_ sky130_fd_sc_hd__a31o_1
X_15577_ net2837 net3440 VGND VGND VPWR VPWR _07649_ sky130_fd_sc_hd__nor2_1
X_12789_ net7932 net1959 net1960 _05060_ _05061_ VGND VGND VPWR VPWR _05062_ sky130_fd_sc_hd__a311oi_1
X_17316_ net6728 VGND VGND VPWR VPWR _09230_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14528_ net9030 _06652_ net676 net2886 VGND VGND VPWR VPWR _00109_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_1_Left_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18296_ _10025_ _09821_ _09820_ VGND VGND VPWR VPWR _10147_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_126_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17247_ net2165 net224 net1800 net9167 VGND VGND VPWR VPWR _00345_ sky130_fd_sc_hd__a22o_1
X_14459_ net9192 _06646_ _06647_ _06648_ VGND VGND VPWR VPWR _00099_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17178_ net618 _09129_ VGND VGND VPWR VPWR _09130_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire990 _07301_ VGND VGND VPWR VPWR net990 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16129_ net3522 net3424 net3429 net3533 VGND VGND VPWR VPWR _08195_ sky130_fd_sc_hd__a211o_1
XFILLER_0_84_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19819_ net1188 _11652_ VGND VGND VPWR VPWR _11653_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22830_ _02729_ _02730_ VGND VGND VPWR VPWR _02731_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22761_ _02685_ VGND VGND VPWR VPWR _00610_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24500_ _04286_ _04305_ _04356_ VGND VGND VPWR VPWR _04357_ sky130_fd_sc_hd__a21o_1
X_21712_ _01617_ _01625_ VGND VGND VPWR VPWR _01723_ sky130_fd_sc_hd__nand2_1
X_25480_ clknet_leaf_52_clk _00360_ net8787 VGND VGND VPWR VPWR svm0.tA\[2\] sky130_fd_sc_hd__dfrtp_1
X_22692_ _02636_ VGND VGND VPWR VPWR _00590_ sky130_fd_sc_hd__clkbuf_1
X_24431_ net4490 _04287_ _04288_ VGND VGND VPWR VPWR _04289_ sky130_fd_sc_hd__o21a_1
Xwire8007 net8008 VGND VGND VPWR VPWR net8007 sky130_fd_sc_hd__buf_1
X_21643_ net1177 _01601_ _01653_ VGND VGND VPWR VPWR _01654_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8018 net8019 VGND VGND VPWR VPWR net8018 sky130_fd_sc_hd__clkbuf_1
Xwire8029 net8030 VGND VGND VPWR VPWR net8029 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_170_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7306 net7307 VGND VGND VPWR VPWR net7306 sky130_fd_sc_hd__buf_1
X_24362_ _04213_ _04220_ VGND VGND VPWR VPWR _04221_ sky130_fd_sc_hd__xnor2_2
Xwire7317 net7318 VGND VGND VPWR VPWR net7317 sky130_fd_sc_hd__buf_1
X_21574_ net5856 net5418 VGND VGND VPWR VPWR _01586_ sky130_fd_sc_hd__nand2_1
XFILLER_0_191_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire7339 matmul0.alpha_pass\[3\] VGND VGND VPWR VPWR net7339 sky130_fd_sc_hd__clkbuf_1
X_23313_ _02946_ _02961_ _03182_ VGND VGND VPWR VPWR _03183_ sky130_fd_sc_hd__o21ai_1
Xwire6605 net6606 VGND VGND VPWR VPWR net6605 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5809 net5829 VGND VGND VPWR VPWR net5809 sky130_fd_sc_hd__buf_1
X_20525_ net1479 _12310_ VGND VGND VPWR VPWR _12311_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6616 net6617 VGND VGND VPWR VPWR net6616 sky130_fd_sc_hd__buf_1
X_24293_ _04067_ net1379 net1380 VGND VGND VPWR VPWR _04153_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_133_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6627 net6628 VGND VGND VPWR VPWR net6627 sky130_fd_sc_hd__clkbuf_1
Xwire6649 net6650 VGND VGND VPWR VPWR net6649 sky130_fd_sc_hd__buf_1
Xwire5904 net5903 VGND VGND VPWR VPWR net5904 sky130_fd_sc_hd__clkbuf_1
X_23244_ _03092_ _03113_ VGND VGND VPWR VPWR _03114_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_104_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5915 net5916 VGND VGND VPWR VPWR net5915 sky130_fd_sc_hd__clkbuf_1
X_20456_ net9191 _12247_ _12248_ _12246_ VGND VGND VPWR VPWR _00497_ sky130_fd_sc_hd__a22o_1
Xwire5926 net5927 VGND VGND VPWR VPWR net5926 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5937 net5939 VGND VGND VPWR VPWR net5937 sky130_fd_sc_hd__buf_1
XFILLER_0_179_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5959 net5960 VGND VGND VPWR VPWR net5959 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23175_ _03038_ _03043_ _03033_ VGND VGND VPWR VPWR _03045_ sky130_fd_sc_hd__a21o_1
X_20387_ _12184_ _12185_ _12151_ _12155_ VGND VGND VPWR VPWR _12186_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_24_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22126_ _02130_ _02131_ VGND VGND VPWR VPWR _02132_ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22057_ _02060_ _02061_ net1710 VGND VGND VPWR VPWR _02064_ sky130_fd_sc_hd__o21ai_1
X_21008_ _01021_ _01023_ VGND VGND VPWR VPWR _01024_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_173_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13830_ _06036_ _06037_ net7721 net1307 VGND VGND VPWR VPWR _06097_ sky130_fd_sc_hd__o211a_1
X_25816_ clknet_leaf_37_clk _00689_ net8750 VGND VGND VPWR VPWR pid_q.prev_error\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13761_ net3676 _06028_ net2948 net7789 net1940 VGND VGND VPWR VPWR _06029_ sky130_fd_sc_hd__o2111ai_1
X_25747_ clknet_leaf_9_clk _00620_ net8560 VGND VGND VPWR VPWR pid_d.kp\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22959_ _02843_ _02846_ VGND VGND VPWR VPWR _02847_ sky130_fd_sc_hd__xnor2_1
X_15500_ net6540 net6594 matmul0.matmul_stage_inst.e\[14\] VGND VGND VPWR VPWR _07573_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_167_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12712_ net7939 net2368 net2365 VGND VGND VPWR VPWR _04985_ sky130_fd_sc_hd__and3_2
X_16480_ _08501_ _08540_ VGND VGND VPWR VPWR _08541_ sky130_fd_sc_hd__xnor2_1
X_13692_ _05954_ _05960_ VGND VGND VPWR VPWR _05961_ sky130_fd_sc_hd__xnor2_1
X_25678_ clknet_leaf_0_clk _00551_ net8405 VGND VGND VPWR VPWR pid_d.curr_error\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_15431_ net3534 VGND VGND VPWR VPWR _07505_ sky130_fd_sc_hd__buf_1
X_24629_ net4823 _04483_ VGND VGND VPWR VPWR _04484_ sky130_fd_sc_hd__nand2_1
X_12643_ _04903_ _04915_ VGND VGND VPWR VPWR _04916_ sky130_fd_sc_hd__xnor2_2
Xfanout8435 net8438 VGND VGND VPWR VPWR net8435 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout8457 net8459 VGND VGND VPWR VPWR net8457 sky130_fd_sc_hd__clkbuf_2
Xfanout8468 net8475 VGND VGND VPWR VPWR net8468 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_182_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout7734 net7754 VGND VGND VPWR VPWR net7734 sky130_fd_sc_hd__buf_1
X_18150_ _09951_ _09997_ _09999_ _10000_ VGND VGND VPWR VPWR _10001_ sky130_fd_sc_hd__o22a_1
X_15362_ _07418_ _07423_ VGND VGND VPWR VPWR _07436_ sky130_fd_sc_hd__xor2_1
Xwire8541 net8542 VGND VGND VPWR VPWR net8541 sky130_fd_sc_hd__clkbuf_1
Xfanout8479 net8529 VGND VGND VPWR VPWR net8479 sky130_fd_sc_hd__buf_1
Xfanout7745 net7752 VGND VGND VPWR VPWR net7745 sky130_fd_sc_hd__buf_1
X_12574_ net4313 pid_q.state\[0\] _04862_ VGND VGND VPWR VPWR _00016_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8552 net8553 VGND VGND VPWR VPWR net8552 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_92_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4250 _05972_ VGND VGND VPWR VPWR net4250 sky130_fd_sc_hd__buf_1
X_17101_ net1478 _09037_ VGND VGND VPWR VPWR _09058_ sky130_fd_sc_hd__nor2_1
Xwire220 net221 VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__buf_1
X_14313_ net5370 _06523_ _06534_ VGND VGND VPWR VPWR _06535_ sky130_fd_sc_hd__o21a_1
Xwire8574 net8573 VGND VGND VPWR VPWR net8574 sky130_fd_sc_hd__buf_1
XFILLER_0_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7840 net7841 VGND VGND VPWR VPWR net7840 sky130_fd_sc_hd__buf_1
Xwire231 _04453_ VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__buf_1
XFILLER_0_123_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18081_ _09754_ _09885_ VGND VGND VPWR VPWR _09932_ sky130_fd_sc_hd__xnor2_2
Xwire8596 net8597 VGND VGND VPWR VPWR net8596 sky130_fd_sc_hd__clkbuf_1
X_15293_ _07343_ _07344_ _07365_ VGND VGND VPWR VPWR _07367_ sky130_fd_sc_hd__a21oi_1
Xwire7862 net7863 VGND VGND VPWR VPWR net7862 sky130_fd_sc_hd__clkbuf_1
Xwire242 _04028_ VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__clkbuf_1
Xmax_length3560 _07038_ VGND VGND VPWR VPWR net3560 sky130_fd_sc_hd__buf_1
Xwire253 _08370_ VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__clkbuf_1
Xwire264 _04388_ VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__clkbuf_1
X_17032_ net1225 VGND VGND VPWR VPWR _08992_ sky130_fd_sc_hd__buf_1
X_14244_ net8062 VGND VGND VPWR VPWR _06499_ sky130_fd_sc_hd__inv_2
Xmax_length3571 net3572 VGND VGND VPWR VPWR net3571 sky130_fd_sc_hd__clkbuf_1
Xwire275 _10746_ VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__buf_1
Xwire286 _05936_ VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__clkbuf_1
Xwire7895 net7896 VGND VGND VPWR VPWR net7895 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire297 _02327_ VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__buf_1
Xmax_length2870 _06820_ VGND VGND VPWR VPWR net2870 sky130_fd_sc_hd__clkbuf_1
X_14175_ net217 _06422_ _06369_ VGND VGND VPWR VPWR _06435_ sky130_fd_sc_hd__a21o_1
Xmax_length2892 _06603_ VGND VGND VPWR VPWR net2892 sky130_fd_sc_hd__buf_1
XFILLER_0_22_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13126_ net734 _05364_ _05365_ VGND VGND VPWR VPWR _05399_ sky130_fd_sc_hd__and3_1
X_18983_ net6352 net6342 VGND VGND VPWR VPWR _10820_ sky130_fd_sc_hd__or2b_1
X_13057_ _05329_ _05209_ _05204_ VGND VGND VPWR VPWR _05330_ sky130_fd_sc_hd__mux2_1
X_17934_ net2561 net2559 net2145 net2143 VGND VGND VPWR VPWR _09785_ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17865_ net4043 _09632_ net3990 VGND VGND VPWR VPWR _09716_ sky130_fd_sc_hd__or3_1
Xwire2180 net2181 VGND VGND VPWR VPWR net2180 sky130_fd_sc_hd__buf_1
Xwire2191 net2192 VGND VGND VPWR VPWR net2191 sky130_fd_sc_hd__buf_1
X_19604_ _11438_ _11440_ VGND VGND VPWR VPWR _11441_ sky130_fd_sc_hd__xor2_2
X_16816_ _08798_ VGND VGND VPWR VPWR _00306_ sky130_fd_sc_hd__clkbuf_1
X_17796_ net3991 _09643_ _09646_ net7120 net7051 VGND VGND VPWR VPWR _09647_ sky130_fd_sc_hd__o221ai_1
Xwire1490 net1491 VGND VGND VPWR VPWR net1490 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19535_ net1060 _11342_ _11351_ VGND VGND VPWR VPWR _11372_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_187_Right_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13959_ _06219_ _06223_ VGND VGND VPWR VPWR _06224_ sky130_fd_sc_hd__xnor2_2
X_16747_ _08762_ VGND VGND VPWR VPWR _00273_ sky130_fd_sc_hd__clkbuf_1
X_19466_ _11301_ _11302_ VGND VGND VPWR VPWR _11303_ sky130_fd_sc_hd__nand2_1
X_16678_ matmul0.matmul_stage_inst.mult1\[8\] VGND VGND VPWR VPWR _08710_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18417_ _10202_ _10198_ _10257_ _10258_ VGND VGND VPWR VPWR _10267_ sky130_fd_sc_hd__o31a_1
XFILLER_0_185_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15629_ _07697_ _07700_ VGND VGND VPWR VPWR _07701_ sky130_fd_sc_hd__xnor2_1
X_19397_ net2108 _11151_ VGND VGND VPWR VPWR _11234_ sky130_fd_sc_hd__or2_1
XFILLER_0_189_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18348_ _10075_ VGND VGND VPWR VPWR _10199_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18279_ _10127_ _10128_ net1074 VGND VGND VPWR VPWR _10130_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_140_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20310_ _12112_ _12114_ VGND VGND VPWR VPWR _12115_ sky130_fd_sc_hd__xor2_1
Xinput50 currT_in[10] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_1
X_21290_ _00819_ _00820_ _00821_ VGND VGND VPWR VPWR _01305_ sky130_fd_sc_hd__o21a_1
Xinput61 currT_in[6] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput72 periodTop[1] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput83 pid_d_addr[11] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_1
X_20241_ _12057_ VGND VGND VPWR VPWR _00473_ sky130_fd_sc_hd__clkbuf_1
Xinput94 pid_d_addr[7] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3809 net3810 VGND VGND VPWR VPWR net3809 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20172_ net6078 _11997_ VGND VGND VPWR VPWR _11998_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24980_ pid_q.kp\[9\] _04720_ net1357 VGND VGND VPWR VPWR _04745_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23931_ net2411 _03794_ VGND VGND VPWR VPWR _03795_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_192_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23862_ _03724_ _03726_ VGND VGND VPWR VPWR _03727_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25601_ clknet_leaf_105_clk _00474_ net8358 VGND VGND VPWR VPWR cordic0.slte0.opB\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_22813_ net4389 net4382 net4321 net4351 VGND VGND VPWR VPWR _02716_ sky130_fd_sc_hd__nor4_1
XFILLER_0_168_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23793_ _03656_ _03658_ VGND VGND VPWR VPWR _03659_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_154_Right_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25532_ clknet_leaf_47_clk _00412_ net8776 VGND VGND VPWR VPWR svm0.state\[2\] sky130_fd_sc_hd__dfrtp_1
X_22744_ net3719 net109 VGND VGND VPWR VPWR _02674_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25463_ clknet_leaf_53_clk _00343_ net8807 VGND VGND VPWR VPWR svm0.tB\[1\] sky130_fd_sc_hd__dfrtp_1
X_22675_ pid_d.ki\[2\] net2439 net2994 pid_d.kp\[2\] VGND VGND VPWR VPWR _02625_ sky130_fd_sc_hd__a22o_1
Xfanout7008 net7026 VGND VGND VPWR VPWR net7008 sky130_fd_sc_hd__buf_1
XFILLER_0_75_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24414_ net2019 net1652 _04271_ VGND VGND VPWR VPWR _04272_ sky130_fd_sc_hd__a21oi_2
X_21626_ _01636_ _01535_ _01637_ VGND VGND VPWR VPWR _01638_ sky130_fd_sc_hd__a21o_1
X_25394_ clknet_leaf_74_clk _00277_ net8466 VGND VGND VPWR VPWR matmul0.b\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_191_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7136 net7137 VGND VGND VPWR VPWR net7136 sky130_fd_sc_hd__buf_1
X_24345_ _04200_ _04203_ VGND VGND VPWR VPWR _04204_ sky130_fd_sc_hd__xnor2_2
Xwire6402 net6403 VGND VGND VPWR VPWR net6402 sky130_fd_sc_hd__buf_1
X_21557_ _01454_ _01459_ _01452_ VGND VGND VPWR VPWR _01569_ sky130_fd_sc_hd__a21bo_1
Xfanout5617 net5623 VGND VGND VPWR VPWR net5617 sky130_fd_sc_hd__buf_1
Xwire6413 net6414 VGND VGND VPWR VPWR net6413 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire7158 net7159 VGND VGND VPWR VPWR net7158 sky130_fd_sc_hd__clkbuf_2
Xfanout5628 net5632 VGND VGND VPWR VPWR net5628 sky130_fd_sc_hd__buf_1
Xwire7169 matmul0.cos\[10\] VGND VGND VPWR VPWR net7169 sky130_fd_sc_hd__buf_1
Xwire6424 cordic0.sin\[7\] VGND VGND VPWR VPWR net6424 sky130_fd_sc_hd__clkbuf_1
Xfanout5639 pid_d.mult0.a\[0\] VGND VGND VPWR VPWR net5639 sky130_fd_sc_hd__buf_1
Xmax_length2122 net2123 VGND VGND VPWR VPWR net2122 sky130_fd_sc_hd__buf_1
Xwire6435 net6436 VGND VGND VPWR VPWR net6435 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6446 net6444 VGND VGND VPWR VPWR net6446 sky130_fd_sc_hd__dlymetal6s2s_1
X_20508_ net6841 net6824 net6790 net6762 net6521 net6491 VGND VGND VPWR VPWR _12295_
+ sky130_fd_sc_hd__mux4_2
X_24276_ net2405 _04135_ VGND VGND VPWR VPWR _04136_ sky130_fd_sc_hd__xnor2_1
Xfanout4916 net4923 VGND VGND VPWR VPWR net4916 sky130_fd_sc_hd__clkbuf_1
X_21488_ _01495_ _01500_ VGND VGND VPWR VPWR _01501_ sky130_fd_sc_hd__xnor2_2
Xwire5723 net5718 VGND VGND VPWR VPWR net5723 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire6468 net6467 VGND VGND VPWR VPWR net6468 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire5734 net5735 VGND VGND VPWR VPWR net5734 sky130_fd_sc_hd__buf_1
X_23227_ _03093_ _03096_ VGND VGND VPWR VPWR _03097_ sky130_fd_sc_hd__xnor2_2
Xwire5745 net5746 VGND VGND VPWR VPWR net5745 sky130_fd_sc_hd__buf_1
XFILLER_0_114_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5756 net5757 VGND VGND VPWR VPWR net5756 sky130_fd_sc_hd__buf_1
X_20439_ net6511 _12232_ VGND VGND VPWR VPWR _12233_ sky130_fd_sc_hd__nor2_1
Xmax_length2188 _08841_ VGND VGND VPWR VPWR net2188 sky130_fd_sc_hd__clkbuf_1
Xwire5767 net5768 VGND VGND VPWR VPWR net5767 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length1465 _09204_ VGND VGND VPWR VPWR net1465 sky130_fd_sc_hd__buf_1
Xwire5778 net5777 VGND VGND VPWR VPWR net5778 sky130_fd_sc_hd__buf_1
Xwire5789 net5790 VGND VGND VPWR VPWR net5789 sky130_fd_sc_hd__clkbuf_1
X_23158_ net5039 net4754 VGND VGND VPWR VPWR _03028_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length1498 _08916_ VGND VGND VPWR VPWR net1498 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22109_ _02095_ _02114_ VGND VGND VPWR VPWR _02115_ sky130_fd_sc_hd__nand2_1
X_15980_ net1518 _08047_ VGND VGND VPWR VPWR _08048_ sky130_fd_sc_hd__xnor2_1
X_23089_ net5001 net4694 _02957_ _02958_ VGND VGND VPWR VPWR _02959_ sky130_fd_sc_hd__a31o_1
XFILLER_0_101_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14931_ _07001_ _07004_ VGND VGND VPWR VPWR _07005_ sky130_fd_sc_hd__xnor2_1
X_17650_ net6704 svm0.tA\[11\] VGND VGND VPWR VPWR _09530_ sky130_fd_sc_hd__or2_1
X_14862_ _06948_ VGND VGND VPWR VPWR _00202_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13813_ net531 net678 VGND VGND VPWR VPWR _06081_ sky130_fd_sc_hd__and2_1
X_16601_ _08650_ VGND VGND VPWR VPWR _00239_ sky130_fd_sc_hd__clkbuf_1
X_17581_ net6712 _09461_ _09462_ VGND VGND VPWR VPWR _09463_ sky130_fd_sc_hd__a21o_1
X_14793_ net3624 net7182 net3618 VGND VGND VPWR VPWR _06913_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_82_Left_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_121_Right_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19320_ net2523 _11054_ VGND VGND VPWR VPWR _11157_ sky130_fd_sc_hd__xor2_2
X_16532_ _08547_ _08591_ VGND VGND VPWR VPWR _08592_ sky130_fd_sc_hd__xor2_1
X_13744_ _05872_ net451 VGND VGND VPWR VPWR _06012_ sky130_fd_sc_hd__and2_1
XFILLER_0_161_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19251_ _11042_ _11041_ VGND VGND VPWR VPWR _11088_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16463_ _08447_ _08464_ _08523_ VGND VGND VPWR VPWR _08524_ sky130_fd_sc_hd__a21o_1
X_13675_ _05875_ _05876_ VGND VGND VPWR VPWR _05944_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18202_ _10051_ _10052_ VGND VGND VPWR VPWR _10053_ sky130_fd_sc_hd__and2_1
X_15414_ net4087 net4086 VGND VGND VPWR VPWR _07488_ sky130_fd_sc_hd__or2_1
X_12626_ svm0.vC\[5\] net2990 net3694 net4275 VGND VGND VPWR VPWR _04899_ sky130_fd_sc_hd__a22oi_1
X_19182_ _11016_ _11013_ VGND VGND VPWR VPWR _11019_ sky130_fd_sc_hd__or2_1
X_16394_ net2791 net2772 VGND VGND VPWR VPWR _08456_ sky130_fd_sc_hd__nor2_1
Xwire8360 net8361 VGND VGND VPWR VPWR net8360 sky130_fd_sc_hd__clkbuf_1
X_18133_ _09914_ _09983_ _09922_ _09917_ VGND VGND VPWR VPWR _09984_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_81_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15345_ net2760 net2756 VGND VGND VPWR VPWR _07419_ sky130_fd_sc_hd__nor2_1
Xwire8371 net8372 VGND VGND VPWR VPWR net8371 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8382 net8380 VGND VGND VPWR VPWR net8382 sky130_fd_sc_hd__clkbuf_2
Xwire8393 net8388 VGND VGND VPWR VPWR net8393 sky130_fd_sc_hd__buf_1
X_18064_ net7087 cordic0.vec\[1\]\[1\] VGND VGND VPWR VPWR _09915_ sky130_fd_sc_hd__nand2_1
Xwire7681 net7679 VGND VGND VPWR VPWR net7681 sky130_fd_sc_hd__buf_1
X_15276_ _07155_ _07158_ _07154_ VGND VGND VPWR VPWR _07350_ sky130_fd_sc_hd__o21ba_1
Xwire7692 net7693 VGND VGND VPWR VPWR net7692 sky130_fd_sc_hd__clkbuf_1
Xhold108 pid_d.curr_error\[15\] VGND VGND VPWR VPWR net9061 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_91_Left_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17015_ net1807 net1483 VGND VGND VPWR VPWR _08976_ sky130_fd_sc_hd__and2_1
X_14227_ _06446_ _06470_ _06404_ VGND VGND VPWR VPWR _06485_ sky130_fd_sc_hd__o21ba_1
Xhold119 svm0.vC\[0\] VGND VGND VPWR VPWR net9072 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6980 cordic0.vec\[1\]\[8\] VGND VGND VPWR VPWR net6980 sky130_fd_sc_hd__buf_1
Xwire6991 net6992 VGND VGND VPWR VPWR net6991 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14158_ _06403_ _06418_ VGND VGND VPWR VPWR _06419_ sky130_fd_sc_hd__xnor2_2
X_13109_ _05253_ _05380_ _05381_ VGND VGND VPWR VPWR _05382_ sky130_fd_sc_hd__a21o_1
X_14089_ _06332_ _06351_ VGND VGND VPWR VPWR _06352_ sky130_fd_sc_hd__xnor2_2
X_18966_ net6203 net6162 VGND VGND VPWR VPWR _10803_ sky130_fd_sc_hd__xnor2_1
X_17917_ _09762_ _09764_ _09766_ _09666_ VGND VGND VPWR VPWR _09768_ sky130_fd_sc_hd__or4_1
X_18897_ _10711_ _10737_ VGND VGND VPWR VPWR _10738_ sky130_fd_sc_hd__xor2_2
X_17848_ net2145 net2143 VGND VGND VPWR VPWR _09699_ sky130_fd_sc_hd__xor2_1
XFILLER_0_178_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17779_ net6996 net3997 VGND VGND VPWR VPWR _09630_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_89_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19518_ _11294_ _11354_ VGND VGND VPWR VPWR _11355_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20790_ net5626 net5730 VGND VGND VPWR VPWR _12561_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19449_ _11284_ _11285_ VGND VGND VPWR VPWR _11286_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22460_ _02402_ _02403_ _02404_ VGND VGND VPWR VPWR _02461_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_173_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21411_ _01423_ _01424_ VGND VGND VPWR VPWR _01425_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22391_ _02262_ _02391_ _02392_ VGND VGND VPWR VPWR _02394_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24130_ net2408 _03990_ VGND VGND VPWR VPWR _03992_ sky130_fd_sc_hd__nand2_1
X_21342_ net5638 net5616 _01350_ _01355_ net5687 VGND VGND VPWR VPWR _01356_ sky130_fd_sc_hd__o32a_1
XFILLER_0_32_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5008 net5009 VGND VGND VPWR VPWR net5008 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24061_ net4640 net4669 _03372_ VGND VGND VPWR VPWR _03924_ sky130_fd_sc_hd__and3_1
Xwire4307 net4309 VGND VGND VPWR VPWR net4307 sky130_fd_sc_hd__clkbuf_1
X_21273_ _01282_ _01287_ VGND VGND VPWR VPWR _01288_ sky130_fd_sc_hd__xnor2_1
Xwire4329 net4330 VGND VGND VPWR VPWR net4329 sky130_fd_sc_hd__clkbuf_1
X_23012_ net5132 net4610 VGND VGND VPWR VPWR _02882_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20224_ net8120 _12043_ VGND VGND VPWR VPWR _12044_ sky130_fd_sc_hd__nor2_1
Xwire3606 _06950_ VGND VGND VPWR VPWR net3606 sky130_fd_sc_hd__clkbuf_2
Xwire3617 _06831_ VGND VGND VPWR VPWR net3617 sky130_fd_sc_hd__clkbuf_1
Xwire3628 net3629 VGND VGND VPWR VPWR net3628 sky130_fd_sc_hd__buf_1
Xwire3639 net3640 VGND VGND VPWR VPWR net3639 sky130_fd_sc_hd__buf_1
Xwire2905 net2906 VGND VGND VPWR VPWR net2905 sky130_fd_sc_hd__clkbuf_1
X_20155_ _11927_ net1055 _11953_ VGND VGND VPWR VPWR _11982_ sky130_fd_sc_hd__or3_1
Xwire2916 net2917 VGND VGND VPWR VPWR net2916 sky130_fd_sc_hd__clkbuf_1
Xwire2927 net2928 VGND VGND VPWR VPWR net2927 sky130_fd_sc_hd__clkbuf_1
Xwire2938 net2939 VGND VGND VPWR VPWR net2938 sky130_fd_sc_hd__clkbuf_1
Xwire2949 _05619_ VGND VGND VPWR VPWR net2949 sky130_fd_sc_hd__buf_1
X_24963_ _04736_ VGND VGND VPWR VPWR _00761_ sky130_fd_sc_hd__clkbuf_1
X_20086_ _11844_ _11873_ VGND VGND VPWR VPWR _11915_ sky130_fd_sc_hd__nand2_1
XFILLER_0_176_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_96_clk clknet_4_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_96_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23914_ _03776_ _03777_ _03758_ VGND VGND VPWR VPWR _03778_ sky130_fd_sc_hd__a21o_1
X_24894_ _04687_ VGND VGND VPWR VPWR _00741_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length8335 net8336 VGND VGND VPWR VPWR net8335 sky130_fd_sc_hd__buf_1
X_23845_ net4669 net4854 VGND VGND VPWR VPWR _03710_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length8379 net8369 VGND VGND VPWR VPWR net8379 sky130_fd_sc_hd__clkbuf_1
Xmax_length6900 net6895 VGND VGND VPWR VPWR net6900 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_169_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23776_ net1666 _03507_ _03503_ VGND VGND VPWR VPWR _03642_ sky130_fd_sc_hd__o21a_1
Xmax_length6933 net6934 VGND VGND VPWR VPWR net6933 sky130_fd_sc_hd__buf_1
X_20988_ _00996_ _01003_ VGND VGND VPWR VPWR _01004_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25515_ clknet_leaf_44_clk _00395_ net8783 VGND VGND VPWR VPWR svm0.counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_184_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22727_ pid_d.ki\[0\] _02653_ net1688 VGND VGND VPWR VPWR _02663_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6988 net6989 VGND VGND VPWR VPWR net6988 sky130_fd_sc_hd__clkbuf_1
X_13460_ net7722 net2331 net2325 VGND VGND VPWR VPWR _05733_ sky130_fd_sc_hd__and3_1
X_25446_ clknet_4_1__leaf_clk _00329_ net8334 VGND VGND VPWR VPWR cordic0.vec\[1\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_22658_ net4364 _02268_ _02600_ net940 VGND VGND VPWR VPWR _02614_ sky130_fd_sc_hd__a211o_1
Xfanout6104 cordic0.vec\[0\]\[12\] VGND VGND VPWR VPWR net6104 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21609_ _01613_ _01620_ VGND VGND VPWR VPWR _01621_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13391_ _05247_ _05245_ VGND VGND VPWR VPWR _05664_ sky130_fd_sc_hd__nor2_1
X_25377_ clknet_leaf_64_clk _00260_ net8663 VGND VGND VPWR VPWR matmul0.alpha_pass\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_22589_ net7294 _02564_ VGND VGND VPWR VPWR _02567_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_20_clk clknet_4_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_16
Xwire6210 net6211 VGND VGND VPWR VPWR net6210 sky130_fd_sc_hd__clkbuf_1
Xfanout6159 net6165 VGND VGND VPWR VPWR net6159 sky130_fd_sc_hd__buf_1
X_15130_ _07149_ VGND VGND VPWR VPWR _07204_ sky130_fd_sc_hd__clkbuf_1
X_24328_ pid_q.prev_int\[10\] VGND VGND VPWR VPWR _04187_ sky130_fd_sc_hd__inv_2
XFILLER_0_161_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout5436 net5452 VGND VGND VPWR VPWR net5436 sky130_fd_sc_hd__clkbuf_1
Xwire6232 net6228 VGND VGND VPWR VPWR net6232 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire6254 net6255 VGND VGND VPWR VPWR net6254 sky130_fd_sc_hd__buf_1
Xfanout4724 pid_q.mult0.a\[3\] VGND VGND VPWR VPWR net4724 sky130_fd_sc_hd__clkbuf_1
Xwire5520 net5521 VGND VGND VPWR VPWR net5520 sky130_fd_sc_hd__clkbuf_1
Xwire5531 net5523 VGND VGND VPWR VPWR net5531 sky130_fd_sc_hd__clkbuf_1
X_15061_ net6540 net6592 VGND VGND VPWR VPWR _07135_ sky130_fd_sc_hd__or2_1
X_24259_ _04048_ net589 VGND VGND VPWR VPWR _04119_ sky130_fd_sc_hd__or2_1
Xwire5542 net5543 VGND VGND VPWR VPWR net5542 sky130_fd_sc_hd__buf_1
Xwire6298 net6300 VGND VGND VPWR VPWR net6298 sky130_fd_sc_hd__buf_1
X_14012_ _06157_ _06215_ _06269_ _06273_ VGND VGND VPWR VPWR _06276_ sky130_fd_sc_hd__a31o_1
Xwire5564 net5567 VGND VGND VPWR VPWR net5564 sky130_fd_sc_hd__buf_1
Xwire4830 net4831 VGND VGND VPWR VPWR net4830 sky130_fd_sc_hd__clkbuf_1
Xfanout4779 pid_q.mult0.a\[0\] VGND VGND VPWR VPWR net4779 sky130_fd_sc_hd__buf_1
Xwire4852 net4853 VGND VGND VPWR VPWR net4852 sky130_fd_sc_hd__buf_1
Xwire5597 net5598 VGND VGND VPWR VPWR net5597 sky130_fd_sc_hd__buf_1
Xwire4863 net4864 VGND VGND VPWR VPWR net4863 sky130_fd_sc_hd__clkbuf_1
X_18820_ _10627_ _10649_ _10662_ VGND VGND VPWR VPWR _10663_ sky130_fd_sc_hd__o21ai_1
Xwire4896 net4894 VGND VGND VPWR VPWR net4896 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18751_ _10520_ _10549_ _10550_ VGND VGND VPWR VPWR _10596_ sky130_fd_sc_hd__o21ai_2
X_15963_ _08025_ _08030_ VGND VGND VPWR VPWR _08031_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_87_clk clknet_4_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_87_clk sky130_fd_sc_hd__clkbuf_16
X_17702_ _04869_ _09577_ VGND VGND VPWR VPWR _09578_ sky130_fd_sc_hd__or2_1
X_14914_ _06987_ VGND VGND VPWR VPWR _06988_ sky130_fd_sc_hd__buf_1
X_15894_ net2647 net2765 VGND VGND VPWR VPWR _07963_ sky130_fd_sc_hd__nor2_1
X_18682_ net6893 net2131 _10475_ VGND VGND VPWR VPWR _10528_ sky130_fd_sc_hd__or3_1
XFILLER_0_175_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17633_ net6699 _09512_ _09513_ VGND VGND VPWR VPWR _09514_ sky130_fd_sc_hd__a21oi_1
X_14845_ matmul0.a\[11\] matmul0.matmul_stage_inst.e\[11\] net3607 VGND VGND VPWR
+ VPWR _06940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17564_ svm0.tC\[1\] VGND VGND VPWR VPWR _09446_ sky130_fd_sc_hd__inv_2
X_14776_ net9040 net2857 net2866 _06901_ VGND VGND VPWR VPWR _00163_ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19303_ net6292 net6244 VGND VGND VPWR VPWR _11140_ sky130_fd_sc_hd__xnor2_2
X_13727_ _05921_ _05924_ _05995_ VGND VGND VPWR VPWR _05996_ sky130_fd_sc_hd__a21oi_1
X_16515_ _08511_ _08513_ VGND VGND VPWR VPWR _08575_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17495_ svm0.delta\[9\] _09383_ VGND VGND VPWR VPWR _09384_ sky130_fd_sc_hd__xnor2_1
X_19234_ net6230 net6340 _11024_ VGND VGND VPWR VPWR _11071_ sky130_fd_sc_hd__o21ba_1
X_13658_ _05806_ _05833_ net681 VGND VGND VPWR VPWR _05928_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16446_ _08389_ _08506_ _08387_ VGND VGND VPWR VPWR _08507_ sky130_fd_sc_hd__a21o_1
XFILLER_0_184_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12609_ net3697 VGND VGND VPWR VPWR _00000_ sky130_fd_sc_hd__clkbuf_1
X_19165_ _11000_ _11001_ VGND VGND VPWR VPWR _11002_ sky130_fd_sc_hd__nand2_1
X_16377_ _08408_ net1079 VGND VGND VPWR VPWR _08439_ sky130_fd_sc_hd__nand2_1
X_13589_ _05771_ _05849_ VGND VGND VPWR VPWR _05859_ sky130_fd_sc_hd__and2b_1
XFILLER_0_54_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_11_clk clknet_4_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_182_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8190 net8191 VGND VGND VPWR VPWR net8190 sky130_fd_sc_hd__clkbuf_1
X_15328_ _07387_ _07401_ VGND VGND VPWR VPWR _07402_ sky130_fd_sc_hd__xnor2_4
X_18116_ net3235 _09867_ _09966_ VGND VGND VPWR VPWR _09967_ sky130_fd_sc_hd__o21ai_1
Xfanout6660 net6671 VGND VGND VPWR VPWR net6660 sky130_fd_sc_hd__buf_1
XFILLER_0_83_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19096_ net2527 _10855_ VGND VGND VPWR VPWR _10933_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18047_ _09856_ _09883_ VGND VGND VPWR VPWR _09898_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15259_ _07297_ _07332_ VGND VGND VPWR VPWR _07333_ sky130_fd_sc_hd__and2_1
X_19998_ net350 _11825_ _11782_ VGND VGND VPWR VPWR _11829_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_129_Left_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18949_ net9073 net2121 net1446 _10786_ VGND VGND VPWR VPWR _00452_ sky130_fd_sc_hd__a31o_1
XFILLER_0_193_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_78_clk clknet_4_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_78_clk sky130_fd_sc_hd__clkbuf_16
X_21960_ net1713 _01967_ VGND VGND VPWR VPWR _01968_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20911_ net1392 net1187 _00926_ VGND VGND VPWR VPWR _00927_ sky130_fd_sc_hd__a21oi_1
X_21891_ net2063 _01897_ VGND VGND VPWR VPWR _01900_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23630_ net4703 net4846 VGND VGND VPWR VPWR _03497_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20842_ _00850_ _00857_ VGND VGND VPWR VPWR _00858_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_166_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23561_ _03427_ _03428_ VGND VGND VPWR VPWR _03429_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20773_ net5596 net5776 VGND VGND VPWR VPWR _12544_ sky130_fd_sc_hd__nand2_1
X_25300_ clknet_leaf_76_clk _00183_ net8460 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.e\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_22512_ _02456_ _02457_ net517 VGND VGND VPWR VPWR _02513_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_138_Left_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23492_ _03357_ _03360_ VGND VGND VPWR VPWR _03361_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_36_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25231_ clknet_leaf_64_clk _00120_ net8661 VGND VGND VPWR VPWR matmul0.start sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire808 _01076_ VGND VGND VPWR VPWR net808 sky130_fd_sc_hd__buf_1
X_22443_ _02228_ net2470 _02444_ net5765 VGND VGND VPWR VPWR _02445_ sky130_fd_sc_hd__a22o_1
Xwire819 _09972_ VGND VGND VPWR VPWR net819 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25162_ clknet_leaf_54_clk _00051_ net8730 VGND VGND VPWR VPWR svm0.periodTop\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_22374_ _02371_ _02376_ VGND VGND VPWR VPWR _02377_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24113_ _03968_ _03974_ VGND VGND VPWR VPWR _03975_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_60_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21325_ _01337_ _01338_ VGND VGND VPWR VPWR _01339_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25093_ net4401 net5172 _04824_ net5174 net4406 VGND VGND VPWR VPWR _04837_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4104 _07132_ VGND VGND VPWR VPWR net4104 sky130_fd_sc_hd__clkbuf_1
Xwire4115 net4117 VGND VGND VPWR VPWR net4115 sky130_fd_sc_hd__buf_1
Xwire4126 net4127 VGND VGND VPWR VPWR net4126 sky130_fd_sc_hd__buf_1
X_24044_ _03899_ _03905_ VGND VGND VPWR VPWR _03907_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4137 net4138 VGND VGND VPWR VPWR net4137 sky130_fd_sc_hd__buf_1
X_21256_ _00844_ _00848_ net2483 VGND VGND VPWR VPWR _01271_ sky130_fd_sc_hd__o21a_1
Xwire4148 net4149 VGND VGND VPWR VPWR net4148 sky130_fd_sc_hd__buf_1
Xwire3403 _07598_ VGND VGND VPWR VPWR net3403 sky130_fd_sc_hd__clkbuf_1
Xwire4159 _07010_ VGND VGND VPWR VPWR net4159 sky130_fd_sc_hd__buf_1
Xwire3414 net3419 VGND VGND VPWR VPWR net3414 sky130_fd_sc_hd__buf_1
Xwire3425 net3426 VGND VGND VPWR VPWR net3425 sky130_fd_sc_hd__buf_1
XFILLER_0_187_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20207_ net9046 net2123 net1445 _12031_ VGND VGND VPWR VPWR _00465_ sky130_fd_sc_hd__a31o_1
Xwire3436 net3437 VGND VGND VPWR VPWR net3436 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_147_Left_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2702 _07368_ VGND VGND VPWR VPWR net2702 sky130_fd_sc_hd__buf_1
Xwire3447 net3448 VGND VGND VPWR VPWR net3447 sky130_fd_sc_hd__buf_1
XFILLER_0_99_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21187_ _01157_ _01161_ _01148_ VGND VGND VPWR VPWR _01203_ sky130_fd_sc_hd__a21bo_1
Xwire3458 net3460 VGND VGND VPWR VPWR net3458 sky130_fd_sc_hd__buf_1
XFILLER_0_25_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2724 net2725 VGND VGND VPWR VPWR net2724 sky130_fd_sc_hd__buf_1
Xwire3469 net3470 VGND VGND VPWR VPWR net3469 sky130_fd_sc_hd__clkbuf_1
Xwire2735 net2736 VGND VGND VPWR VPWR net2735 sky130_fd_sc_hd__buf_1
Xwire2746 net2747 VGND VGND VPWR VPWR net2746 sky130_fd_sc_hd__buf_1
X_20138_ net1439 _11965_ VGND VGND VPWR VPWR _11966_ sky130_fd_sc_hd__nor2_1
Xwire2757 _07204_ VGND VGND VPWR VPWR net2757 sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_69_clk clknet_4_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_69_clk sky130_fd_sc_hd__clkbuf_16
Xwire2768 net2769 VGND VGND VPWR VPWR net2768 sky130_fd_sc_hd__clkbuf_2
X_24946_ pid_q.ki\[11\] _04724_ net1636 VGND VGND VPWR VPWR _04725_ sky130_fd_sc_hd__mux2_1
X_12960_ _05224_ _05232_ VGND VGND VPWR VPWR _05233_ sky130_fd_sc_hd__nor2_1
X_20069_ _11863_ net2494 VGND VGND VPWR VPWR _11898_ sky130_fd_sc_hd__nor2_1
Xmax_length8121 net8120 VGND VGND VPWR VPWR net8121 sky130_fd_sc_hd__clkbuf_2
X_24877_ pid_q.ki\[7\] net2397 net3009 pid_q.kp\[7\] VGND VGND VPWR VPWR _04676_ sky130_fd_sc_hd__a22o_1
X_12891_ _05160_ _05161_ _05162_ _05163_ VGND VGND VPWR VPWR _05164_ sky130_fd_sc_hd__a211o_1
XFILLER_0_99_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14630_ net8992 _06797_ _06523_ VGND VGND VPWR VPWR _00121_ sky130_fd_sc_hd__o21a_1
Xmax_length7431 matmul0.matmul_stage_inst.b\[4\] VGND VGND VPWR VPWR net7431 sky130_fd_sc_hd__clkbuf_1
X_23828_ _03685_ _03692_ VGND VGND VPWR VPWR _03693_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_157_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length7464 net7465 VGND VGND VPWR VPWR net7464 sky130_fd_sc_hd__buf_1
XFILLER_0_157_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14561_ net5223 _06731_ VGND VGND VPWR VPWR _06738_ sky130_fd_sc_hd__and2_1
X_23759_ net4636 net4899 VGND VGND VPWR VPWR _03625_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_156_Left_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length7497 net7498 VGND VGND VPWR VPWR net7497 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6763 net6764 VGND VGND VPWR VPWR net6763 sky130_fd_sc_hd__buf_1
XFILLER_0_71_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13512_ _05698_ net622 _05782_ VGND VGND VPWR VPWR _05783_ sky130_fd_sc_hd__o21a_1
X_16300_ net491 _08299_ _08297_ VGND VGND VPWR VPWR _08364_ sky130_fd_sc_hd__a21oi_1
X_17280_ _08646_ net4067 VGND VGND VPWR VPWR _09195_ sky130_fd_sc_hd__nor2_1
X_14492_ _06674_ _06675_ VGND VGND VPWR VPWR _06676_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16231_ _08256_ _08295_ VGND VGND VPWR VPWR _08296_ sky130_fd_sc_hd__xor2_2
XFILLER_0_82_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13443_ net7745 net1963 _05506_ VGND VGND VPWR VPWR _05716_ sky130_fd_sc_hd__and3_1
X_25429_ clknet_leaf_98_clk _00312_ net8384 VGND VGND VPWR VPWR matmul0.sin\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16162_ _08138_ _08148_ VGND VGND VPWR VPWR _08228_ sky130_fd_sc_hd__nand2_1
X_13374_ _05538_ _05638_ VGND VGND VPWR VPWR _05647_ sky130_fd_sc_hd__nand2_1
XFILLER_0_181_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15113_ _07116_ _07117_ VGND VGND VPWR VPWR _07187_ sky130_fd_sc_hd__xnor2_1
Xwire6062 net6058 VGND VGND VPWR VPWR net6062 sky130_fd_sc_hd__buf_1
X_16093_ _08158_ _08159_ VGND VGND VPWR VPWR _08160_ sky130_fd_sc_hd__nor2_1
Xwire6073 net6074 VGND VGND VPWR VPWR net6073 sky130_fd_sc_hd__buf_1
Xmax_length995 _06542_ VGND VGND VPWR VPWR net995 sky130_fd_sc_hd__buf_1
Xwire6095 net6091 VGND VGND VPWR VPWR net6095 sky130_fd_sc_hd__buf_1
X_19921_ net3916 _11748_ _11751_ _11752_ VGND VGND VPWR VPWR _11753_ sky130_fd_sc_hd__o211a_1
X_15044_ net4195 net4193 VGND VGND VPWR VPWR _07118_ sky130_fd_sc_hd__or2_1
Xwire5361 net5362 VGND VGND VPWR VPWR net5361 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_165_Left_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5372 pid_d.kp\[15\] VGND VGND VPWR VPWR net5372 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5383 net5384 VGND VGND VPWR VPWR net5383 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4660 net4668 VGND VGND VPWR VPWR net4660 sky130_fd_sc_hd__clkbuf_1
Xwire4671 net4672 VGND VGND VPWR VPWR net4671 sky130_fd_sc_hd__clkbuf_1
X_19852_ net3165 _11680_ _11682_ _11683_ _11684_ VGND VGND VPWR VPWR _11685_ sky130_fd_sc_hd__o221a_1
Xwire4682 net4683 VGND VGND VPWR VPWR net4682 sky130_fd_sc_hd__clkbuf_1
Xwire4693 net4694 VGND VGND VPWR VPWR net4693 sky130_fd_sc_hd__buf_1
X_18803_ _10636_ _10646_ VGND VGND VPWR VPWR _10647_ sky130_fd_sc_hd__xnor2_2
Xwire3970 net3971 VGND VGND VPWR VPWR net3970 sky130_fd_sc_hd__buf_1
X_19783_ _11609_ net604 _11542_ VGND VGND VPWR VPWR _11617_ sky130_fd_sc_hd__nand3b_1
Xwire3981 net3982 VGND VGND VPWR VPWR net3981 sky130_fd_sc_hd__buf_1
X_16995_ net6460 net2189 _08953_ _08956_ VGND VGND VPWR VPWR _08957_ sky130_fd_sc_hd__o31a_1
Xwire3992 _09636_ VGND VGND VPWR VPWR net3992 sky130_fd_sc_hd__clkbuf_1
X_18734_ net6784 _10349_ VGND VGND VPWR VPWR _10579_ sky130_fd_sc_hd__xnor2_2
X_15946_ _07926_ _08012_ _08013_ VGND VGND VPWR VPWR _08014_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_0_clk clknet_4_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_16
X_18665_ net1437 net246 VGND VGND VPWR VPWR _10512_ sky130_fd_sc_hd__nor2_1
X_15877_ net1845 net1842 VGND VGND VPWR VPWR _07946_ sky130_fd_sc_hd__nor2_1
X_17616_ net6739 svm0.tB\[0\] VGND VGND VPWR VPWR _09497_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_174_Left_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14828_ matmul0.a\[3\] matmul0.matmul_stage_inst.e\[3\] net3610 VGND VGND VPWR VPWR
+ _06931_ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18596_ net6771 net2129 _10443_ net6818 VGND VGND VPWR VPWR _10444_ sky130_fd_sc_hd__o22a_1
XFILLER_0_25_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17547_ _09420_ _09424_ _09428_ VGND VGND VPWR VPWR _09429_ sky130_fd_sc_hd__nor3_1
XFILLER_0_19_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14759_ net8955 net2867 _06889_ VGND VGND VPWR VPWR _00158_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_74_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17478_ net6718 net2576 VGND VGND VPWR VPWR _09370_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19217_ net6271 net6224 VGND VGND VPWR VPWR _11054_ sky130_fd_sc_hd__xor2_2
XFILLER_0_73_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16429_ _08490_ VGND VGND VPWR VPWR _00227_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19148_ net6267 net6300 VGND VGND VPWR VPWR _10985_ sky130_fd_sc_hd__and2b_1
XFILLER_0_14_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_183_Left_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19079_ net6268 _10911_ VGND VGND VPWR VPWR _10916_ sky130_fd_sc_hd__nand2_1
X_21110_ _01119_ _01125_ VGND VGND VPWR VPWR _01126_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_23_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22090_ _02093_ _02094_ VGND VGND VPWR VPWR _02097_ sky130_fd_sc_hd__and2_1
XFILLER_0_140_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21041_ _01055_ _01056_ net3841 VGND VGND VPWR VPWR _01057_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2009 net2010 VGND VGND VPWR VPWR net2009 sky130_fd_sc_hd__buf_1
XFILLER_0_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1308 net1309 VGND VGND VPWR VPWR net1308 sky130_fd_sc_hd__buf_1
XFILLER_0_157_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1319 _05687_ VGND VGND VPWR VPWR net1319 sky130_fd_sc_hd__buf_1
X_24800_ net259 VGND VGND VPWR VPWR _04625_ sky130_fd_sc_hd__inv_2
X_25780_ clknet_leaf_73_clk _00653_ net8499 VGND VGND VPWR VPWR matmul0.beta_pass\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_22992_ matmul0.beta_pass\[15\] _08750_ net6575 VGND VGND VPWR VPWR _02864_ sky130_fd_sc_hd__mux2_1
X_24731_ _04562_ net8012 _04552_ net8017 _04555_ VGND VGND VPWR VPWR _04564_ sky130_fd_sc_hd__a221o_1
X_21943_ _01948_ _01950_ VGND VGND VPWR VPWR _01951_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24662_ net9178 net1377 _04513_ VGND VGND VPWR VPWR _00683_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21874_ net1048 net1172 VGND VGND VPWR VPWR _01883_ sky130_fd_sc_hd__nor2_1
X_23613_ net7527 _03393_ net514 net7468 net2414 VGND VGND VPWR VPWR _03481_ sky130_fd_sc_hd__a221o_1
X_20825_ net5774 net5570 VGND VGND VPWR VPWR _00841_ sky130_fd_sc_hd__nand2_1
X_24593_ pid_q.prev_error\[13\] net5166 VGND VGND VPWR VPWR _04449_ sky130_fd_sc_hd__nor2_1
X_23544_ net4597 net4996 VGND VGND VPWR VPWR _03412_ sky130_fd_sc_hd__nand2_1
Xwire8926 net8927 VGND VGND VPWR VPWR net8926 sky130_fd_sc_hd__clkbuf_1
X_20756_ net5491 net5906 VGND VGND VPWR VPWR _12527_ sky130_fd_sc_hd__nand2_1
Xwire8937 net8938 VGND VGND VPWR VPWR net8937 sky130_fd_sc_hd__clkbuf_1
Xwire8948 net8949 VGND VGND VPWR VPWR net8948 sky130_fd_sc_hd__clkbuf_1
Xwire605 _10413_ VGND VGND VPWR VPWR net605 sky130_fd_sc_hd__dlymetal6s2s_1
X_23475_ _03272_ _03273_ _03274_ VGND VGND VPWR VPWR _03344_ sky130_fd_sc_hd__o21a_1
XFILLER_0_52_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20687_ net3143 _12461_ _12462_ VGND VGND VPWR VPWR _00514_ sky130_fd_sc_hd__a21oi_1
Xmax_length4679 net4673 VGND VGND VPWR VPWR net4679 sky130_fd_sc_hd__buf_1
Xwire627 _05685_ VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25214_ clknet_leaf_61_clk _00103_ net8717 VGND VGND VPWR VPWR svm0.vC\[2\] sky130_fd_sc_hd__dfrtp_1
Xwire649 net650 VGND VGND VPWR VPWR net649 sky130_fd_sc_hd__clkbuf_1
X_22426_ _02424_ _02427_ VGND VGND VPWR VPWR _02428_ sky130_fd_sc_hd__xor2_1
XFILLER_0_66_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25145_ clknet_leaf_104_clk _00034_ net8363 VGND VGND VPWR VPWR cordic0.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_22357_ _02290_ _02295_ _02359_ VGND VGND VPWR VPWR _02360_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21308_ _00860_ _00875_ _01322_ VGND VGND VPWR VPWR _01323_ sky130_fd_sc_hd__o21a_1
X_13090_ _05262_ _05277_ _05264_ VGND VGND VPWR VPWR _05363_ sky130_fd_sc_hd__a21bo_1
X_25076_ net5176 VGND VGND VPWR VPWR _04822_ sky130_fd_sc_hd__inv_2
X_22288_ net5465 net5670 VGND VGND VPWR VPWR _02292_ sky130_fd_sc_hd__nand2_1
Xwire3200 net3201 VGND VGND VPWR VPWR net3200 sky130_fd_sc_hd__buf_1
Xwire3211 net3212 VGND VGND VPWR VPWR net3211 sky130_fd_sc_hd__buf_1
X_24027_ _03872_ _03889_ VGND VGND VPWR VPWR _03890_ sky130_fd_sc_hd__xnor2_1
Xhold280 cordic0.cos\[13\] VGND VGND VPWR VPWR net9233 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3222 net3224 VGND VGND VPWR VPWR net3222 sky130_fd_sc_hd__buf_1
X_21239_ net759 _01253_ VGND VGND VPWR VPWR _01254_ sky130_fd_sc_hd__nor2_1
Xhold291 svm0.calc_ready VGND VGND VPWR VPWR net9244 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3233 _10047_ VGND VGND VPWR VPWR net3233 sky130_fd_sc_hd__buf_1
Xwire3244 _09737_ VGND VGND VPWR VPWR net3244 sky130_fd_sc_hd__clkbuf_1
Xwire2510 _11158_ VGND VGND VPWR VPWR net2510 sky130_fd_sc_hd__buf_1
Xwire3255 net3256 VGND VGND VPWR VPWR net3255 sky130_fd_sc_hd__buf_1
Xwire2521 _10980_ VGND VGND VPWR VPWR net2521 sky130_fd_sc_hd__buf_1
Xwire2532 net2533 VGND VGND VPWR VPWR net2532 sky130_fd_sc_hd__buf_1
XFILLER_0_46_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2543 _10177_ VGND VGND VPWR VPWR net2543 sky130_fd_sc_hd__buf_1
Xwire3288 net3289 VGND VGND VPWR VPWR net3288 sky130_fd_sc_hd__clkbuf_1
Xwire3299 net3300 VGND VGND VPWR VPWR net3299 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2565 _09563_ VGND VGND VPWR VPWR net2565 sky130_fd_sc_hd__clkbuf_1
X_15800_ _07778_ _07779_ _07781_ VGND VGND VPWR VPWR _07870_ sky130_fd_sc_hd__a21o_1
Xwire1820 net1821 VGND VGND VPWR VPWR net1820 sky130_fd_sc_hd__buf_1
Xwire2576 net2577 VGND VGND VPWR VPWR net2576 sky130_fd_sc_hd__buf_1
Xwire1831 net1833 VGND VGND VPWR VPWR net1831 sky130_fd_sc_hd__dlymetal6s2s_1
X_13992_ _06249_ _06256_ VGND VGND VPWR VPWR _06257_ sky130_fd_sc_hd__xor2_1
Xwire1842 net1843 VGND VGND VPWR VPWR net1842 sky130_fd_sc_hd__buf_1
X_16780_ _08779_ VGND VGND VPWR VPWR _00289_ sky130_fd_sc_hd__clkbuf_1
Xwire2587 _09158_ VGND VGND VPWR VPWR net2587 sky130_fd_sc_hd__buf_1
Xwire2598 _09033_ VGND VGND VPWR VPWR net2598 sky130_fd_sc_hd__buf_1
Xwire1853 _07621_ VGND VGND VPWR VPWR net1853 sky130_fd_sc_hd__buf_1
Xwire1864 _07491_ VGND VGND VPWR VPWR net1864 sky130_fd_sc_hd__buf_1
X_12943_ net1974 net1971 VGND VGND VPWR VPWR _05216_ sky130_fd_sc_hd__and2_1
X_15731_ net888 _07667_ _07801_ VGND VGND VPWR VPWR _07802_ sky130_fd_sc_hd__a21oi_2
Xwire1875 net1876 VGND VGND VPWR VPWR net1875 sky130_fd_sc_hd__clkbuf_2
X_24929_ _04713_ VGND VGND VPWR VPWR _00750_ sky130_fd_sc_hd__clkbuf_1
Xwire1886 net1887 VGND VGND VPWR VPWR net1886 sky130_fd_sc_hd__buf_1
Xwire1897 _07068_ VGND VGND VPWR VPWR net1897 sky130_fd_sc_hd__clkbuf_1
X_18450_ net6988 net7076 VGND VGND VPWR VPWR _10300_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12874_ _05032_ _05084_ _05146_ VGND VGND VPWR VPWR _05147_ sky130_fd_sc_hd__o21a_1
X_15662_ _07710_ _07733_ VGND VGND VPWR VPWR _07734_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17401_ _09303_ net616 net1461 _09306_ VGND VGND VPWR VPWR _00383_ sky130_fd_sc_hd__a31o_1
XFILLER_0_157_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14613_ _06512_ net6443 VGND VGND VPWR VPWR _06785_ sky130_fd_sc_hd__or2_1
XFILLER_0_139_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15593_ _07617_ _07663_ _07664_ VGND VGND VPWR VPWR _07665_ sky130_fd_sc_hd__o21ai_1
X_18381_ net7012 _09909_ VGND VGND VPWR VPWR _10232_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17332_ _09207_ _09244_ _09245_ VGND VGND VPWR VPWR _09246_ sky130_fd_sc_hd__mux2_1
X_14544_ net7278 net5250 _06711_ VGND VGND VPWR VPWR _06723_ sky130_fd_sc_hd__or3_1
XFILLER_0_28_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length6571 net6567 VGND VGND VPWR VPWR net6571 sky130_fd_sc_hd__buf_1
XFILLER_0_138_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17263_ net2156 VGND VGND VPWR VPWR _09194_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14475_ _06660_ _06661_ VGND VGND VPWR VPWR _06662_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19002_ net6267 net6300 VGND VGND VPWR VPWR _10839_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13426_ _05590_ net844 VGND VGND VPWR VPWR _05699_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16214_ _08277_ _08278_ VGND VGND VPWR VPWR _08279_ sky130_fd_sc_hd__nor2_1
X_17194_ net2597 _09143_ VGND VGND VPWR VPWR _09144_ sky130_fd_sc_hd__or2_1
XFILLER_0_183_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16145_ _08131_ _08136_ net776 VGND VGND VPWR VPWR _08211_ sky130_fd_sc_hd__o21a_1
X_13357_ net1330 _05536_ _05524_ VGND VGND VPWR VPWR _05630_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_106_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16076_ _08141_ _08142_ net3460 VGND VGND VPWR VPWR _08143_ sky130_fd_sc_hd__a21oi_1
X_13288_ net733 _05559_ _05560_ VGND VGND VPWR VPWR _05561_ sky130_fd_sc_hd__a21o_1
X_15027_ net4181 net4179 VGND VGND VPWR VPWR _07101_ sky130_fd_sc_hd__or2_1
X_19904_ net3127 net351 VGND VGND VPWR VPWR _11736_ sky130_fd_sc_hd__nor2_1
Xwire5191 net5192 VGND VGND VPWR VPWR net5191 sky130_fd_sc_hd__clkbuf_1
Xwire4490 net4487 VGND VGND VPWR VPWR net4490 sky130_fd_sc_hd__dlymetal6s2s_1
X_19835_ _11601_ _11604_ _11668_ VGND VGND VPWR VPWR _11669_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19766_ _11500_ _11530_ _11529_ VGND VGND VPWR VPWR _11601_ sky130_fd_sc_hd__a21o_1
X_16978_ net1918 net878 net8069 VGND VGND VPWR VPWR _08941_ sky130_fd_sc_hd__o21a_1
Xinput4 angle_in[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
XFILLER_0_78_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18717_ _10493_ net1195 _10562_ VGND VGND VPWR VPWR _10563_ sky130_fd_sc_hd__o21ai_1
X_15929_ _07892_ _07905_ VGND VGND VPWR VPWR _07998_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19697_ _11443_ _11470_ _11441_ VGND VGND VPWR VPWR _11533_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18648_ _10441_ net1069 _10494_ VGND VGND VPWR VPWR _10495_ sky130_fd_sc_hd__a21o_1
XFILLER_0_93_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18579_ net6934 _10364_ _10424_ _10425_ _10426_ VGND VGND VPWR VPWR _10427_ sky130_fd_sc_hd__a41o_1
XFILLER_0_15_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20610_ net1396 _12384_ _12388_ _12366_ _12390_ VGND VGND VPWR VPWR _12391_ sky130_fd_sc_hd__o221a_1
XFILLER_0_145_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21590_ net1177 _01601_ VGND VGND VPWR VPWR _01602_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_188_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20541_ net1484 net2082 net2079 net3193 VGND VGND VPWR VPWR _12326_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6809 net6807 VGND VGND VPWR VPWR net6809 sky130_fd_sc_hd__clkbuf_2
X_23260_ _03114_ _03129_ VGND VGND VPWR VPWR _03130_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20472_ net8044 _12224_ _12258_ cordic0.slte0.opA\[17\] net2178 VGND VGND VPWR VPWR
+ _12262_ sky130_fd_sc_hd__a32o_1
XFILLER_0_172_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22211_ net5726 net5409 VGND VGND VPWR VPWR _02216_ sky130_fd_sc_hd__nand2_1
X_23191_ _03053_ _03056_ _03060_ VGND VGND VPWR VPWR _03061_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_131_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22142_ _02038_ _02049_ _02036_ VGND VGND VPWR VPWR _02148_ sky130_fd_sc_hd__o21a_1
XFILLER_0_168_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22073_ net802 _02079_ VGND VGND VPWR VPWR _02080_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25901_ clknet_leaf_17_clk _00774_ net8630 VGND VGND VPWR VPWR pid_q.kp\[13\] sky130_fd_sc_hd__dfrtp_1
X_21024_ _01037_ _01038_ _01039_ VGND VGND VPWR VPWR _01040_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_22_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1105 net1106 VGND VGND VPWR VPWR net1105 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1116 _07428_ VGND VGND VPWR VPWR net1116 sky130_fd_sc_hd__buf_1
Xwire1127 _05780_ VGND VGND VPWR VPWR net1127 sky130_fd_sc_hd__clkbuf_2
X_25832_ clknet_leaf_36_clk _00705_ net8753 VGND VGND VPWR VPWR pid_q.curr_error\[8\]
+ sky130_fd_sc_hd__dfrtp_2
Xwire1138 net1139 VGND VGND VPWR VPWR net1138 sky130_fd_sc_hd__buf_1
XFILLER_0_96_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1149 net1151 VGND VGND VPWR VPWR net1149 sky130_fd_sc_hd__buf_1
X_22975_ _02855_ VGND VGND VPWR VPWR _00654_ sky130_fd_sc_hd__clkbuf_1
X_25763_ clknet_leaf_67_clk _00636_ net8455 VGND VGND VPWR VPWR pid_d.out\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_184_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24714_ pid_q.curr_error\[2\] net1368 net1365 net1010 VGND VGND VPWR VPWR _00699_
+ sky130_fd_sc_hd__a22o_1
X_21926_ net5710 net5499 VGND VGND VPWR VPWR _01934_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25694_ clknet_leaf_121_clk _00567_ net8395 VGND VGND VPWR VPWR pid_d.mult0.b\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24645_ net263 _04498_ _04499_ VGND VGND VPWR VPWR _04500_ sky130_fd_sc_hd__o21a_1
X_21857_ net5839 VGND VGND VPWR VPWR _01866_ sky130_fd_sc_hd__inv_2
Xfanout8617 net8622 VGND VGND VPWR VPWR net8617 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_77_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20808_ _12504_ _12505_ _12506_ VGND VGND VPWR VPWR _00824_ sky130_fd_sc_hd__o21ai_1
X_24576_ net4894 net4871 _04347_ VGND VGND VPWR VPWR _04432_ sky130_fd_sc_hd__a21o_1
Xfanout7905 net7925 VGND VGND VPWR VPWR net7905 sky130_fd_sc_hd__buf_1
X_12590_ _04865_ _04872_ VGND VGND VPWR VPWR _04873_ sky130_fd_sc_hd__nor2_1
Xmax_length5144 net5145 VGND VGND VPWR VPWR net5144 sky130_fd_sc_hd__clkbuf_1
X_21788_ _01797_ VGND VGND VPWR VPWR _01798_ sky130_fd_sc_hd__clkbuf_1
Xwire8723 net8724 VGND VGND VPWR VPWR net8723 sky130_fd_sc_hd__clkbuf_2
Xmax_length5166 pid_q.curr_error\[13\] VGND VGND VPWR VPWR net5166 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire8734 net8735 VGND VGND VPWR VPWR net8734 sky130_fd_sc_hd__clkbuf_1
X_23527_ net5129 net4512 VGND VGND VPWR VPWR _03395_ sky130_fd_sc_hd__nand2_1
Xwire8745 net8743 VGND VGND VPWR VPWR net8745 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20739_ net5545 net5838 VGND VGND VPWR VPWR _12510_ sky130_fd_sc_hd__nand2_1
Xwire402 _07922_ VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire413 net414 VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__buf_1
XFILLER_0_136_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire424 _08240_ VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__buf_1
Xwire8789 net8786 VGND VGND VPWR VPWR net8789 sky130_fd_sc_hd__buf_1
X_14260_ net4236 _06513_ net3666 VGND VGND VPWR VPWR _06514_ sky130_fd_sc_hd__o21ba_1
Xwire435 net436 VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__clkbuf_1
X_23458_ _03265_ _03266_ _03267_ VGND VGND VPWR VPWR _03327_ sky130_fd_sc_hd__o21ai_1
Xmax_length3742 _03705_ VGND VGND VPWR VPWR net3742 sky130_fd_sc_hd__buf_1
Xwire446 net447 VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire457 net458 VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__buf_1
XFILLER_0_107_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire468 net469 VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__clkbuf_1
X_13211_ _05431_ _05479_ VGND VGND VPWR VPWR _05484_ sky130_fd_sc_hd__and2_1
X_22409_ _02337_ _02409_ _02410_ VGND VGND VPWR VPWR _02411_ sky130_fd_sc_hd__a21o_1
Xmax_length3775 _02541_ VGND VGND VPWR VPWR net3775 sky130_fd_sc_hd__buf_1
Xwire479 net480 VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__clkbuf_1
X_14191_ _06411_ VGND VGND VPWR VPWR _06451_ sky130_fd_sc_hd__inv_2
X_23389_ _03256_ _03258_ VGND VGND VPWR VPWR _03259_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25128_ clknet_leaf_51_clk _00017_ net8809 VGND VGND VPWR VPWR svm0.tC\[0\] sky130_fd_sc_hd__dfrtp_1
X_13142_ _05413_ _05414_ VGND VGND VPWR VPWR _05415_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13073_ _05345_ VGND VGND VPWR VPWR _05346_ sky130_fd_sc_hd__buf_1
X_25059_ net1628 _04807_ net2147 VGND VGND VPWR VPWR _04808_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17950_ net7022 _09800_ _09637_ VGND VGND VPWR VPWR _09801_ sky130_fd_sc_hd__a21oi_1
Xwire3030 _04857_ VGND VGND VPWR VPWR net3030 sky130_fd_sc_hd__buf_1
XFILLER_0_104_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3041 _03971_ VGND VGND VPWR VPWR net3041 sky130_fd_sc_hd__clkbuf_2
X_16901_ net6372 VGND VGND VPWR VPWR _08865_ sky130_fd_sc_hd__inv_2
Xwire3052 net3053 VGND VGND VPWR VPWR net3052 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_168_Right_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire3063 _02867_ VGND VGND VPWR VPWR net3063 sky130_fd_sc_hd__buf_1
XFILLER_0_40_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17881_ net3245 _09731_ VGND VGND VPWR VPWR _09732_ sky130_fd_sc_hd__xnor2_1
Xwire3074 net3075 VGND VGND VPWR VPWR net3074 sky130_fd_sc_hd__clkbuf_1
Xwire2340 _04930_ VGND VGND VPWR VPWR net2340 sky130_fd_sc_hd__clkbuf_1
Xwire3085 _02599_ VGND VGND VPWR VPWR net3085 sky130_fd_sc_hd__buf_1
Xwire2351 net2352 VGND VGND VPWR VPWR net2351 sky130_fd_sc_hd__buf_1
X_19620_ _11454_ _11456_ VGND VGND VPWR VPWR _11457_ sky130_fd_sc_hd__xnor2_1
Xwire3096 net3097 VGND VGND VPWR VPWR net3096 sky130_fd_sc_hd__clkbuf_1
X_16832_ net6427 matmul0.sin\[4\] _08803_ VGND VGND VPWR VPWR _08807_ sky130_fd_sc_hd__mux2_1
Xwire2362 net2364 VGND VGND VPWR VPWR net2362 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2373 net2376 VGND VGND VPWR VPWR net2373 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2384 _00011_ VGND VGND VPWR VPWR net2384 sky130_fd_sc_hd__buf_1
Xwire1650 _04283_ VGND VGND VPWR VPWR net1650 sky130_fd_sc_hd__buf_2
Xwire2395 net2396 VGND VGND VPWR VPWR net2395 sky130_fd_sc_hd__buf_1
Xwire1661 _03631_ VGND VGND VPWR VPWR net1661 sky130_fd_sc_hd__clkbuf_1
X_19551_ _11384_ _11386_ VGND VGND VPWR VPWR _11388_ sky130_fd_sc_hd__or2_1
XFILLER_0_189_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16763_ matmul0.a_in\[1\] matmul0.a\[1\] net3378 VGND VGND VPWR VPWR _08771_ sky130_fd_sc_hd__mux2_1
Xwire1672 net1673 VGND VGND VPWR VPWR net1672 sky130_fd_sc_hd__clkbuf_1
X_13975_ _06173_ net1965 net1583 _06177_ _06239_ VGND VGND VPWR VPWR _06240_ sky130_fd_sc_hd__a41o_1
Xwire1683 net1684 VGND VGND VPWR VPWR net1683 sky130_fd_sc_hd__clkbuf_1
Xwire1694 net1695 VGND VGND VPWR VPWR net1694 sky130_fd_sc_hd__clkbuf_1
X_18502_ _10349_ _10350_ VGND VGND VPWR VPWR _10351_ sky130_fd_sc_hd__nor2_1
X_15714_ net3398 _07656_ _07784_ VGND VGND VPWR VPWR _07785_ sky130_fd_sc_hd__o21a_1
XFILLER_0_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12926_ net1140 net1004 VGND VGND VPWR VPWR _05199_ sky130_fd_sc_hd__xnor2_2
X_19482_ net6297 net6359 _10851_ VGND VGND VPWR VPWR _11319_ sky130_fd_sc_hd__or3b_1
XFILLER_0_87_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16694_ _08722_ _08718_ _08723_ VGND VGND VPWR VPWR _08724_ sky130_fd_sc_hd__a21o_1
X_18433_ _10222_ _10224_ net6827 VGND VGND VPWR VPWR _10283_ sky130_fd_sc_hd__o21ai_1
X_15645_ _07716_ VGND VGND VPWR VPWR _07717_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_180_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12857_ net7272 _04892_ net3695 net2991 net7548 VGND VGND VPWR VPWR _05130_ sky130_fd_sc_hd__a32oi_1
XFILLER_0_29_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18364_ _10208_ _10211_ _10214_ _10209_ VGND VGND VPWR VPWR _10215_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12788_ net4260 net7876 _04974_ _04975_ VGND VGND VPWR VPWR _05061_ sky130_fd_sc_hd__and4_1
X_15576_ net2830 net3488 VGND VGND VPWR VPWR _07648_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17315_ net6714 net7764 VGND VGND VPWR VPWR _09229_ sky130_fd_sc_hd__xor2_1
XFILLER_0_7_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14527_ net726 _06706_ VGND VGND VPWR VPWR _06707_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18295_ _10139_ _10142_ _10143_ _10145_ VGND VGND VPWR VPWR _10146_ sky130_fd_sc_hd__a211o_1
XFILLER_0_113_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17246_ net2165 net285 net1800 net9204 VGND VGND VPWR VPWR _00344_ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14458_ _06530_ matmul0.op_in\[0\] _06541_ net6443 net4235 VGND VGND VPWR VPWR _06648_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_25_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13409_ _05652_ _05656_ VGND VGND VPWR VPWR _05682_ sky130_fd_sc_hd__and2b_1
X_14389_ net5312 net1297 net2895 net4471 _06594_ VGND VGND VPWR VPWR _06595_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17177_ net6891 net670 _09127_ _09128_ VGND VGND VPWR VPWR _09129_ sky130_fd_sc_hd__o211a_1
Xwire980 _08269_ VGND VGND VPWR VPWR net980 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire991 _07168_ VGND VGND VPWR VPWR net991 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap735 _05245_ VGND VGND VPWR VPWR net735 sky130_fd_sc_hd__buf_1
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16128_ net3492 net2697 net3442 net3516 VGND VGND VPWR VPWR _08194_ sky130_fd_sc_hd__a211o_1
XFILLER_0_84_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16059_ _08120_ _08125_ VGND VGND VPWR VPWR _08126_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_135_Right_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19818_ net1747 _11651_ VGND VGND VPWR VPWR _11652_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_102_Left_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19749_ _11581_ _11583_ VGND VGND VPWR VPWR _11584_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_194_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22760_ pid_d.ki\[11\] net3068 net2037 VGND VGND VPWR VPWR _02685_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21711_ _01652_ _01721_ VGND VGND VPWR VPWR _01722_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_188_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22691_ _02635_ net5532 net2447 VGND VGND VPWR VPWR _02636_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24430_ net4895 net4504 _04200_ VGND VGND VPWR VPWR _04288_ sky130_fd_sc_hd__or3_1
X_21642_ net1177 _01601_ net1178 VGND VGND VPWR VPWR _01653_ sky130_fd_sc_hd__o21ba_1
Xwire8008 net8009 VGND VGND VPWR VPWR net8008 sky130_fd_sc_hd__clkbuf_1
Xwire8019 net8020 VGND VGND VPWR VPWR net8019 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24361_ net2019 net1652 VGND VGND VPWR VPWR _04220_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21573_ net5816 net5458 VGND VGND VPWR VPWR _01585_ sky130_fd_sc_hd__nand2_1
Xwire7307 net7308 VGND VGND VPWR VPWR net7307 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7318 net7319 VGND VGND VPWR VPWR net7318 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7329 net7330 VGND VGND VPWR VPWR net7329 sky130_fd_sc_hd__buf_1
X_23312_ _02946_ _02961_ _02948_ VGND VGND VPWR VPWR _03182_ sky130_fd_sc_hd__a21o_1
Xmax_length3027 _04870_ VGND VGND VPWR VPWR net3027 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20524_ net2082 net2084 VGND VGND VPWR VPWR _12310_ sky130_fd_sc_hd__or2_1
X_24292_ _04143_ _04151_ VGND VGND VPWR VPWR _04152_ sky130_fd_sc_hd__xnor2_2
Xwire6606 net6607 VGND VGND VPWR VPWR net6606 sky130_fd_sc_hd__clkbuf_1
Xwire6617 net6613 VGND VGND VPWR VPWR net6617 sky130_fd_sc_hd__buf_1
XFILLER_0_172_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire6628 net6626 VGND VGND VPWR VPWR net6628 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6639 net6640 VGND VGND VPWR VPWR net6639 sky130_fd_sc_hd__buf_1
X_23243_ _03104_ _03112_ VGND VGND VPWR VPWR _03113_ sky130_fd_sc_hd__xnor2_1
Xwire5905 net5906 VGND VGND VPWR VPWR net5905 sky130_fd_sc_hd__buf_1
XFILLER_0_133_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length1603 _05057_ VGND VGND VPWR VPWR net1603 sky130_fd_sc_hd__buf_1
Xwire5916 net5912 VGND VGND VPWR VPWR net5916 sky130_fd_sc_hd__buf_1
X_20455_ cordic0.slte0.opA\[14\] _06509_ VGND VGND VPWR VPWR _12248_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5927 pid_d.mult0.b\[2\] VGND VGND VPWR VPWR net5927 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5949 net5951 VGND VGND VPWR VPWR net5949 sky130_fd_sc_hd__buf_1
X_23174_ _03033_ _03038_ _03043_ VGND VGND VPWR VPWR _03044_ sky130_fd_sc_hd__nand3_1
X_20386_ net1054 _12169_ _12183_ VGND VGND VPWR VPWR _12185_ sky130_fd_sc_hd__and3_1
X_22125_ net5720 net5437 VGND VGND VPWR VPWR _02131_ sky130_fd_sc_hd__nand2_1
X_22056_ _01948_ _01950_ _02062_ VGND VGND VPWR VPWR _02063_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_102_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21007_ _01022_ _00963_ VGND VGND VPWR VPWR _01023_ sky130_fd_sc_hd__xnor2_1
X_25815_ clknet_leaf_37_clk _00688_ net8749 VGND VGND VPWR VPWR pid_q.prev_error\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13760_ net7741 net3670 VGND VGND VPWR VPWR _06028_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22958_ _02830_ _02844_ _02845_ VGND VGND VPWR VPWR _02846_ sky130_fd_sc_hd__a21oi_1
X_25746_ clknet_leaf_8_clk _00619_ net8554 VGND VGND VPWR VPWR pid_d.kp\[4\] sky130_fd_sc_hd__dfrtp_1
X_12711_ _04980_ _04981_ _04983_ VGND VGND VPWR VPWR _04984_ sky130_fd_sc_hd__o21ai_4
X_21909_ net5978 VGND VGND VPWR VPWR _01917_ sky130_fd_sc_hd__inv_2
X_13691_ _05957_ net782 VGND VGND VPWR VPWR _05960_ sky130_fd_sc_hd__xor2_1
X_25677_ clknet_leaf_4_clk _00550_ net8563 VGND VGND VPWR VPWR pid_d.prev_error\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_22889_ net8895 _02783_ VGND VGND VPWR VPWR _02784_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8414 net8537 VGND VGND VPWR VPWR net8414 sky130_fd_sc_hd__buf_1
X_12642_ _04908_ _04914_ VGND VGND VPWR VPWR _04915_ sky130_fd_sc_hd__xnor2_1
X_15430_ _07398_ _07400_ _07503_ VGND VGND VPWR VPWR _07504_ sky130_fd_sc_hd__a21o_1
X_24628_ net4514 _04482_ _04478_ _04475_ VGND VGND VPWR VPWR _04483_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout7724 svm0.periodTop\[9\] VGND VGND VPWR VPWR net7724 sky130_fd_sc_hd__buf_1
X_15361_ _07412_ _07415_ _07431_ _07433_ _07434_ VGND VGND VPWR VPWR _07435_ sky130_fd_sc_hd__o311a_1
Xwire8520 net8523 VGND VGND VPWR VPWR net8520 sky130_fd_sc_hd__clkbuf_1
X_24559_ net4809 VGND VGND VPWR VPWR _04415_ sky130_fd_sc_hd__inv_2
X_12573_ net7478 net8863 VGND VGND VPWR VPWR _04862_ sky130_fd_sc_hd__or2b_1
Xwire8531 net8532 VGND VGND VPWR VPWR net8531 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_66_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8542 net8543 VGND VGND VPWR VPWR net8542 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8553 net8551 VGND VGND VPWR VPWR net8553 sky130_fd_sc_hd__clkbuf_2
Xmax_length4240 net4241 VGND VGND VPWR VPWR net4240 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17100_ _09053_ net3326 _09056_ net2602 _08955_ VGND VGND VPWR VPWR _09057_ sky130_fd_sc_hd__o221a_1
Xwire7830 net7833 VGND VGND VPWR VPWR net7830 sky130_fd_sc_hd__clkbuf_1
X_14312_ net6451 net6456 net8319 VGND VGND VPWR VPWR _06534_ sky130_fd_sc_hd__or3_1
Xwire210 net211 VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_1
Xwire221 net222 VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__buf_1
X_15292_ _07343_ _07344_ _07365_ VGND VGND VPWR VPWR _07366_ sky130_fd_sc_hd__and3_1
X_18080_ net3306 _09711_ VGND VGND VPWR VPWR _09931_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire7841 net7842 VGND VGND VPWR VPWR net7841 sky130_fd_sc_hd__clkbuf_1
Xwire8586 net8587 VGND VGND VPWR VPWR net8586 sky130_fd_sc_hd__buf_1
Xwire232 net233 VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8597 net8598 VGND VGND VPWR VPWR net8597 sky130_fd_sc_hd__clkbuf_1
Xwire7852 net7853 VGND VGND VPWR VPWR net7852 sky130_fd_sc_hd__clkbuf_1
Xwire243 _12014_ VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__buf_1
Xwire254 _06361_ VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__buf_1
Xwire7863 net7864 VGND VGND VPWR VPWR net7863 sky130_fd_sc_hd__clkbuf_1
X_14243_ net152 _06496_ _06498_ VGND VGND VPWR VPWR _00033_ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17031_ net1480 VGND VGND VPWR VPWR _08991_ sky130_fd_sc_hd__buf_1
Xwire7885 net7886 VGND VGND VPWR VPWR net7885 sky130_fd_sc_hd__buf_1
Xwire276 net277 VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__clkbuf_1
Xwire287 net288 VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__buf_1
Xwire7896 net7897 VGND VGND VPWR VPWR net7896 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire298 net299 VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length2860 net2861 VGND VGND VPWR VPWR net2860 sky130_fd_sc_hd__buf_1
X_14174_ _06432_ _06433_ _06394_ VGND VGND VPWR VPWR _06434_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length2882 net2883 VGND VGND VPWR VPWR net2882 sky130_fd_sc_hd__buf_1
XFILLER_0_22_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13125_ _05364_ _05365_ net734 VGND VGND VPWR VPWR _05398_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_131_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18982_ net2530 _10818_ VGND VGND VPWR VPWR _10819_ sky130_fd_sc_hd__xnor2_2
X_13056_ net790 _05208_ VGND VGND VPWR VPWR _05329_ sky130_fd_sc_hd__nand2_1
X_17933_ net2561 net2559 VGND VGND VPWR VPWR _09784_ sky130_fd_sc_hd__nand2_1
X_17864_ _08985_ net3258 _09707_ VGND VGND VPWR VPWR _09715_ sky130_fd_sc_hd__o21a_1
XFILLER_0_139_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2170 _09070_ VGND VGND VPWR VPWR net2170 sky130_fd_sc_hd__clkbuf_1
X_19603_ net6012 _11439_ VGND VGND VPWR VPWR _11440_ sky130_fd_sc_hd__nand2_1
Xwire2181 net2188 VGND VGND VPWR VPWR net2181 sky130_fd_sc_hd__buf_1
X_16815_ cordic0.cos\[10\] matmul0.cos\[10\] net3368 VGND VGND VPWR VPWR _08798_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2192 net2193 VGND VGND VPWR VPWR net2192 sky130_fd_sc_hd__buf_1
XFILLER_0_108_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17795_ _09644_ _09645_ net7082 VGND VGND VPWR VPWR _09646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1480 net1481 VGND VGND VPWR VPWR net1480 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1491 net1493 VGND VGND VPWR VPWR net1491 sky130_fd_sc_hd__buf_1
X_19534_ _11306_ _11300_ VGND VGND VPWR VPWR _11371_ sky130_fd_sc_hd__and2b_1
X_16746_ net7566 matmul0.b\[9\] net3380 VGND VGND VPWR VPWR _08762_ sky130_fd_sc_hd__mux2_1
X_13958_ _06220_ _06222_ VGND VGND VPWR VPWR _06223_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_177_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12909_ _05176_ _05181_ VGND VGND VPWR VPWR _05182_ sky130_fd_sc_hd__xor2_1
X_19465_ _11254_ _11300_ VGND VGND VPWR VPWR _11302_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16677_ _08709_ VGND VGND VPWR VPWR _00256_ sky130_fd_sc_hd__clkbuf_1
X_13889_ _06080_ _06142_ _06154_ VGND VGND VPWR VPWR _06155_ sky130_fd_sc_hd__a21oi_1
X_18416_ net716 net715 _10257_ _10265_ VGND VGND VPWR VPWR _10266_ sky130_fd_sc_hd__or4_1
X_15628_ _07698_ _07699_ VGND VGND VPWR VPWR _07700_ sky130_fd_sc_hd__xor2_1
XFILLER_0_173_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19396_ _11231_ _11232_ VGND VGND VPWR VPWR _11233_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18347_ _10192_ _10194_ _10197_ VGND VGND VPWR VPWR _10198_ sky130_fd_sc_hd__a21o_1
X_15559_ _07541_ _07502_ _07504_ VGND VGND VPWR VPWR _07632_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_86_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18278_ net1074 _10127_ _10128_ VGND VGND VPWR VPWR _10129_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput40 currB_in[1] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
X_17229_ _09176_ VGND VGND VPWR VPWR _09177_ sky130_fd_sc_hd__buf_1
XFILLER_0_3_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput51 currT_in[11] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput62 currT_in[7] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput73 periodTop[2] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput84 pid_d_addr[12] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_1
X_20240_ _12056_ cordic0.slte0.opB\[8\] net2936 VGND VGND VPWR VPWR _12057_ sky130_fd_sc_hd__mux2_1
Xinput95 pid_d_addr[8] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20171_ net6004 net3137 _11754_ _11996_ net6072 VGND VGND VPWR VPWR _11997_ sky130_fd_sc_hd__a32o_1
XFILLER_0_161_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_110_Left_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23930_ _03788_ _03793_ VGND VGND VPWR VPWR _03794_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_165_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23861_ _03595_ _03597_ _03725_ VGND VGND VPWR VPWR _03726_ sky130_fd_sc_hd__o21ai_1
Xmax_length8517 net8510 VGND VGND VPWR VPWR net8517 sky130_fd_sc_hd__buf_1
XFILLER_0_165_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25600_ clknet_leaf_105_clk _00473_ net8358 VGND VGND VPWR VPWR cordic0.slte0.opB\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_22812_ net4299 net2464 VGND VGND VPWR VPWR _02715_ sky130_fd_sc_hd__nor2_1
XFILLER_0_196_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23792_ net744 _03559_ _03657_ VGND VGND VPWR VPWR _03658_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_189_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25531_ clknet_leaf_35_clk _00411_ net8764 VGND VGND VPWR VPWR svm0.state\[1\] sky130_fd_sc_hd__dfrtp_2
X_22743_ _02673_ VGND VGND VPWR VPWR _00604_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_177_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25462_ clknet_leaf_53_clk _00342_ net8804 VGND VGND VPWR VPWR svm0.tB\[0\] sky130_fd_sc_hd__dfrtp_1
X_22674_ net3705 VGND VGND VPWR VPWR _02624_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24413_ net2019 net1652 _04213_ VGND VGND VPWR VPWR _04271_ sky130_fd_sc_hd__o21a_1
XFILLER_0_191_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21625_ _01636_ _01535_ pid_d.prev_error\[3\] VGND VGND VPWR VPWR _01637_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_30_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25393_ clknet_leaf_80_clk _00276_ net8497 VGND VGND VPWR VPWR matmul0.b\[12\] sky130_fd_sc_hd__dfrtp_1
Xwire7115 net7116 VGND VGND VPWR VPWR net7115 sky130_fd_sc_hd__buf_1
X_24344_ _04201_ _04202_ VGND VGND VPWR VPWR _04203_ sky130_fd_sc_hd__xnor2_1
Xwire7126 net7128 VGND VGND VPWR VPWR net7126 sky130_fd_sc_hd__buf_1
XFILLER_0_74_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21556_ _01556_ _01567_ VGND VGND VPWR VPWR _01568_ sky130_fd_sc_hd__xnor2_1
Xwire7137 net7134 VGND VGND VPWR VPWR net7137 sky130_fd_sc_hd__buf_1
XFILLER_0_62_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6403 cordic0.slte0.opB\[10\] VGND VGND VPWR VPWR net6403 sky130_fd_sc_hd__clkbuf_1
Xwire7148 matmul0.sin\[13\] VGND VGND VPWR VPWR net7148 sky130_fd_sc_hd__clkbuf_2
Xwire6414 net6415 VGND VGND VPWR VPWR net6414 sky130_fd_sc_hd__clkbuf_1
Xwire7159 matmul0.sin\[2\] VGND VGND VPWR VPWR net7159 sky130_fd_sc_hd__buf_1
XFILLER_0_7_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6425 net6426 VGND VGND VPWR VPWR net6425 sky130_fd_sc_hd__clkbuf_1
X_20507_ net6461 _12268_ net2492 _12293_ VGND VGND VPWR VPWR _12294_ sky130_fd_sc_hd__o31a_1
X_24275_ _04131_ _04134_ VGND VGND VPWR VPWR _04135_ sky130_fd_sc_hd__xnor2_2
Xwire6436 net6437 VGND VGND VPWR VPWR net6436 sky130_fd_sc_hd__clkbuf_1
Xwire5702 net5705 VGND VGND VPWR VPWR net5702 sky130_fd_sc_hd__buf_1
X_21487_ net1725 _01499_ VGND VGND VPWR VPWR _01500_ sky130_fd_sc_hd__xnor2_1
Xwire5713 net5714 VGND VGND VPWR VPWR net5713 sky130_fd_sc_hd__clkbuf_1
Xwire6458 net6459 VGND VGND VPWR VPWR net6458 sky130_fd_sc_hd__buf_1
X_23226_ _03094_ _03095_ VGND VGND VPWR VPWR _03096_ sky130_fd_sc_hd__xnor2_1
Xwire5735 net5736 VGND VGND VPWR VPWR net5735 sky130_fd_sc_hd__buf_1
X_20438_ net6493 net2166 VGND VGND VPWR VPWR _12232_ sky130_fd_sc_hd__nand2_1
Xwire5746 net5749 VGND VGND VPWR VPWR net5746 sky130_fd_sc_hd__buf_1
Xwire5757 net5751 VGND VGND VPWR VPWR net5757 sky130_fd_sc_hd__clkbuf_1
Xwire5768 net5769 VGND VGND VPWR VPWR net5768 sky130_fd_sc_hd__buf_1
Xwire5779 net5780 VGND VGND VPWR VPWR net5779 sky130_fd_sc_hd__buf_1
X_23157_ net4983 net4776 VGND VGND VPWR VPWR _03027_ sky130_fd_sc_hd__nand2_1
X_20369_ cordic0.slte0.opA\[7\] _12168_ VGND VGND VPWR VPWR _12169_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22108_ net471 _02003_ _02004_ _02097_ VGND VGND VPWR VPWR _02114_ sky130_fd_sc_hd__a211o_1
X_23088_ _02890_ _02891_ VGND VGND VPWR VPWR _02958_ sky130_fd_sc_hd__nor2_1
X_22039_ _01942_ _01943_ _01944_ VGND VGND VPWR VPWR _02046_ sky130_fd_sc_hd__o21a_1
X_14930_ net4171 net4167 net4196 net4194 VGND VGND VPWR VPWR _07004_ sky130_fd_sc_hd__o22a_1
XFILLER_0_54_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14861_ net7187 matmul0.matmul_stage_inst.f\[3\] net3609 VGND VGND VPWR VPWR _06948_
+ sky130_fd_sc_hd__mux2_1
X_16600_ matmul0.matmul_stage_inst.mult2\[7\] net354 net2616 VGND VGND VPWR VPWR _08650_
+ sky130_fd_sc_hd__mux2_1
X_13812_ net531 net678 VGND VGND VPWR VPWR _06080_ sky130_fd_sc_hd__or2_1
X_17580_ net6712 _09461_ svm0.tC\[8\] VGND VGND VPWR VPWR _09462_ sky130_fd_sc_hd__o21ba_1
X_14792_ net9007 net2871 _06912_ VGND VGND VPWR VPWR _00168_ sky130_fd_sc_hd__a21o_1
XFILLER_0_159_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16531_ _08589_ _08590_ VGND VGND VPWR VPWR _08591_ sky130_fd_sc_hd__or2b_1
XFILLER_0_97_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13743_ net9147 net1126 net223 net1926 VGND VGND VPWR VPWR _00020_ sky130_fd_sc_hd__a22o_1
X_25729_ clknet_leaf_8_clk _00602_ net8553 VGND VGND VPWR VPWR pid_d.ki\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_196_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19250_ _11085_ _11086_ VGND VGND VPWR VPWR _11087_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16462_ _08447_ _08464_ _08522_ VGND VGND VPWR VPWR _08523_ sky130_fd_sc_hd__o21a_1
X_13674_ net7770 net1306 _05875_ _05876_ VGND VGND VPWR VPWR _05943_ sky130_fd_sc_hd__a22o_1
X_18201_ _10049_ _10050_ net2547 VGND VGND VPWR VPWR _10052_ sky130_fd_sc_hd__a21o_1
X_15413_ net2778 net3428 net3426 net2781 VGND VGND VPWR VPWR _07487_ sky130_fd_sc_hd__o211a_1
X_12625_ net6749 net6599 net5268 VGND VGND VPWR VPWR _04898_ sky130_fd_sc_hd__and3_1
Xfanout7521 pid_q.state\[1\] VGND VGND VPWR VPWR net7521 sky130_fd_sc_hd__buf_1
X_19181_ net3187 _10922_ _11013_ _11016_ _11017_ VGND VGND VPWR VPWR _11018_ sky130_fd_sc_hd__a32o_1
XFILLER_0_6_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16393_ net2750 _08454_ VGND VGND VPWR VPWR _08455_ sky130_fd_sc_hd__nor2_1
XFILLER_0_182_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8350 net8351 VGND VGND VPWR VPWR net8350 sky130_fd_sc_hd__buf_1
X_18132_ _09916_ _09921_ _09982_ VGND VGND VPWR VPWR _09983_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_170_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8361 net8359 VGND VGND VPWR VPWR net8361 sky130_fd_sc_hd__dlymetal6s2s_1
X_15344_ _07416_ _07417_ VGND VGND VPWR VPWR _07418_ sky130_fd_sc_hd__nand2_1
Xwire8372 net8373 VGND VGND VPWR VPWR net8372 sky130_fd_sc_hd__clkbuf_1
Xfanout6831 net6834 VGND VGND VPWR VPWR net6831 sky130_fd_sc_hd__buf_1
XFILLER_0_54_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18063_ _09905_ _09913_ VGND VGND VPWR VPWR _09914_ sky130_fd_sc_hd__xor2_2
XFILLER_0_41_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire7671 net7673 VGND VGND VPWR VPWR net7671 sky130_fd_sc_hd__buf_1
X_15275_ _07345_ _07348_ VGND VGND VPWR VPWR _07349_ sky130_fd_sc_hd__xnor2_1
Xwire7682 net7683 VGND VGND VPWR VPWR net7682 sky130_fd_sc_hd__buf_1
Xwire7693 net7694 VGND VGND VPWR VPWR net7693 sky130_fd_sc_hd__clkbuf_1
X_17014_ net2173 net1806 VGND VGND VPWR VPWR _08975_ sky130_fd_sc_hd__or2_1
Xhold109 cordic0.sin\[10\] VGND VGND VPWR VPWR net9062 sky130_fd_sc_hd__dlygate4sd3_1
X_14226_ net1119 _06470_ _06483_ VGND VGND VPWR VPWR _06484_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6992 net6985 VGND VGND VPWR VPWR net6992 sky130_fd_sc_hd__buf_1
XFILLER_0_1_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14157_ _06411_ _06417_ VGND VGND VPWR VPWR _06418_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13108_ _05255_ _05260_ VGND VGND VPWR VPWR _05381_ sky130_fd_sc_hd__nor2_1
X_14088_ _06349_ _06350_ VGND VGND VPWR VPWR _06351_ sky130_fd_sc_hd__nand2_1
X_18965_ net6232 net6264 VGND VGND VPWR VPWR _10802_ sky130_fd_sc_hd__or2b_1
XFILLER_0_185_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13039_ net791 net736 _05126_ VGND VGND VPWR VPWR _05312_ sky130_fd_sc_hd__a21o_1
X_17916_ _09762_ _09764_ _09766_ _09666_ VGND VGND VPWR VPWR _09767_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18896_ net6794 _10714_ _10736_ net6860 VGND VGND VPWR VPWR _10737_ sky130_fd_sc_hd__a22o_1
X_17847_ _09693_ _09695_ _09697_ VGND VGND VPWR VPWR _09698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_179_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17778_ _09612_ net1448 VGND VGND VPWR VPWR _09629_ sky130_fd_sc_hd__xnor2_2
X_19517_ net2522 _11295_ _11296_ VGND VGND VPWR VPWR _11354_ sky130_fd_sc_hd__o21ai_1
X_16729_ net7574 matmul0.b\[1\] net3702 VGND VGND VPWR VPWR _08753_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19448_ _11282_ _11283_ _11261_ VGND VGND VPWR VPWR _11285_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_158_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19379_ _11210_ _11212_ VGND VGND VPWR VPWR _11216_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21410_ _01420_ net757 VGND VGND VPWR VPWR _01424_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22390_ _02262_ _02391_ _02392_ VGND VGND VPWR VPWR _02393_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21341_ net5654 _01354_ _01349_ VGND VGND VPWR VPWR _01355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5009 net5010 VGND VGND VPWR VPWR net5009 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24060_ _03795_ _03800_ _03801_ VGND VGND VPWR VPWR _03923_ sky130_fd_sc_hd__o21a_1
X_21272_ _01284_ _01286_ VGND VGND VPWR VPWR _01287_ sky130_fd_sc_hd__xor2_1
Xwire4308 _04866_ VGND VGND VPWR VPWR net4308 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4319 net4318 VGND VGND VPWR VPWR net4319 sky130_fd_sc_hd__buf_1
X_23011_ net5087 net4623 VGND VGND VPWR VPWR _02881_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20223_ net8953 net8119 net8 net8100 VGND VGND VPWR VPWR _12043_ sky130_fd_sc_hd__and4_1
XFILLER_0_40_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3607 net3608 VGND VGND VPWR VPWR net3607 sky130_fd_sc_hd__clkbuf_2
Xwire3618 net3619 VGND VGND VPWR VPWR net3618 sky130_fd_sc_hd__buf_1
Xwire3629 _06800_ VGND VGND VPWR VPWR net3629 sky130_fd_sc_hd__buf_1
Xwire2906 net2907 VGND VGND VPWR VPWR net2906 sky130_fd_sc_hd__clkbuf_1
X_20154_ _11911_ _11920_ VGND VGND VPWR VPWR _11981_ sky130_fd_sc_hd__or2_1
Xwire2917 net2918 VGND VGND VPWR VPWR net2917 sky130_fd_sc_hd__clkbuf_1
Xwire2928 net2929 VGND VGND VPWR VPWR net2928 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2939 net2940 VGND VGND VPWR VPWR net2939 sky130_fd_sc_hd__clkbuf_1
X_24962_ pid_q.kp\[0\] _04694_ _04735_ VGND VGND VPWR VPWR _04736_ sky130_fd_sc_hd__mux2_1
X_20085_ net350 _11839_ VGND VGND VPWR VPWR _11914_ sky130_fd_sc_hd__nand2_1
X_23913_ _03656_ _03677_ _03676_ VGND VGND VPWR VPWR _03777_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24893_ _04686_ pid_q.mult0.a\[12\] net1998 VGND VGND VPWR VPWR _04687_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23844_ net4688 net4827 VGND VGND VPWR VPWR _03709_ sky130_fd_sc_hd__nand2_1
Xmax_length8347 net8343 VGND VGND VPWR VPWR net8347 sky130_fd_sc_hd__buf_1
XFILLER_0_196_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length7635 net7636 VGND VGND VPWR VPWR net7635 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_178_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23775_ net1019 net1018 _03640_ VGND VGND VPWR VPWR _03641_ sky130_fd_sc_hd__o21a_1
XFILLER_0_192_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20987_ _00998_ _01002_ VGND VGND VPWR VPWR _01003_ sky130_fd_sc_hd__xnor2_1
X_25514_ clknet_leaf_43_clk _00394_ net8783 VGND VGND VPWR VPWR svm0.counter\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_22726_ net2037 VGND VGND VPWR VPWR _02662_ sky130_fd_sc_hd__clkbuf_1
Xmax_length6967 net6968 VGND VGND VPWR VPWR net6967 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_177_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6978 net6973 VGND VGND VPWR VPWR net6978 sky130_fd_sc_hd__buf_1
X_22657_ net9156 _02599_ _02613_ net337 net8890 VGND VGND VPWR VPWR _00578_ sky130_fd_sc_hd__o221a_1
X_25445_ clknet_leaf_117_clk _00328_ net8332 VGND VGND VPWR VPWR cordic0.vec\[1\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21608_ net5416 net5893 _01513_ VGND VGND VPWR VPWR _01620_ sky130_fd_sc_hd__a21oi_1
X_13390_ _05401_ _05662_ VGND VGND VPWR VPWR _05663_ sky130_fd_sc_hd__xor2_1
XFILLER_0_168_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25376_ clknet_leaf_58_clk _00259_ net8726 VGND VGND VPWR VPWR matmul0.alpha_pass\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout6127 net6135 VGND VGND VPWR VPWR net6127 sky130_fd_sc_hd__buf_1
XFILLER_0_8_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22588_ net7294 _02564_ VGND VGND VPWR VPWR _02566_ sky130_fd_sc_hd__or2_1
Xfanout6138 net6147 VGND VGND VPWR VPWR net6138 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24327_ _02869_ _04118_ _04186_ VGND VGND VPWR VPWR _00675_ sky130_fd_sc_hd__o21a_1
Xwire6222 net6220 VGND VGND VPWR VPWR net6222 sky130_fd_sc_hd__buf_1
X_21539_ net702 _01546_ VGND VGND VPWR VPWR _01551_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6244 net6246 VGND VGND VPWR VPWR net6244 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire5510 net5511 VGND VGND VPWR VPWR net5510 sky130_fd_sc_hd__buf_1
Xfanout5459 pid_d.mult0.a\[11\] VGND VGND VPWR VPWR net5459 sky130_fd_sc_hd__clkbuf_1
Xwire6255 net6253 VGND VGND VPWR VPWR net6255 sky130_fd_sc_hd__buf_1
X_15060_ _07133_ VGND VGND VPWR VPWR _07134_ sky130_fd_sc_hd__buf_1
XFILLER_0_160_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5521 net5522 VGND VGND VPWR VPWR net5521 sky130_fd_sc_hd__clkbuf_1
X_24258_ _04117_ _02868_ VGND VGND VPWR VPWR _04118_ sky130_fd_sc_hd__nor2_1
Xwire6266 net6267 VGND VGND VPWR VPWR net6266 sky130_fd_sc_hd__buf_1
Xwire6277 net6278 VGND VGND VPWR VPWR net6277 sky130_fd_sc_hd__buf_1
XFILLER_0_49_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6288 net6289 VGND VGND VPWR VPWR net6288 sky130_fd_sc_hd__buf_1
Xwire5543 net5544 VGND VGND VPWR VPWR net5543 sky130_fd_sc_hd__buf_1
X_14011_ _05862_ net321 net320 _06274_ VGND VGND VPWR VPWR _06275_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_120_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5554 net5555 VGND VGND VPWR VPWR net5554 sky130_fd_sc_hd__clkbuf_1
X_23209_ net5104 net4736 VGND VGND VPWR VPWR _03079_ sky130_fd_sc_hd__nor2_1
Xwire4820 net4814 VGND VGND VPWR VPWR net4820 sky130_fd_sc_hd__clkbuf_1
Xwire6299 net6300 VGND VGND VPWR VPWR net6299 sky130_fd_sc_hd__buf_1
Xmax_length1252 net1253 VGND VGND VPWR VPWR net1252 sky130_fd_sc_hd__buf_1
XFILLER_0_120_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5565 net5566 VGND VGND VPWR VPWR net5565 sky130_fd_sc_hd__buf_1
Xwire4831 net4832 VGND VGND VPWR VPWR net4831 sky130_fd_sc_hd__clkbuf_1
X_24189_ _04003_ _04014_ _04049_ VGND VGND VPWR VPWR _04050_ sky130_fd_sc_hd__o21ai_1
Xwire5576 net5577 VGND VGND VPWR VPWR net5576 sky130_fd_sc_hd__clkbuf_1
Xwire4842 net4843 VGND VGND VPWR VPWR net4842 sky130_fd_sc_hd__buf_1
Xwire5587 net5588 VGND VGND VPWR VPWR net5587 sky130_fd_sc_hd__clkbuf_1
Xwire4853 net4857 VGND VGND VPWR VPWR net4853 sky130_fd_sc_hd__buf_1
Xwire5598 net5599 VGND VGND VPWR VPWR net5598 sky130_fd_sc_hd__buf_1
Xwire4875 net4876 VGND VGND VPWR VPWR net4875 sky130_fd_sc_hd__buf_1
XFILLER_0_105_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4886 net4887 VGND VGND VPWR VPWR net4886 sky130_fd_sc_hd__clkbuf_1
X_18750_ _10572_ _10594_ VGND VGND VPWR VPWR _10595_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_179_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15962_ _08026_ _08029_ VGND VGND VPWR VPWR _08030_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_175_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17701_ _09576_ VGND VGND VPWR VPWR _09577_ sky130_fd_sc_hd__buf_1
X_14913_ net4222 net4220 VGND VGND VPWR VPWR _06987_ sky130_fd_sc_hd__or2_1
X_18681_ net3296 _10525_ _10526_ _10475_ VGND VGND VPWR VPWR _10527_ sky130_fd_sc_hd__or4b_1
X_15893_ net987 _07857_ _07858_ VGND VGND VPWR VPWR _07962_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_175_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17632_ net6699 _09512_ svm0.tB\[12\] VGND VGND VPWR VPWR _09513_ sky130_fd_sc_hd__o21ba_1
X_14844_ net4283 VGND VGND VPWR VPWR _06939_ sky130_fd_sc_hd__buf_1
XFILLER_0_172_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17563_ net6712 svm0.tC\[8\] VGND VGND VPWR VPWR _09445_ sky130_fd_sc_hd__xnor2_1
X_14775_ matmul0.sin\[11\] _06900_ VGND VGND VPWR VPWR _06901_ sky130_fd_sc_hd__xor2_1
XFILLER_0_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19302_ _11134_ _11135_ _11138_ VGND VGND VPWR VPWR _11139_ sky130_fd_sc_hd__mux2_1
X_16514_ net2665 _08511_ _08573_ VGND VGND VPWR VPWR _08574_ sky130_fd_sc_hd__a21o_1
X_13726_ _05921_ _05924_ _05925_ VGND VGND VPWR VPWR _05995_ sky130_fd_sc_hd__o21ba_1
X_17494_ _09303_ net770 _09382_ VGND VGND VPWR VPWR _09383_ sky130_fd_sc_hd__a21o_1
XFILLER_0_112_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19233_ net1422 _11069_ VGND VGND VPWR VPWR _11070_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8041 net8046 VGND VGND VPWR VPWR net8041 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16445_ net2772 net2621 net2204 VGND VGND VPWR VPWR _08506_ sky130_fd_sc_hd__or3_1
X_13657_ _05921_ _05926_ VGND VGND VPWR VPWR _05927_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_13_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19164_ net6119 net6155 net6069 _10997_ _10998_ VGND VGND VPWR VPWR _11001_ sky130_fd_sc_hd__a311o_1
X_12608_ net4279 VGND VGND VPWR VPWR _04884_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16376_ net1081 _08436_ _08437_ VGND VGND VPWR VPWR _08438_ sky130_fd_sc_hd__o21ba_1
X_13588_ net504 VGND VGND VPWR VPWR _05858_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8180 net8181 VGND VGND VPWR VPWR net8180 sky130_fd_sc_hd__clkbuf_1
X_18115_ _09965_ _09860_ net2550 _09878_ VGND VGND VPWR VPWR _09966_ sky130_fd_sc_hd__o31ai_1
Xwire8191 net8192 VGND VGND VPWR VPWR net8191 sky130_fd_sc_hd__clkbuf_1
X_15327_ _07398_ _07400_ VGND VGND VPWR VPWR _07401_ sky130_fd_sc_hd__xor2_2
X_19095_ net3208 _10929_ _10931_ net3202 VGND VGND VPWR VPWR _10932_ sky130_fd_sc_hd__o22a_1
XFILLER_0_170_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6672 net6674 VGND VGND VPWR VPWR net6672 sky130_fd_sc_hd__buf_1
XFILLER_0_2_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7490 net7491 VGND VGND VPWR VPWR net7490 sky130_fd_sc_hd__buf_1
X_18046_ _09887_ _09893_ _09896_ VGND VGND VPWR VPWR _09897_ sky130_fd_sc_hd__a21o_1
X_15258_ _07331_ _07295_ _07278_ VGND VGND VPWR VPWR _07332_ sky130_fd_sc_hd__mux2_1
X_14209_ _06439_ _06442_ VGND VGND VPWR VPWR _06468_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15189_ _07215_ _07216_ VGND VGND VPWR VPWR _07263_ sky130_fd_sc_hd__and2b_1
X_19997_ _11826_ _11827_ _11783_ net3127 VGND VGND VPWR VPWR _11828_ sky130_fd_sc_hd__o211ai_1
X_18948_ _10784_ _10785_ net2133 VGND VGND VPWR VPWR _10786_ sky130_fd_sc_hd__o21a_1
XFILLER_0_146_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18879_ _10713_ _10720_ VGND VGND VPWR VPWR _10721_ sky130_fd_sc_hd__xnor2_1
X_20910_ _00916_ _00925_ VGND VGND VPWR VPWR _00926_ sky130_fd_sc_hd__xnor2_1
X_21890_ _01896_ _01898_ VGND VGND VPWR VPWR _01899_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20841_ net3842 _00856_ VGND VGND VPWR VPWR _00857_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23560_ net4641 net4944 VGND VGND VPWR VPWR _03428_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20772_ net5578 net5794 VGND VGND VPWR VPWR _12543_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22511_ _02509_ _02511_ VGND VGND VPWR VPWR _02512_ sky130_fd_sc_hd__xnor2_1
X_23491_ _03358_ _03359_ VGND VGND VPWR VPWR _03360_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_175_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22442_ net3829 net2470 VGND VGND VPWR VPWR _02444_ sky130_fd_sc_hd__or2_1
X_25230_ clknet_leaf_65_clk _00119_ net8655 VGND VGND VPWR VPWR cordic0.in_valid sky130_fd_sc_hd__dfrtp_1
Xwire809 net810 VGND VGND VPWR VPWR net809 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length407 net408 VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__clkbuf_1
X_25161_ clknet_leaf_45_clk _00050_ net8785 VGND VGND VPWR VPWR pid_q.target\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_22373_ net2476 _02375_ VGND VGND VPWR VPWR _02376_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_190_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24112_ net3040 _03973_ VGND VGND VPWR VPWR _03974_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21324_ pid_d.curr_int\[0\] pid_d.prev_int\[0\] pid_d.prev_int\[1\] net5984 VGND
+ VGND VPWR VPWR _01338_ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25092_ net5171 VGND VGND VPWR VPWR _04836_ sky130_fd_sc_hd__inv_2
Xwire4105 net4106 VGND VGND VPWR VPWR net4105 sky130_fd_sc_hd__buf_1
X_24043_ _03899_ _03905_ VGND VGND VPWR VPWR _03906_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4116 net4117 VGND VGND VPWR VPWR net4116 sky130_fd_sc_hd__buf_1
Xwire4127 _07036_ VGND VGND VPWR VPWR net4127 sky130_fd_sc_hd__buf_1
X_21255_ _01261_ _01269_ VGND VGND VPWR VPWR _01270_ sky130_fd_sc_hd__xnor2_2
Xwire4138 _07029_ VGND VGND VPWR VPWR net4138 sky130_fd_sc_hd__buf_1
Xwire3404 net3406 VGND VGND VPWR VPWR net3404 sky130_fd_sc_hd__buf_1
Xwire4149 net4150 VGND VGND VPWR VPWR net4149 sky130_fd_sc_hd__buf_1
X_20206_ net1785 _12030_ VGND VGND VPWR VPWR _12031_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3426 _07486_ VGND VGND VPWR VPWR net3426 sky130_fd_sc_hd__buf_1
X_21186_ _01167_ _01187_ _01197_ _01201_ VGND VGND VPWR VPWR _01202_ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3437 net3438 VGND VGND VPWR VPWR net3437 sky130_fd_sc_hd__buf_1
Xwire2703 _07354_ VGND VGND VPWR VPWR net2703 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2714 _07305_ VGND VGND VPWR VPWR net2714 sky130_fd_sc_hd__buf_1
Xwire2725 _07268_ VGND VGND VPWR VPWR net2725 sky130_fd_sc_hd__buf_1
X_20137_ net274 _11964_ VGND VGND VPWR VPWR _11965_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2736 _07240_ VGND VGND VPWR VPWR net2736 sky130_fd_sc_hd__clkbuf_1
Xwire2747 net2748 VGND VGND VPWR VPWR net2747 sky130_fd_sc_hd__buf_1
Xwire2758 net2759 VGND VGND VPWR VPWR net2758 sky130_fd_sc_hd__buf_1
Xwire2769 net2770 VGND VGND VPWR VPWR net2769 sky130_fd_sc_hd__clkbuf_1
X_24945_ net8866 net132 VGND VGND VPWR VPWR _04724_ sky130_fd_sc_hd__and2b_1
X_20068_ _11887_ _11896_ VGND VGND VPWR VPWR _11897_ sky130_fd_sc_hd__xor2_2
X_24876_ _04675_ VGND VGND VPWR VPWR _00735_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12890_ net7804 net1610 _05091_ VGND VGND VPWR VPWR _05163_ sky130_fd_sc_hd__a21oi_2
X_23827_ _03688_ _03691_ VGND VGND VPWR VPWR _03692_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14560_ net7257 net5222 _06731_ VGND VGND VPWR VPWR _06737_ sky130_fd_sc_hd__or3_1
XFILLER_0_56_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23758_ net4616 net4922 VGND VGND VPWR VPWR _03624_ sky130_fd_sc_hd__nand2_1
X_13511_ _05698_ net622 net625 VGND VGND VPWR VPWR _05782_ sky130_fd_sc_hd__a21o_1
XFILLER_0_137_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22709_ _02647_ pid_d.mult0.a\[13\] net3094 VGND VGND VPWR VPWR _02648_ sky130_fd_sc_hd__mux2_1
X_14491_ net7324 net5279 VGND VGND VPWR VPWR _06675_ sky130_fd_sc_hd__xnor2_2
X_23689_ net933 _03555_ VGND VGND VPWR VPWR _03556_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16230_ _08267_ _08294_ VGND VGND VPWR VPWR _08295_ sky130_fd_sc_hd__xnor2_2
X_13442_ _05506_ _05507_ net7769 net1584 VGND VGND VPWR VPWR _05715_ sky130_fd_sc_hd__o211a_1
X_25428_ clknet_leaf_97_clk _00311_ net8380 VGND VGND VPWR VPWR matmul0.sin\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13373_ net1130 _05643_ VGND VGND VPWR VPWR _05646_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_141_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16161_ _08138_ _08148_ VGND VGND VPWR VPWR _08227_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25359_ clknet_leaf_56_clk _00242_ net8718 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult2\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire6030 net6028 VGND VGND VPWR VPWR net6030 sky130_fd_sc_hd__clkbuf_2
X_15112_ _06964_ _07061_ VGND VGND VPWR VPWR _07186_ sky130_fd_sc_hd__nor2_1
Xwire6052 net6057 VGND VGND VPWR VPWR net6052 sky130_fd_sc_hd__buf_1
X_16092_ net572 _08157_ VGND VGND VPWR VPWR _08159_ sky130_fd_sc_hd__nor2_1
Xfanout4533 net4546 VGND VGND VPWR VPWR net4533 sky130_fd_sc_hd__clkbuf_1
Xwire6074 net6075 VGND VGND VPWR VPWR net6074 sky130_fd_sc_hd__clkbuf_1
Xwire5340 pid_d.out\[11\] VGND VGND VPWR VPWR net5340 sky130_fd_sc_hd__buf_1
Xwire6085 net6084 VGND VGND VPWR VPWR net6085 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_181_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5351 net5352 VGND VGND VPWR VPWR net5351 sky130_fd_sc_hd__clkbuf_1
X_19920_ net6110 _11686_ _11690_ VGND VGND VPWR VPWR _11752_ sky130_fd_sc_hd__or3_1
XFILLER_0_32_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15043_ net4176 net4174 net4205 net4204 VGND VGND VPWR VPWR _07117_ sky130_fd_sc_hd__o22a_1
Xwire5362 pid_d.out\[6\] VGND VGND VPWR VPWR net5362 sky130_fd_sc_hd__clkbuf_1
Xwire5373 pid_d.ki\[15\] VGND VGND VPWR VPWR net5373 sky130_fd_sc_hd__clkbuf_1
Xfanout4577 pid_q.mult0.a\[10\] VGND VGND VPWR VPWR net4577 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout4588 net4594 VGND VGND VPWR VPWR net4588 sky130_fd_sc_hd__buf_1
XFILLER_0_43_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4650 net4652 VGND VGND VPWR VPWR net4650 sky130_fd_sc_hd__clkbuf_1
Xwire5395 net5396 VGND VGND VPWR VPWR net5395 sky130_fd_sc_hd__buf_1
X_19851_ net6127 net2506 _11642_ VGND VGND VPWR VPWR _11684_ sky130_fd_sc_hd__or3_1
Xwire4661 net4667 VGND VGND VPWR VPWR net4661 sky130_fd_sc_hd__clkbuf_1
Xwire4672 pid_q.mult0.a\[6\] VGND VGND VPWR VPWR net4672 sky130_fd_sc_hd__clkbuf_1
Xwire4683 net4684 VGND VGND VPWR VPWR net4683 sky130_fd_sc_hd__buf_1
Xwire4694 net4695 VGND VGND VPWR VPWR net4694 sky130_fd_sc_hd__buf_1
Xwire3960 net3961 VGND VGND VPWR VPWR net3960 sky130_fd_sc_hd__buf_1
X_18802_ _10644_ _10645_ VGND VGND VPWR VPWR _10646_ sky130_fd_sc_hd__or2b_1
X_19782_ _11542_ net604 _11609_ VGND VGND VPWR VPWR _11616_ sky130_fd_sc_hd__or3b_1
X_16994_ _08836_ net4057 _08955_ VGND VGND VPWR VPWR _08956_ sky130_fd_sc_hd__a21o_1
Xwire3982 net3983 VGND VGND VPWR VPWR net3982 sky130_fd_sc_hd__buf_1
Xwire3993 _09634_ VGND VGND VPWR VPWR net3993 sky130_fd_sc_hd__buf_1
X_18733_ _10533_ _10573_ _10574_ _10577_ net6975 VGND VGND VPWR VPWR _10578_ sky130_fd_sc_hd__a32o_1
X_15945_ _07995_ _07987_ VGND VGND VPWR VPWR _08013_ sky130_fd_sc_hd__and2b_1
X_18664_ _10502_ _10510_ VGND VGND VPWR VPWR _10511_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15876_ _07769_ _07943_ _07944_ VGND VGND VPWR VPWR _07945_ sky130_fd_sc_hd__o21a_1
XFILLER_0_188_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17615_ net6734 svm0.tB\[2\] VGND VGND VPWR VPWR _09496_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14827_ _06930_ VGND VGND VPWR VPWR _00185_ sky130_fd_sc_hd__clkbuf_1
X_18595_ net6771 net2129 net3281 VGND VGND VPWR VPWR _10443_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17546_ net6698 _09425_ _09427_ VGND VGND VPWR VPWR _09428_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14758_ net7448 _06887_ _06888_ net7454 net3621 VGND VGND VPWR VPWR _06889_ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13709_ _05971_ _05977_ VGND VGND VPWR VPWR _05978_ sky130_fd_sc_hd__xnor2_1
X_17477_ net3273 _09368_ net6661 VGND VGND VPWR VPWR _09369_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14689_ net7155 _06836_ VGND VGND VPWR VPWR _06837_ sky130_fd_sc_hd__xnor2_1
X_19216_ net3205 net6225 net3901 _11049_ _11052_ VGND VGND VPWR VPWR _11053_ sky130_fd_sc_hd__a32o_1
XFILLER_0_6_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16428_ matmul0.matmul_stage_inst.mult1\[12\] net209 net3475 VGND VGND VPWR VPWR
+ _08490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19147_ _10983_ _10797_ VGND VGND VPWR VPWR _10984_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16359_ _08339_ _08347_ _08349_ VGND VGND VPWR VPWR _08422_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19078_ net6357 net3908 _10829_ _10912_ net6249 VGND VGND VPWR VPWR _10915_ sky130_fd_sc_hd__o221a_1
XFILLER_0_14_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6491 net6497 VGND VGND VPWR VPWR net6491 sky130_fd_sc_hd__clkbuf_2
X_18029_ net4043 net3943 VGND VGND VPWR VPWR _09880_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21040_ net5541 _01032_ _01033_ VGND VGND VPWR VPWR _01056_ sky130_fd_sc_hd__or3_1
Xwire1309 _05779_ VGND VGND VPWR VPWR net1309 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22991_ _02863_ VGND VGND VPWR VPWR _00662_ sky130_fd_sc_hd__clkbuf_1
X_24730_ net8012 _04557_ _04562_ VGND VGND VPWR VPWR _04563_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21942_ _01847_ _01848_ _01949_ VGND VGND VPWR VPWR _01950_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_173_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24661_ pid_q.curr_error\[2\] net2382 net1372 VGND VGND VPWR VPWR _04513_ sky130_fd_sc_hd__and3_1
X_21873_ _01880_ _01881_ VGND VGND VPWR VPWR _01882_ sky130_fd_sc_hd__and2_1
XFILLER_0_173_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length6005 net6006 VGND VGND VPWR VPWR net6005 sky130_fd_sc_hd__buf_1
XFILLER_0_55_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23612_ _03478_ _03479_ net7510 VGND VGND VPWR VPWR _03480_ sky130_fd_sc_hd__o21a_1
Xmax_length6027 net6024 VGND VGND VPWR VPWR net6027 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_82_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20824_ net5795 net5544 VGND VGND VPWR VPWR _00840_ sky130_fd_sc_hd__nand2_2
X_24592_ _04446_ _04447_ VGND VGND VPWR VPWR _04448_ sky130_fd_sc_hd__or2b_1
Xmax_length5304 net5305 VGND VGND VPWR VPWR net5304 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23543_ net4619 net4962 VGND VGND VPWR VPWR _03411_ sky130_fd_sc_hd__nand2_2
Xwire8905 net8906 VGND VGND VPWR VPWR net8905 sky130_fd_sc_hd__buf_1
X_20755_ net5931 net5472 VGND VGND VPWR VPWR _12526_ sky130_fd_sc_hd__nand2_2
Xwire8916 net8917 VGND VGND VPWR VPWR net8916 sky130_fd_sc_hd__buf_1
XFILLER_0_147_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8927 net112 VGND VGND VPWR VPWR net8927 sky130_fd_sc_hd__clkbuf_1
Xwire8938 net8939 VGND VGND VPWR VPWR net8938 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23474_ _03283_ _03284_ _03342_ VGND VGND VPWR VPWR _03343_ sky130_fd_sc_hd__a21oi_1
Xwire8949 net8950 VGND VGND VPWR VPWR net8949 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20686_ net6077 net1496 _12460_ VGND VGND VPWR VPWR _12462_ sky130_fd_sc_hd__and3_1
Xwire606 net607 VGND VGND VPWR VPWR net606 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire617 _09135_ VGND VGND VPWR VPWR net617 sky130_fd_sc_hd__clkbuf_2
Xwire628 _05635_ VGND VGND VPWR VPWR net628 sky130_fd_sc_hd__buf_1
XFILLER_0_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire639 _03488_ VGND VGND VPWR VPWR net639 sky130_fd_sc_hd__buf_1
XFILLER_0_162_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22425_ net3777 _02425_ _02426_ VGND VGND VPWR VPWR _02427_ sky130_fd_sc_hd__or3_1
XFILLER_0_134_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25213_ clknet_leaf_61_clk _00102_ net8717 VGND VGND VPWR VPWR svm0.vC\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3946 _09879_ VGND VGND VPWR VPWR net3946 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22356_ _02290_ _02295_ _02288_ VGND VGND VPWR VPWR _02359_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_149_Right_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25144_ clknet_leaf_65_clk _00033_ net8655 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__dfstp_1
XFILLER_0_21_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21307_ _00860_ _00875_ net1052 VGND VGND VPWR VPWR _01322_ sky130_fd_sc_hd__a21bo_1
X_25075_ net4418 net1633 net291 net1629 _04821_ VGND VGND VPWR VPWR _00788_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22287_ _01317_ net5646 VGND VGND VPWR VPWR _02291_ sky130_fd_sc_hd__nand2_2
X_24026_ _03885_ _03888_ VGND VGND VPWR VPWR _03889_ sky130_fd_sc_hd__xor2_1
Xwire3201 _10871_ VGND VGND VPWR VPWR net3201 sky130_fd_sc_hd__buf_1
Xhold270 pid_q.prev_int\[9\] VGND VGND VPWR VPWR net9223 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3212 _10821_ VGND VGND VPWR VPWR net3212 sky130_fd_sc_hd__buf_1
X_21238_ net705 net703 VGND VGND VPWR VPWR _01253_ sky130_fd_sc_hd__and2_1
Xwire3223 net3224 VGND VGND VPWR VPWR net3223 sky130_fd_sc_hd__buf_1
Xhold281 pid_d.ki\[7\] VGND VGND VPWR VPWR net9234 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3234 _09955_ VGND VGND VPWR VPWR net3234 sky130_fd_sc_hd__buf_1
Xhold292 cordic0.sin\[6\] VGND VGND VPWR VPWR net9245 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3245 _09730_ VGND VGND VPWR VPWR net3245 sky130_fd_sc_hd__clkbuf_2
Xwire2511 _11149_ VGND VGND VPWR VPWR net2511 sky130_fd_sc_hd__buf_1
Xwire3256 _09649_ VGND VGND VPWR VPWR net3256 sky130_fd_sc_hd__dlymetal6s2s_1
X_21169_ net5628 net5882 _01181_ VGND VGND VPWR VPWR _01185_ sky130_fd_sc_hd__a21o_1
Xwire2522 _10978_ VGND VGND VPWR VPWR net2522 sky130_fd_sc_hd__buf_1
Xwire3267 net3268 VGND VGND VPWR VPWR net3267 sky130_fd_sc_hd__buf_1
Xwire3278 net3279 VGND VGND VPWR VPWR net3278 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2533 net2534 VGND VGND VPWR VPWR net2533 sky130_fd_sc_hd__clkbuf_2
Xwire2544 _10099_ VGND VGND VPWR VPWR net2544 sky130_fd_sc_hd__buf_1
Xwire1810 net1811 VGND VGND VPWR VPWR net1810 sky130_fd_sc_hd__clkbuf_1
Xwire2555 net2556 VGND VGND VPWR VPWR net2555 sky130_fd_sc_hd__clkbuf_2
Xwire2566 _09517_ VGND VGND VPWR VPWR net2566 sky130_fd_sc_hd__clkbuf_1
Xwire1821 _08911_ VGND VGND VPWR VPWR net1821 sky130_fd_sc_hd__buf_1
Xwire2577 net2578 VGND VGND VPWR VPWR net2577 sky130_fd_sc_hd__buf_1
X_13991_ _06251_ _06255_ VGND VGND VPWR VPWR _06256_ sky130_fd_sc_hd__xnor2_1
Xwire1832 net1833 VGND VGND VPWR VPWR net1832 sky130_fd_sc_hd__clkbuf_1
Xwire1843 net1844 VGND VGND VPWR VPWR net1843 sky130_fd_sc_hd__clkbuf_1
Xwire2588 net2589 VGND VGND VPWR VPWR net2588 sky130_fd_sc_hd__buf_1
XFILLER_0_137_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2599 _09004_ VGND VGND VPWR VPWR net2599 sky130_fd_sc_hd__buf_1
Xwire1854 net1855 VGND VGND VPWR VPWR net1854 sky130_fd_sc_hd__buf_1
XFILLER_0_99_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15730_ net888 _07667_ _07708_ VGND VGND VPWR VPWR _07801_ sky130_fd_sc_hd__o21a_1
Xwire1865 _07482_ VGND VGND VPWR VPWR net1865 sky130_fd_sc_hd__buf_1
X_24928_ pid_q.ki\[5\] _04712_ net1360 VGND VGND VPWR VPWR _04713_ sky130_fd_sc_hd__mux2_1
X_12942_ net7939 net2356 net1978 VGND VGND VPWR VPWR _05215_ sky130_fd_sc_hd__and3_1
Xwire1876 _07363_ VGND VGND VPWR VPWR net1876 sky130_fd_sc_hd__clkbuf_1
Xwire1887 net1888 VGND VGND VPWR VPWR net1887 sky130_fd_sc_hd__clkbuf_1
Xwire1898 net1899 VGND VGND VPWR VPWR net1898 sky130_fd_sc_hd__clkbuf_2
X_15661_ _07712_ _07732_ VGND VGND VPWR VPWR _07733_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24859_ _04663_ VGND VGND VPWR VPWR _00730_ sky130_fd_sc_hd__clkbuf_1
X_12873_ _05144_ _05145_ VGND VGND VPWR VPWR _05146_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17400_ net613 _09305_ _09303_ VGND VGND VPWR VPWR _09306_ sky130_fd_sc_hd__a21oi_1
X_14612_ _06512_ net6443 VGND VGND VPWR VPWR _06784_ sky130_fd_sc_hd__nand2_1
X_18380_ net7043 _09704_ net3241 VGND VGND VPWR VPWR _10231_ sky130_fd_sc_hd__mux2_1
Xmax_length7273 net7274 VGND VGND VPWR VPWR net7273 sky130_fd_sc_hd__clkbuf_1
X_15592_ net1854 net1853 VGND VGND VPWR VPWR _07664_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17331_ net6730 net7828 VGND VGND VPWR VPWR _09245_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14543_ net7278 _06711_ VGND VGND VPWR VPWR _06722_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6594 net6595 VGND VGND VPWR VPWR net6594 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_139_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17262_ _09192_ VGND VGND VPWR VPWR _09193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14474_ _06659_ _06657_ _06658_ VGND VGND VPWR VPWR _06661_ sky130_fd_sc_hd__and3_1
XFILLER_0_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19001_ net6295 net3898 VGND VGND VPWR VPWR _10838_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length5893 net5894 VGND VGND VPWR VPWR net5893 sky130_fd_sc_hd__buf_1
X_16213_ net2655 net3442 net2697 net3522 VGND VGND VPWR VPWR _08278_ sky130_fd_sc_hd__o211a_1
X_13425_ _05695_ net728 VGND VGND VPWR VPWR _05698_ sky130_fd_sc_hd__xnor2_2
X_17193_ net2592 net3305 VGND VGND VPWR VPWR _09143_ sky130_fd_sc_hd__nand2_1
X_16144_ net774 _08209_ VGND VGND VPWR VPWR _08210_ sky130_fd_sc_hd__xnor2_1
X_13356_ _05509_ _05627_ _05628_ VGND VGND VPWR VPWR _05629_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_116_Right_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16075_ net2662 _08028_ VGND VGND VPWR VPWR _08142_ sky130_fd_sc_hd__nand2_1
X_13287_ _05467_ _05468_ _05465_ _05464_ VGND VGND VPWR VPWR _05560_ sky130_fd_sc_hd__o211a_1
Xfanout4352 net4369 VGND VGND VPWR VPWR net4352 sky130_fd_sc_hd__buf_1
Xwire5170 net5171 VGND VGND VPWR VPWR net5170 sky130_fd_sc_hd__clkbuf_2
Xwire5181 net5182 VGND VGND VPWR VPWR net5181 sky130_fd_sc_hd__buf_1
X_19903_ _11720_ _11734_ VGND VGND VPWR VPWR _11735_ sky130_fd_sc_hd__nor2_1
X_15026_ _07099_ VGND VGND VPWR VPWR _07100_ sky130_fd_sc_hd__clkbuf_1
Xwire5192 matmul0.beta_pass\[15\] VGND VGND VPWR VPWR net5192 sky130_fd_sc_hd__buf_1
Xwire4480 pid_q.ki\[9\] VGND VGND VPWR VPWR net4480 sky130_fd_sc_hd__clkbuf_1
Xwire4491 net4487 VGND VGND VPWR VPWR net4491 sky130_fd_sc_hd__buf_1
X_19834_ _11601_ _11604_ _11600_ VGND VGND VPWR VPWR _11668_ sky130_fd_sc_hd__o21a_1
XFILLER_0_127_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3790 net3791 VGND VGND VPWR VPWR net3790 sky130_fd_sc_hd__clkbuf_1
X_16977_ _08923_ _08939_ VGND VGND VPWR VPWR _08940_ sky130_fd_sc_hd__xor2_1
X_19765_ _11574_ _11599_ VGND VGND VPWR VPWR _11600_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_39_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput5 angle_in[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
X_15928_ _07926_ _07996_ VGND VGND VPWR VPWR _07997_ sky130_fd_sc_hd__xnor2_1
X_18716_ _10493_ net1195 _10495_ VGND VGND VPWR VPWR _10562_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_190_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19696_ _11500_ _11531_ VGND VGND VPWR VPWR _11532_ sky130_fd_sc_hd__xnor2_2
X_18647_ _10441_ net1069 net1070 VGND VGND VPWR VPWR _10494_ sky130_fd_sc_hd__o21ba_1
X_15859_ net2700 net2761 net2671 _07837_ VGND VGND VPWR VPWR _07928_ sky130_fd_sc_hd__o31a_1
XFILLER_0_143_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18578_ net6934 _10171_ _10364_ VGND VGND VPWR VPWR _10426_ sky130_fd_sc_hd__nor3_1
XFILLER_0_59_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17529_ net6686 _09268_ _09411_ VGND VGND VPWR VPWR _09413_ sky130_fd_sc_hd__or3_1
XFILLER_0_4_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20540_ _12323_ _12324_ net2079 VGND VGND VPWR VPWR _12325_ sky130_fd_sc_hd__a21o_1
XFILLER_0_145_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20471_ net3353 net9153 _12260_ _12261_ VGND VGND VPWR VPWR _00499_ sky130_fd_sc_hd__a211o_1
XFILLER_0_171_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22210_ net5747 net5404 VGND VGND VPWR VPWR _02215_ sky130_fd_sc_hd__nand2_2
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23190_ _03057_ _03059_ VGND VGND VPWR VPWR _03060_ sky130_fd_sc_hd__xnor2_1
Xmax_length1818 net1819 VGND VGND VPWR VPWR net1818 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22141_ net1389 _02146_ VGND VGND VPWR VPWR _02147_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22072_ net2062 net945 VGND VGND VPWR VPWR _02079_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_112_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25900_ clknet_leaf_17_clk _00773_ net8628 VGND VGND VPWR VPWR pid_q.kp\[12\] sky130_fd_sc_hd__dfrtp_1
X_21023_ net5640 net5820 VGND VGND VPWR VPWR _01039_ sky130_fd_sc_hd__and2_1
XFILLER_0_61_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1106 net1107 VGND VGND VPWR VPWR net1106 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25831_ clknet_leaf_36_clk _00704_ net8752 VGND VGND VPWR VPWR pid_q.curr_error\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1117 _07163_ VGND VGND VPWR VPWR net1117 sky130_fd_sc_hd__buf_1
Xwire1128 _05712_ VGND VGND VPWR VPWR net1128 sky130_fd_sc_hd__buf_1
Xwire1139 _05377_ VGND VGND VPWR VPWR net1139 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25762_ clknet_leaf_95_clk _00635_ net8455 VGND VGND VPWR VPWR pid_d.out\[3\] sky130_fd_sc_hd__dfrtp_2
X_22974_ matmul0.beta_pass\[6\] net972 net6573 VGND VGND VPWR VPWR _02855_ sky130_fd_sc_hd__mux2_1
X_24713_ net8023 net1158 VGND VGND VPWR VPWR _04549_ sky130_fd_sc_hd__xnor2_1
X_21925_ net5719 net5479 VGND VGND VPWR VPWR _01933_ sky130_fd_sc_hd__nand2_2
X_25693_ clknet_leaf_3_clk _00566_ net8569 VGND VGND VPWR VPWR pid_d.curr_error\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_24644_ _04441_ net631 VGND VGND VPWR VPWR _04499_ sky130_fd_sc_hd__nand2_1
XFILLER_0_179_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21856_ net5406 net5376 _01864_ net5839 VGND VGND VPWR VPWR _01865_ sky130_fd_sc_hd__o22a_1
XFILLER_0_167_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout8629 net8642 VGND VGND VPWR VPWR net8629 sky130_fd_sc_hd__buf_1
XFILLER_0_132_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20807_ _00819_ _00822_ VGND VGND VPWR VPWR _00823_ sky130_fd_sc_hd__xnor2_1
X_24575_ net4918 net4896 VGND VGND VPWR VPWR _04431_ sky130_fd_sc_hd__xnor2_1
X_21787_ net5896 net3108 net5385 VGND VGND VPWR VPWR _01797_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4400 pid_q.out\[14\] VGND VGND VPWR VPWR net4400 sky130_fd_sc_hd__buf_1
Xwire8713 net8712 VGND VGND VPWR VPWR net8713 sky130_fd_sc_hd__buf_1
Xwire8724 net8725 VGND VGND VPWR VPWR net8724 sky130_fd_sc_hd__clkbuf_1
X_23526_ net5163 net4496 VGND VGND VPWR VPWR _03394_ sky130_fd_sc_hd__nand2_1
Xwire8735 net8736 VGND VGND VPWR VPWR net8735 sky130_fd_sc_hd__clkbuf_1
Xwire8746 net8743 VGND VGND VPWR VPWR net8746 sky130_fd_sc_hd__buf_1
X_20738_ net5525 net5867 VGND VGND VPWR VPWR _12509_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire403 _06365_ VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__buf_1
Xwire8757 net8758 VGND VGND VPWR VPWR net8757 sky130_fd_sc_hd__buf_1
Xmax_length5189 net5190 VGND VGND VPWR VPWR net5189 sky130_fd_sc_hd__clkbuf_2
Xwire8768 net8767 VGND VGND VPWR VPWR net8768 sky130_fd_sc_hd__buf_1
XFILLER_0_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4466 pid_q.out\[2\] VGND VGND VPWR VPWR net4466 sky130_fd_sc_hd__buf_1
Xwire414 _01907_ VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__clkbuf_1
Xwire8779 net8780 VGND VGND VPWR VPWR net8779 sky130_fd_sc_hd__buf_1
Xwire425 _07924_ VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__buf_1
Xmax_length4477 pid_q.kp\[9\] VGND VGND VPWR VPWR net4477 sky130_fd_sc_hd__clkbuf_1
X_23457_ _03322_ _03325_ VGND VGND VPWR VPWR _03326_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_136_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20669_ _12431_ _12434_ net6109 VGND VGND VPWR VPWR _12446_ sky130_fd_sc_hd__o21a_1
Xwire436 net437 VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__clkbuf_1
Xwire447 _07640_ VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__clkbuf_1
Xwire458 net459 VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13210_ _05431_ _05479_ VGND VGND VPWR VPWR _05483_ sky130_fd_sc_hd__and2b_1
Xwire469 net470 VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__clkbuf_1
X_22408_ _02337_ _02409_ net551 VGND VGND VPWR VPWR _02410_ sky130_fd_sc_hd__o21ba_1
X_14190_ _06439_ _06449_ VGND VGND VPWR VPWR _06450_ sky130_fd_sc_hd__xnor2_2
X_23388_ _03223_ net2428 _03257_ VGND VGND VPWR VPWR _03258_ sky130_fd_sc_hd__o21ai_1
Xmax_length3787 net3788 VGND VGND VPWR VPWR net3787 sky130_fd_sc_hd__buf_1
XFILLER_0_115_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13141_ net7845 net2304 net2964 VGND VGND VPWR VPWR _05414_ sky130_fd_sc_hd__and3_1
X_25127_ net9134 _04849_ net2391 net5974 VGND VGND VPWR VPWR _00808_ sky130_fd_sc_hd__a22o_1
X_22339_ net3829 net2472 net5762 VGND VGND VPWR VPWR _02342_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13072_ _05343_ _05344_ _05052_ VGND VGND VPWR VPWR _05345_ sky130_fd_sc_hd__o21ai_1
X_25058_ net3732 _04806_ VGND VGND VPWR VPWR _04807_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3020 net3021 VGND VGND VPWR VPWR net3020 sky130_fd_sc_hd__buf_1
Xwire3031 net3032 VGND VGND VPWR VPWR net3031 sky130_fd_sc_hd__buf_1
X_16900_ net6371 _08861_ _08863_ VGND VGND VPWR VPWR _08864_ sky130_fd_sc_hd__o21ai_1
Xwire3042 _03791_ VGND VGND VPWR VPWR net3042 sky130_fd_sc_hd__clkbuf_1
X_24009_ _03870_ _03871_ net3741 VGND VGND VPWR VPWR _03872_ sky130_fd_sc_hd__a21oi_1
Xwire3053 net3054 VGND VGND VPWR VPWR net3053 sky130_fd_sc_hd__buf_1
X_17880_ net3977 _09664_ VGND VGND VPWR VPWR _09731_ sky130_fd_sc_hd__nor2_1
Xwire3064 net3067 VGND VGND VPWR VPWR net3064 sky130_fd_sc_hd__buf_1
Xwire3075 _02678_ VGND VGND VPWR VPWR net3075 sky130_fd_sc_hd__clkbuf_1
Xwire2330 net2331 VGND VGND VPWR VPWR net2330 sky130_fd_sc_hd__buf_1
XFILLER_0_40_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2341 net2342 VGND VGND VPWR VPWR net2341 sky130_fd_sc_hd__buf_1
X_16831_ _08806_ VGND VGND VPWR VPWR _00313_ sky130_fd_sc_hd__clkbuf_1
Xwire3097 net3098 VGND VGND VPWR VPWR net3097 sky130_fd_sc_hd__clkbuf_1
Xwire2352 net2353 VGND VGND VPWR VPWR net2352 sky130_fd_sc_hd__clkbuf_1
Xwire2374 net2375 VGND VGND VPWR VPWR net2374 sky130_fd_sc_hd__buf_1
XFILLER_0_189_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1640 net1641 VGND VGND VPWR VPWR net1640 sky130_fd_sc_hd__buf_1
Xwire2385 _04858_ VGND VGND VPWR VPWR net2385 sky130_fd_sc_hd__buf_1
X_19550_ _11384_ _11386_ VGND VGND VPWR VPWR _11387_ sky130_fd_sc_hd__nand2_1
Xwire1651 _04281_ VGND VGND VPWR VPWR net1651 sky130_fd_sc_hd__clkbuf_4
Xwire2396 _04753_ VGND VGND VPWR VPWR net2396 sky130_fd_sc_hd__buf_1
X_16762_ net4291 VGND VGND VPWR VPWR _08770_ sky130_fd_sc_hd__clkbuf_2
Xwire1662 _03599_ VGND VGND VPWR VPWR net1662 sky130_fd_sc_hd__buf_1
X_13974_ net7642 net1311 _06238_ VGND VGND VPWR VPWR _06239_ sky130_fd_sc_hd__and3_1
Xwire1673 _03364_ VGND VGND VPWR VPWR net1673 sky130_fd_sc_hd__clkbuf_1
Xwire1684 net1685 VGND VGND VPWR VPWR net1684 sky130_fd_sc_hd__clkbuf_1
X_18501_ net3286 net6799 VGND VGND VPWR VPWR _10350_ sky130_fd_sc_hd__nor2_1
X_15713_ net2735 _07133_ net3398 net3411 net2685 VGND VGND VPWR VPWR _07784_ sky130_fd_sc_hd__a32o_1
Xwire1695 net1696 VGND VGND VPWR VPWR net1695 sky130_fd_sc_hd__clkbuf_1
X_12925_ _05196_ _05107_ _05197_ VGND VGND VPWR VPWR _05198_ sky130_fd_sc_hd__a21o_1
X_19481_ _10851_ _11264_ _11317_ VGND VGND VPWR VPWR _11318_ sky130_fd_sc_hd__o21a_1
X_16693_ _08722_ _08718_ matmul0.matmul_stage_inst.mult2\[10\] VGND VGND VPWR VPWR
+ _08723_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_158_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18432_ net3966 _10224_ VGND VGND VPWR VPWR _10282_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_14_Left_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15644_ net2821 net3426 net2696 VGND VGND VPWR VPWR _07716_ sky130_fd_sc_hd__and3_1
X_12856_ net2966 VGND VGND VPWR VPWR _05129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length7070 net7071 VGND VGND VPWR VPWR net7070 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18363_ _10212_ _10213_ net6842 VGND VGND VPWR VPWR _10214_ sky130_fd_sc_hd__mux2_1
X_15575_ net2799 net3427 VGND VGND VPWR VPWR _07647_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12787_ _04959_ _05059_ VGND VGND VPWR VPWR _05060_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17314_ _09221_ _09222_ _09225_ _09227_ VGND VGND VPWR VPWR _09228_ sky130_fd_sc_hd__o31a_1
X_14526_ net1625 _06705_ VGND VGND VPWR VPWR _06706_ sky130_fd_sc_hd__nand2_1
X_18294_ net963 _10144_ _09836_ VGND VGND VPWR VPWR _10145_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_113_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17245_ net2165 net288 net1800 net9054 VGND VGND VPWR VPWR _00343_ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14457_ net6454 matmul0.op_in\[0\] _06513_ net6447 VGND VGND VPWR VPWR _06647_ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13408_ net452 _05660_ _05673_ _05676_ _05680_ VGND VGND VPWR VPWR _05681_ sky130_fd_sc_hd__o32a_1
XFILLER_0_52_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17176_ net6901 _09102_ _09126_ VGND VGND VPWR VPWR _09128_ sky130_fd_sc_hd__or3_1
X_14388_ net8198 net3636 VGND VGND VPWR VPWR _06594_ sky130_fd_sc_hd__and2_1
Xwire970 net971 VGND VGND VPWR VPWR net970 sky130_fd_sc_hd__buf_1
Xwire981 net982 VGND VGND VPWR VPWR net981 sky130_fd_sc_hd__buf_1
XFILLER_0_84_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire992 net993 VGND VGND VPWR VPWR net992 sky130_fd_sc_hd__buf_1
XFILLER_0_141_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16127_ _08121_ _08122_ _08192_ VGND VGND VPWR VPWR _08193_ sky130_fd_sc_hd__o21a_1
X_13339_ _05606_ net1320 VGND VGND VPWR VPWR _05612_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_23_Left_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16058_ _08121_ _08124_ VGND VGND VPWR VPWR _08125_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15009_ _07079_ _07081_ _07076_ VGND VGND VPWR VPWR _07083_ sky130_fd_sc_hd__a21oi_1
X_19817_ net2500 _11650_ VGND VGND VPWR VPWR _11651_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19748_ net2104 _11582_ VGND VGND VPWR VPWR _11583_ sky130_fd_sc_hd__xor2_1
XFILLER_0_56_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19679_ net6200 _11466_ VGND VGND VPWR VPWR _11515_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21710_ _01718_ _01720_ VGND VGND VPWR VPWR _01721_ sky130_fd_sc_hd__xnor2_1
X_22690_ pid_d.ki\[7\] net2440 net2993 pid_d.kp\[7\] VGND VGND VPWR VPWR _02635_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21641_ _01603_ _01650_ _01651_ VGND VGND VPWR VPWR _01652_ sky130_fd_sc_hd__a21o_1
Xwire8009 net8010 VGND VGND VPWR VPWR net8009 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24360_ net2405 _04135_ _04218_ VGND VGND VPWR VPWR _04219_ sky130_fd_sc_hd__a21oi_1
X_21572_ net1727 _01477_ _01478_ VGND VGND VPWR VPWR _01584_ sky130_fd_sc_hd__o21ai_1
Xwire7308 net7309 VGND VGND VPWR VPWR net7308 sky130_fd_sc_hd__clkbuf_1
Xmax_length3006 _00000_ VGND VGND VPWR VPWR net3006 sky130_fd_sc_hd__buf_1
XFILLER_0_170_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7319 net7320 VGND VGND VPWR VPWR net7319 sky130_fd_sc_hd__clkbuf_1
X_23311_ net697 net755 VGND VGND VPWR VPWR _03181_ sky130_fd_sc_hd__or2_1
Xmax_length3017 net3018 VGND VGND VPWR VPWR net3017 sky130_fd_sc_hd__buf_1
X_20523_ net6324 _12304_ VGND VGND VPWR VPWR _12309_ sky130_fd_sc_hd__nand2_1
X_24291_ _04144_ _04150_ VGND VGND VPWR VPWR _04151_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6607 net6608 VGND VGND VPWR VPWR net6607 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length2316 _05035_ VGND VGND VPWR VPWR net2316 sky130_fd_sc_hd__buf_1
XFILLER_0_104_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23242_ _03107_ _03111_ VGND VGND VPWR VPWR _03112_ sky130_fd_sc_hd__xnor2_2
X_20454_ net1830 _12246_ net8044 VGND VGND VPWR VPWR _12247_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5906 net5907 VGND VGND VPWR VPWR net5906 sky130_fd_sc_hd__clkbuf_2
Xmax_length1626 _04860_ VGND VGND VPWR VPWR net1626 sky130_fd_sc_hd__buf_1
X_23173_ _03035_ _03037_ _03042_ VGND VGND VPWR VPWR _03043_ sky130_fd_sc_hd__a21o_1
X_20385_ net1054 _12169_ _12183_ VGND VGND VPWR VPWR _12184_ sky130_fd_sc_hd__nor3_1
XFILLER_0_31_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22124_ net5745 net5411 VGND VGND VPWR VPWR _02130_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput150 net150 VGND VGND VPWR VPWR pwmB_out sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22055_ _01948_ _01950_ _01946_ VGND VGND VPWR VPWR _02062_ sky130_fd_sc_hd__a21bo_1
X_21006_ _00966_ _00944_ VGND VGND VPWR VPWR _01022_ sky130_fd_sc_hd__xnor2_1
X_25814_ clknet_leaf_32_clk _00687_ net8680 VGND VGND VPWR VPWR pid_q.prev_error\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25745_ clknet_leaf_8_clk _00618_ net8553 VGND VGND VPWR VPWR pid_d.kp\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22957_ pid_d.out\[14\] pid_d.curr_int\[14\] VGND VGND VPWR VPWR _02845_ sky130_fd_sc_hd__nor2_1
X_12710_ _04980_ _04981_ _04982_ VGND VGND VPWR VPWR _04983_ sky130_fd_sc_hd__a21o_1
X_21908_ pid_d.prev_int\[7\] VGND VGND VPWR VPWR _01916_ sky130_fd_sc_hd__inv_2
X_13690_ _05900_ _05902_ _05958_ VGND VGND VPWR VPWR _05959_ sky130_fd_sc_hd__a21o_1
X_25676_ clknet_leaf_6_clk _00549_ net8561 VGND VGND VPWR VPWR pid_d.prev_error\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22888_ net346 net2033 _02782_ VGND VGND VPWR VPWR _02783_ sky130_fd_sc_hd__a21o_1
XFILLER_0_194_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24627_ net3745 net4807 _04475_ VGND VGND VPWR VPWR _04482_ sky130_fd_sc_hd__a21o_1
X_12641_ net7825 net2357 net1979 VGND VGND VPWR VPWR _04914_ sky130_fd_sc_hd__and3_1
X_21839_ net5784 net5431 VGND VGND VPWR VPWR _01848_ sky130_fd_sc_hd__nand2_1
Xfanout8426 net8432 VGND VGND VPWR VPWR net8426 sky130_fd_sc_hd__buf_1
Xfanout8459 net8484 VGND VGND VPWR VPWR net8459 sky130_fd_sc_hd__clkbuf_2
X_15360_ _07412_ _07432_ _07415_ VGND VGND VPWR VPWR _07434_ sky130_fd_sc_hd__or3b_1
Xwire8521 net8522 VGND VGND VPWR VPWR net8521 sky130_fd_sc_hd__clkbuf_1
X_24558_ _04342_ _04353_ _04413_ VGND VGND VPWR VPWR _04414_ sky130_fd_sc_hd__o21a_1
X_12572_ net7531 VGND VGND VPWR VPWR _04861_ sky130_fd_sc_hd__inv_2
Xwire8532 net8533 VGND VGND VPWR VPWR net8532 sky130_fd_sc_hd__clkbuf_2
Xwire8543 net8544 VGND VGND VPWR VPWR net8543 sky130_fd_sc_hd__clkbuf_1
X_14311_ _06532_ VGND VGND VPWR VPWR _06533_ sky130_fd_sc_hd__buf_1
Xwire200 _04382_ VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__buf_1
X_23509_ _03376_ _03377_ VGND VGND VPWR VPWR _03378_ sky130_fd_sc_hd__nand2_1
Xfanout7769 net7774 VGND VGND VPWR VPWR net7769 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_124_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire211 net212 VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_1
Xwire222 _06216_ VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__clkbuf_1
Xwire8576 net8577 VGND VGND VPWR VPWR net8576 sky130_fd_sc_hd__clkbuf_1
X_15291_ net1274 _07364_ VGND VGND VPWR VPWR _07365_ sky130_fd_sc_hd__xnor2_1
X_24489_ _04344_ _04345_ VGND VGND VPWR VPWR _04346_ sky130_fd_sc_hd__xor2_1
Xwire7842 net7835 VGND VGND VPWR VPWR net7842 sky130_fd_sc_hd__clkbuf_1
Xwire8587 net8588 VGND VGND VPWR VPWR net8587 sky130_fd_sc_hd__buf_1
XFILLER_0_136_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire233 net234 VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkbuf_1
Xwire7853 net7854 VGND VGND VPWR VPWR net7853 sky130_fd_sc_hd__buf_1
Xwire8598 net8599 VGND VGND VPWR VPWR net8598 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17030_ net1809 VGND VGND VPWR VPWR _08990_ sky130_fd_sc_hd__buf_1
Xwire244 _11987_ VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__buf_1
Xwire255 _06360_ VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__buf_1
Xwire7864 net7865 VGND VGND VPWR VPWR net7864 sky130_fd_sc_hd__clkbuf_1
X_14242_ net152 _06497_ net6451 VGND VGND VPWR VPWR _06498_ sky130_fd_sc_hd__a21o_1
Xwire7875 net7876 VGND VGND VPWR VPWR net7875 sky130_fd_sc_hd__buf_1
Xwire266 net267 VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__clkbuf_1
Xwire7886 net7887 VGND VGND VPWR VPWR net7886 sky130_fd_sc_hd__clkbuf_1
Xwire277 net278 VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__clkbuf_1
Xmax_length3584 net3585 VGND VGND VPWR VPWR net3584 sky130_fd_sc_hd__buf_1
Xwire288 net289 VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__buf_1
Xwire299 net300 VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__buf_1
XFILLER_0_180_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14173_ net217 _06369_ _06422_ _06421_ VGND VGND VPWR VPWR _06433_ sky130_fd_sc_hd__a31o_1
XFILLER_0_104_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2894 net2895 VGND VGND VPWR VPWR net2894 sky130_fd_sc_hd__buf_1
X_13124_ _05379_ _05396_ VGND VGND VPWR VPWR _05397_ sky130_fd_sc_hd__xnor2_1
X_18981_ _10795_ net3214 VGND VGND VPWR VPWR _10818_ sky130_fd_sc_hd__xnor2_1
X_13055_ _05079_ _05327_ _05002_ VGND VGND VPWR VPWR _05328_ sky130_fd_sc_hd__or3_1
X_17932_ net2559 _09782_ _09780_ _09678_ VGND VGND VPWR VPWR _09783_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_178_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17863_ net7064 net2142 _09713_ VGND VGND VPWR VPWR _09714_ sky130_fd_sc_hd__a21oi_1
Xwire2160 _09191_ VGND VGND VPWR VPWR net2160 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2171 net2172 VGND VGND VPWR VPWR net2171 sky130_fd_sc_hd__clkbuf_2
X_19602_ net6087 net6045 VGND VGND VPWR VPWR _11439_ sky130_fd_sc_hd__nand2_1
Xwire2182 net2183 VGND VGND VPWR VPWR net2182 sky130_fd_sc_hd__clkbuf_1
X_16814_ _08797_ VGND VGND VPWR VPWR _00305_ sky130_fd_sc_hd__clkbuf_1
Xwire2193 net2194 VGND VGND VPWR VPWR net2193 sky130_fd_sc_hd__clkbuf_1
X_17794_ net7108 net7133 VGND VGND VPWR VPWR _09645_ sky130_fd_sc_hd__xor2_1
XFILLER_0_75_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1481 net1482 VGND VGND VPWR VPWR net1481 sky130_fd_sc_hd__buf_1
X_19533_ _11254_ _11369_ VGND VGND VPWR VPWR _11370_ sky130_fd_sc_hd__and2_1
X_16745_ _08761_ VGND VGND VPWR VPWR _00272_ sky130_fd_sc_hd__clkbuf_1
X_13957_ net7642 _06221_ VGND VGND VPWR VPWR _06222_ sky130_fd_sc_hd__nand2_1
Xwire1492 net1494 VGND VGND VPWR VPWR net1492 sky130_fd_sc_hd__clkbuf_1
X_12908_ _05177_ _05180_ VGND VGND VPWR VPWR _05181_ sky130_fd_sc_hd__xnor2_2
X_19464_ _11254_ _11300_ VGND VGND VPWR VPWR _11301_ sky130_fd_sc_hd__or2_1
X_16676_ net7281 net720 net6549 VGND VGND VPWR VPWR _08709_ sky130_fd_sc_hd__mux2_1
X_13888_ _06081_ _06142_ net532 VGND VGND VPWR VPWR _06154_ sky130_fd_sc_hd__o21a_1
XFILLER_0_124_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15627_ net3513 net3508 net4216 net4214 VGND VGND VPWR VPWR _07699_ sky130_fd_sc_hd__o22a_1
X_18415_ _10192_ _10195_ VGND VGND VPWR VPWR _10265_ sky130_fd_sc_hd__xnor2_1
X_12839_ net7931 net1958 net1957 _05111_ VGND VGND VPWR VPWR _05112_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19395_ _11168_ _11184_ VGND VGND VPWR VPWR _11232_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18346_ _10192_ _10193_ _10131_ VGND VGND VPWR VPWR _10197_ sky130_fd_sc_hd__o21a_1
X_15558_ _07629_ _07630_ VGND VGND VPWR VPWR _07631_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14509_ _06655_ _06689_ _06690_ net893 net9005 VGND VGND VPWR VPWR _00107_ sky130_fd_sc_hd__a32o_1
X_18277_ _10115_ _10116_ _10126_ VGND VGND VPWR VPWR _10128_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15489_ _07475_ _07554_ VGND VGND VPWR VPWR _07562_ sky130_fd_sc_hd__and2b_1
X_17228_ net6799 VGND VGND VPWR VPWR _09176_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput30 currA_in[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput41 currB_in[2] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_1
Xinput52 currT_in[12] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_1
Xinput63 currT_in[8] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput74 periodTop[3] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_1
X_17159_ net2595 _09095_ _09111_ net6484 VGND VGND VPWR VPWR _09112_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput85 pid_d_addr[13] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_1
Xinput96 pid_d_addr[9] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20170_ net6100 net6042 VGND VGND VPWR VPWR _11996_ sky130_fd_sc_hd__nor2_1
XFILLER_0_196_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23860_ _03595_ _03597_ _03593_ VGND VGND VPWR VPWR _03725_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_74_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length8529 net8518 VGND VGND VPWR VPWR net8529 sky130_fd_sc_hd__clkbuf_1
X_22811_ _02714_ VGND VGND VPWR VPWR _00631_ sky130_fd_sc_hd__clkbuf_1
X_23791_ net744 _03559_ _03562_ VGND VGND VPWR VPWR _03657_ sky130_fd_sc_hd__o21a_1
Xmax_length7839 net7840 VGND VGND VPWR VPWR net7839 sky130_fd_sc_hd__clkbuf_1
X_25530_ clknet_leaf_35_clk _00410_ net8764 VGND VGND VPWR VPWR svm0.state\[0\] sky130_fd_sc_hd__dfrtp_1
X_22742_ pid_d.ki\[5\] _02672_ net1689 VGND VGND VPWR VPWR _02673_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25461_ clknet_leaf_68_clk _00001_ net8454 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.start
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_181_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22673_ _02623_ VGND VGND VPWR VPWR _00584_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24412_ _04222_ _04225_ _04269_ VGND VGND VPWR VPWR _04270_ sky130_fd_sc_hd__o21a_1
X_21624_ net5970 VGND VGND VPWR VPWR _01636_ sky130_fd_sc_hd__inv_2
XFILLER_0_192_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25392_ clknet_leaf_82_clk _00275_ net8508 VGND VGND VPWR VPWR matmul0.b\[11\] sky130_fd_sc_hd__dfrtp_1
Xwire7105 net7103 VGND VGND VPWR VPWR net7105 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire7116 net7117 VGND VGND VPWR VPWR net7116 sky130_fd_sc_hd__buf_1
XFILLER_0_75_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24343_ net4895 net4504 VGND VGND VPWR VPWR _04202_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21555_ _01561_ _01566_ VGND VGND VPWR VPWR _01567_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_191_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7138 net7134 VGND VGND VPWR VPWR net7138 sky130_fd_sc_hd__buf_1
Xwire6404 net6405 VGND VGND VPWR VPWR net6404 sky130_fd_sc_hd__buf_1
Xwire7149 net7150 VGND VGND VPWR VPWR net7149 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire6415 cordic0.slte0.opB\[6\] VGND VGND VPWR VPWR net6415 sky130_fd_sc_hd__buf_1
XFILLER_0_160_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20506_ _08836_ net3849 net3345 net6766 VGND VGND VPWR VPWR _12293_ sky130_fd_sc_hd__a211o_1
X_24274_ _04132_ _04133_ VGND VGND VPWR VPWR _04134_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6437 net6438 VGND VGND VPWR VPWR net6437 sky130_fd_sc_hd__clkbuf_1
X_21486_ _01379_ _01384_ _01498_ VGND VGND VPWR VPWR _01499_ sky130_fd_sc_hd__a21o_1
Xwire5703 net5704 VGND VGND VPWR VPWR net5703 sky130_fd_sc_hd__buf_1
Xmax_length2146 _09577_ VGND VGND VPWR VPWR net2146 sky130_fd_sc_hd__buf_1
Xwire5714 net5715 VGND VGND VPWR VPWR net5714 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2157 net2158 VGND VGND VPWR VPWR net2157 sky130_fd_sc_hd__buf_1
X_23225_ net5038 net4717 VGND VGND VPWR VPWR _03095_ sky130_fd_sc_hd__nand2_1
Xwire5725 net5729 VGND VGND VPWR VPWR net5725 sky130_fd_sc_hd__clkbuf_1
X_20437_ net6370 _12230_ _12231_ VGND VGND VPWR VPWR _00495_ sky130_fd_sc_hd__a21bo_1
Xwire5736 net5737 VGND VGND VPWR VPWR net5736 sky130_fd_sc_hd__clkbuf_1
Xwire5747 net5748 VGND VGND VPWR VPWR net5747 sky130_fd_sc_hd__buf_1
XFILLER_0_114_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5769 net5766 VGND VGND VPWR VPWR net5769 sky130_fd_sc_hd__buf_1
XFILLER_0_28_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23156_ _03014_ _03025_ VGND VGND VPWR VPWR _03026_ sky130_fd_sc_hd__xnor2_2
X_20368_ net2608 _12167_ VGND VGND VPWR VPWR _12168_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22107_ _02111_ _02112_ VGND VGND VPWR VPWR _02113_ sky130_fd_sc_hd__xnor2_1
X_23087_ _02890_ _02891_ VGND VGND VPWR VPWR _02957_ sky130_fd_sc_hd__nand2_1
X_20299_ cordic0.slte0.opA\[1\] net2281 _12103_ VGND VGND VPWR VPWR _12105_ sky130_fd_sc_hd__or3_1
XFILLER_0_101_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22038_ _01933_ _01935_ _02044_ VGND VGND VPWR VPWR _02045_ sky130_fd_sc_hd__a21oi_2
X_14860_ _06947_ VGND VGND VPWR VPWR _00201_ sky130_fd_sc_hd__clkbuf_1
X_13811_ net780 _05987_ _06078_ VGND VGND VPWR VPWR _06079_ sky130_fd_sc_hd__o21ai_1
X_14791_ net3624 matmul0.cos\[0\] net2878 net2855 VGND VGND VPWR VPWR _06912_ sky130_fd_sc_hd__o211a_1
X_23989_ _03852_ _03764_ pid_q.prev_error\[5\] VGND VGND VPWR VPWR _03853_ sky130_fd_sc_hd__o21ba_1
X_16530_ _08548_ _08588_ VGND VGND VPWR VPWR _08590_ sky130_fd_sc_hd__or2_1
X_13742_ net404 _06010_ VGND VGND VPWR VPWR _06011_ sky130_fd_sc_hd__xnor2_1
X_25728_ clknet_leaf_8_clk _00601_ net8551 VGND VGND VPWR VPWR pid_d.ki\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16461_ net976 VGND VGND VPWR VPWR _08522_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13673_ _05938_ _05941_ VGND VGND VPWR VPWR _05942_ sky130_fd_sc_hd__xnor2_2
X_25659_ clknet_leaf_25_clk _00532_ net8579 VGND VGND VPWR VPWR pid_d.curr_int\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_128_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18200_ net2547 _10049_ _10050_ VGND VGND VPWR VPWR _10051_ sky130_fd_sc_hd__nand3_1
XFILLER_0_156_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15412_ net4095 net4094 VGND VGND VPWR VPWR _07486_ sky130_fd_sc_hd__or2_1
XFILLER_0_167_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12624_ _04896_ VGND VGND VPWR VPWR _04897_ sky130_fd_sc_hd__buf_6
X_19180_ _10958_ _10959_ _11012_ VGND VGND VPWR VPWR _11017_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16392_ net2772 net2642 VGND VGND VPWR VPWR _08454_ sky130_fd_sc_hd__nand2_1
XFILLER_0_182_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18131_ _09916_ _09921_ _09922_ VGND VGND VPWR VPWR _09982_ sky130_fd_sc_hd__or3b_1
Xwire8340 net8338 VGND VGND VPWR VPWR net8340 sky130_fd_sc_hd__dlymetal6s2s_1
X_15343_ net2811 net2782 net3487 net2716 VGND VGND VPWR VPWR _07417_ sky130_fd_sc_hd__a211o_1
XFILLER_0_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8373 net8369 VGND VGND VPWR VPWR net8373 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6843 cordic0.vec\[1\]\[14\] VGND VGND VPWR VPWR net6843 sky130_fd_sc_hd__clkbuf_1
Xwire8384 net8383 VGND VGND VPWR VPWR net8384 sky130_fd_sc_hd__buf_1
XFILLER_0_81_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7650 net7649 VGND VGND VPWR VPWR net7650 sky130_fd_sc_hd__buf_1
X_18062_ _09908_ _09912_ VGND VGND VPWR VPWR _09913_ sky130_fd_sc_hd__xnor2_1
Xfanout6854 net6869 VGND VGND VPWR VPWR net6854 sky130_fd_sc_hd__buf_1
Xwire8395 net8394 VGND VGND VPWR VPWR net8395 sky130_fd_sc_hd__clkbuf_2
Xwire7661 net7663 VGND VGND VPWR VPWR net7661 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_0_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15274_ _07346_ _07347_ VGND VGND VPWR VPWR _07348_ sky130_fd_sc_hd__xnor2_1
Xwire7672 net7674 VGND VGND VPWR VPWR net7672 sky130_fd_sc_hd__buf_1
XFILLER_0_123_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6876 net6878 VGND VGND VPWR VPWR net6876 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17013_ net3345 _08968_ _08972_ _08973_ net5993 VGND VGND VPWR VPWR _08974_ sky130_fd_sc_hd__a32o_1
Xfanout6887 cordic0.vec\[1\]\[12\] VGND VGND VPWR VPWR net6887 sky130_fd_sc_hd__buf_1
Xwire7694 net7697 VGND VGND VPWR VPWR net7694 sky130_fd_sc_hd__clkbuf_1
X_14225_ net1119 _06470_ net7626 VGND VGND VPWR VPWR _06483_ sky130_fd_sc_hd__a21o_1
Xwire6960 cordic0.vec\[1\]\[9\] VGND VGND VPWR VPWR net6960 sky130_fd_sc_hd__buf_1
Xwire6971 net6972 VGND VGND VPWR VPWR net6971 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6982 net6984 VGND VGND VPWR VPWR net6982 sky130_fd_sc_hd__buf_1
X_14156_ _06415_ _06416_ VGND VGND VPWR VPWR _06417_ sky130_fd_sc_hd__or2_1
XFILLER_0_186_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13107_ _05255_ _05260_ VGND VGND VPWR VPWR _05380_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14087_ _06346_ _06348_ VGND VGND VPWR VPWR _06350_ sky130_fd_sc_hd__or2_1
X_18964_ net6222 net6241 VGND VGND VPWR VPWR _10801_ sky130_fd_sc_hd__and2_1
X_13038_ net791 net736 VGND VGND VPWR VPWR _05311_ sky130_fd_sc_hd__or2_1
X_17915_ _09653_ _09668_ net1781 _09765_ VGND VGND VPWR VPWR _09766_ sky130_fd_sc_hd__a22o_1
X_18895_ net3283 net3934 VGND VGND VPWR VPWR _10736_ sky130_fd_sc_hd__nand2_1
XFILLER_0_178_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17846_ net7027 net3970 VGND VGND VPWR VPWR _09697_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_135_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17777_ _08985_ _09627_ VGND VGND VPWR VPWR _09628_ sky130_fd_sc_hd__xnor2_1
X_14989_ net4210 net4208 VGND VGND VPWR VPWR _07063_ sky130_fd_sc_hd__or2_1
XFILLER_0_178_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19516_ net1060 _11352_ VGND VGND VPWR VPWR _11353_ sky130_fd_sc_hd__xnor2_2
X_16728_ _08752_ VGND VGND VPWR VPWR _00264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19447_ _11261_ _11282_ _11283_ VGND VGND VPWR VPWR _11284_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16659_ _08692_ _08688_ _08693_ VGND VGND VPWR VPWR _08694_ sky130_fd_sc_hd__a21o_1
XFILLER_0_146_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19378_ net2509 _11213_ _11214_ net6276 VGND VGND VPWR VPWR _11215_ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18329_ _10168_ _10179_ VGND VGND VPWR VPWR _10180_ sky130_fd_sc_hd__xnor2_1
Xfanout8790 net8801 VGND VGND VPWR VPWR net8790 sky130_fd_sc_hd__buf_1
XFILLER_0_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21340_ net5638 net5654 VGND VGND VPWR VPWR _01354_ sky130_fd_sc_hd__or2b_1
XFILLER_0_71_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21271_ _00840_ _00841_ _01285_ VGND VGND VPWR VPWR _01286_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_114_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23010_ _02876_ _02879_ VGND VGND VPWR VPWR _02880_ sky130_fd_sc_hd__xnor2_1
X_20222_ _12042_ VGND VGND VPWR VPWR _00469_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3619 net3620 VGND VGND VPWR VPWR net3619 sky130_fd_sc_hd__buf_1
X_20153_ _11934_ _11979_ _11954_ VGND VGND VPWR VPWR _11980_ sky130_fd_sc_hd__a21o_1
Xwire2907 net2908 VGND VGND VPWR VPWR net2907 sky130_fd_sc_hd__clkbuf_1
Xwire2918 net2919 VGND VGND VPWR VPWR net2918 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2929 net2930 VGND VGND VPWR VPWR net2929 sky130_fd_sc_hd__clkbuf_1
X_24961_ net1635 VGND VGND VPWR VPWR _04735_ sky130_fd_sc_hd__buf_1
X_20084_ _11910_ _11912_ VGND VGND VPWR VPWR _11913_ sky130_fd_sc_hd__nand2_1
X_23912_ _03759_ VGND VGND VPWR VPWR _03776_ sky130_fd_sc_hd__inv_2
X_24892_ pid_q.ki\[12\] net3710 net3700 pid_q.kp\[12\] VGND VGND VPWR VPWR _04686_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23843_ net1660 _03707_ VGND VGND VPWR VPWR _03708_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_196_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23774_ net1019 net1018 _03509_ VGND VGND VPWR VPWR _03640_ sky130_fd_sc_hd__a21bo_1
X_20986_ net5547 net5884 _01001_ VGND VGND VPWR VPWR _01002_ sky130_fd_sc_hd__and3_1
XFILLER_0_196_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25513_ clknet_leaf_43_clk _00393_ net8783 VGND VGND VPWR VPWR svm0.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6935 net6932 VGND VGND VPWR VPWR net6935 sky130_fd_sc_hd__clkbuf_1
X_22725_ _02654_ net3764 net2434 VGND VGND VPWR VPWR _02661_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_67_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6957 net6952 VGND VGND VPWR VPWR net6957 sky130_fd_sc_hd__buf_1
XFILLER_0_95_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25444_ clknet_leaf_114_clk _00327_ net8333 VGND VGND VPWR VPWR cordic0.vec\[1\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_22656_ net3089 _02584_ _02600_ VGND VGND VPWR VPWR _02613_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21607_ net948 _01515_ _01618_ VGND VGND VPWR VPWR _01619_ sky130_fd_sc_hd__a21o_1
XFILLER_0_180_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25375_ clknet_leaf_57_clk _00258_ net8716 VGND VGND VPWR VPWR matmul0.alpha_pass\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22587_ _02548_ _02564_ _02565_ net2044 net8957 VGND VGND VPWR VPWR _00556_ sky130_fd_sc_hd__a32o_1
Xwire6201 net6200 VGND VGND VPWR VPWR net6201 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_168_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24326_ net7464 net238 _04185_ _04118_ VGND VGND VPWR VPWR _04186_ sky130_fd_sc_hd__a211o_1
XFILLER_0_90_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21538_ _01329_ _01423_ _01548_ VGND VGND VPWR VPWR _01550_ sky130_fd_sc_hd__a21o_1
Xwire6234 net6235 VGND VGND VPWR VPWR net6234 sky130_fd_sc_hd__clkbuf_1
Xwire5500 net5502 VGND VGND VPWR VPWR net5500 sky130_fd_sc_hd__buf_1
Xwire6245 net6246 VGND VGND VPWR VPWR net6245 sky130_fd_sc_hd__clkbuf_2
Xfanout4715 net4725 VGND VGND VPWR VPWR net4715 sky130_fd_sc_hd__buf_1
Xwire5511 net5505 VGND VGND VPWR VPWR net5511 sky130_fd_sc_hd__buf_1
Xwire5522 pid_d.mult0.a\[8\] VGND VGND VPWR VPWR net5522 sky130_fd_sc_hd__clkbuf_1
X_24257_ pid_q.curr_int\[10\] VGND VGND VPWR VPWR _04117_ sky130_fd_sc_hd__inv_2
Xwire6267 net6264 VGND VGND VPWR VPWR net6267 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_120_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21469_ net1729 _01370_ _01481_ VGND VGND VPWR VPWR _01482_ sky130_fd_sc_hd__a21o_1
Xwire5533 net5534 VGND VGND VPWR VPWR net5533 sky130_fd_sc_hd__clkbuf_1
Xwire6278 net6279 VGND VGND VPWR VPWR net6278 sky130_fd_sc_hd__clkbuf_1
X_14010_ _06156_ _06273_ VGND VGND VPWR VPWR _06274_ sky130_fd_sc_hd__nor2_1
Xwire6289 net6286 VGND VGND VPWR VPWR net6289 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire5544 net5545 VGND VGND VPWR VPWR net5544 sky130_fd_sc_hd__buf_1
Xfanout4759 net4764 VGND VGND VPWR VPWR net4759 sky130_fd_sc_hd__clkbuf_1
X_23208_ _03076_ _03077_ VGND VGND VPWR VPWR _03078_ sky130_fd_sc_hd__xnor2_1
Xwire5555 pid_d.mult0.a\[6\] VGND VGND VPWR VPWR net5555 sky130_fd_sc_hd__clkbuf_1
Xwire5566 net5567 VGND VGND VPWR VPWR net5566 sky130_fd_sc_hd__buf_1
Xwire4832 net4840 VGND VGND VPWR VPWR net4832 sky130_fd_sc_hd__buf_1
X_24188_ _04003_ _04014_ _04005_ VGND VGND VPWR VPWR _04049_ sky130_fd_sc_hd__a21o_1
Xwire5577 net5578 VGND VGND VPWR VPWR net5577 sky130_fd_sc_hd__buf_1
Xwire5588 net5589 VGND VGND VPWR VPWR net5588 sky130_fd_sc_hd__clkbuf_1
Xwire4854 net4855 VGND VGND VPWR VPWR net4854 sky130_fd_sc_hd__clkbuf_1
Xwire5599 net5595 VGND VGND VPWR VPWR net5599 sky130_fd_sc_hd__buf_1
X_23139_ _02965_ _03008_ VGND VGND VPWR VPWR _03009_ sky130_fd_sc_hd__xor2_1
Xwire4865 net4866 VGND VGND VPWR VPWR net4865 sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_length1297 net1298 VGND VGND VPWR VPWR net1297 sky130_fd_sc_hd__clkbuf_2
Xwire4876 net4877 VGND VGND VPWR VPWR net4876 sky130_fd_sc_hd__buf_1
Xwire4887 net4888 VGND VGND VPWR VPWR net4887 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4898 net4897 VGND VGND VPWR VPWR net4898 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15961_ _08027_ _08028_ VGND VGND VPWR VPWR _08029_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17700_ net7489 net3270 net8864 VGND VGND VPWR VPWR _09576_ sky130_fd_sc_hd__o21a_1
X_14912_ net4196 net4194 net3595 net3593 VGND VGND VPWR VPWR _06986_ sky130_fd_sc_hd__o22a_1
X_15892_ net984 _07960_ VGND VGND VPWR VPWR _07961_ sky130_fd_sc_hd__xor2_1
X_18680_ net3231 net2131 VGND VGND VPWR VPWR _10526_ sky130_fd_sc_hd__and2_1
X_17631_ _09510_ _09511_ _09488_ _09489_ VGND VGND VPWR VPWR _09512_ sky130_fd_sc_hd__o2bb2a_1
X_14843_ _06938_ VGND VGND VPWR VPWR _00193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17562_ _09393_ svm0.tC\[11\] _09441_ _09443_ VGND VGND VPWR VPWR _09444_ sky130_fd_sc_hd__a211o_1
Xmax_length8871 net8872 VGND VGND VPWR VPWR net8871 sky130_fd_sc_hd__buf_1
XFILLER_0_58_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14774_ matmul0.sin\[10\] net1908 net3616 VGND VGND VPWR VPWR _06900_ sky130_fd_sc_hd__o21a_1
X_19301_ _11136_ _11137_ net3887 VGND VGND VPWR VPWR _11138_ sky130_fd_sc_hd__mux2_1
X_16513_ net2665 _08511_ _08513_ VGND VGND VPWR VPWR _08573_ sky130_fd_sc_hd__o21a_1
X_13725_ _05925_ _05929_ VGND VGND VPWR VPWR _05994_ sky130_fd_sc_hd__nand2_1
X_17493_ _09303_ net770 net4027 VGND VGND VPWR VPWR _09382_ sky130_fd_sc_hd__o21a_1
XFILLER_0_169_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19232_ _11033_ _11068_ VGND VGND VPWR VPWR _11069_ sky130_fd_sc_hd__xnor2_1
X_16444_ _08453_ VGND VGND VPWR VPWR _08505_ sky130_fd_sc_hd__inv_2
XFILLER_0_195_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13656_ _05924_ _05925_ VGND VGND VPWR VPWR _05926_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout8064 cordic0.state\[0\] VGND VGND VPWR VPWR net8064 sky130_fd_sc_hd__buf_1
XFILLER_0_186_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19163_ _10995_ _10961_ _10999_ VGND VGND VPWR VPWR _11000_ sky130_fd_sc_hd__or3_1
X_12607_ matmul0.matmul_stage_inst.state\[0\] matmul0.matmul_stage_inst.start VGND
+ VGND VPWR VPWR _04883_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16375_ _08408_ net1087 net1079 VGND VGND VPWR VPWR _08437_ sky130_fd_sc_hd__mux2_1
X_13587_ svm0.tC\[1\] net1127 net287 net1927 VGND VGND VPWR VPWR _00018_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8170 net8171 VGND VGND VPWR VPWR net8170 sky130_fd_sc_hd__clkbuf_1
X_18114_ net3235 VGND VGND VPWR VPWR _09965_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15326_ net2256 net2252 _07399_ VGND VGND VPWR VPWR _07400_ sky130_fd_sc_hd__a21o_1
Xwire8181 net8182 VGND VGND VPWR VPWR net8181 sky130_fd_sc_hd__clkbuf_1
X_19094_ net6268 net3192 net3885 net6319 VGND VGND VPWR VPWR _10931_ sky130_fd_sc_hd__o22a_1
Xwire8192 net8193 VGND VGND VPWR VPWR net8192 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7480 net7482 VGND VGND VPWR VPWR net7480 sky130_fd_sc_hd__buf_1
X_18045_ _09887_ _09893_ _09895_ VGND VGND VPWR VPWR _09896_ sky130_fd_sc_hd__o21ba_1
Xwire7491 net7492 VGND VGND VPWR VPWR net7491 sky130_fd_sc_hd__clkbuf_1
X_15257_ net1276 _07296_ _07292_ VGND VGND VPWR VPWR _07331_ sky130_fd_sc_hd__o21a_1
X_14208_ _06439_ _06442_ VGND VGND VPWR VPWR _06467_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6790 net6791 VGND VGND VPWR VPWR net6790 sky130_fd_sc_hd__clkbuf_1
Xfanout5994 net6015 VGND VGND VPWR VPWR net5994 sky130_fd_sc_hd__clkbuf_1
X_15188_ _07259_ _07255_ _07235_ VGND VGND VPWR VPWR _07262_ sky130_fd_sc_hd__nor3_1
X_14139_ _06349_ net834 _06375_ VGND VGND VPWR VPWR _06400_ sky130_fd_sc_hd__a21o_1
X_19996_ _11782_ VGND VGND VPWR VPWR _11827_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18947_ net6375 net207 VGND VGND VPWR VPWR _10785_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18878_ _10718_ _10719_ VGND VGND VPWR VPWR _10720_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_6_Left_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17829_ net7065 net7032 VGND VGND VPWR VPWR _09680_ sky130_fd_sc_hd__nand2_1
X_20840_ _00852_ _00855_ VGND VGND VPWR VPWR _00856_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_178_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20771_ net5612 net5760 VGND VGND VPWR VPWR _12542_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22510_ _02451_ _02450_ _02510_ VGND VGND VPWR VPWR _02511_ sky130_fd_sc_hd__o21a_1
XFILLER_0_71_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23490_ net4749 net4845 VGND VGND VPWR VPWR _03359_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22441_ net2060 _02442_ VGND VGND VPWR VPWR _02443_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_88_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25160_ clknet_leaf_44_clk _00049_ net8785 VGND VGND VPWR VPWR pid_q.target\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_190_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22372_ net5380 _02374_ VGND VGND VPWR VPWR _02375_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24111_ _03879_ _03881_ _03972_ VGND VGND VPWR VPWR _03973_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_72_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21323_ net5984 pid_d.prev_int\[1\] VGND VGND VPWR VPWR _01337_ sky130_fd_sc_hd__or2_1
X_25091_ net198 _04829_ _04834_ _04835_ VGND VGND VPWR VPWR _00790_ sky130_fd_sc_hd__o211ai_1
Xwire4106 net4107 VGND VGND VPWR VPWR net4106 sky130_fd_sc_hd__clkbuf_1
X_24042_ _03903_ _03904_ VGND VGND VPWR VPWR _03905_ sky130_fd_sc_hd__or2_1
Xwire4117 net4118 VGND VGND VPWR VPWR net4117 sky130_fd_sc_hd__buf_1
X_21254_ _01263_ _01268_ VGND VGND VPWR VPWR _01269_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4128 net4129 VGND VGND VPWR VPWR net4128 sky130_fd_sc_hd__clkbuf_1
Xwire4139 _07025_ VGND VGND VPWR VPWR net4139 sky130_fd_sc_hd__buf_1
X_20205_ net179 _12029_ VGND VGND VPWR VPWR _12030_ sky130_fd_sc_hd__xnor2_1
Xwire3416 net3417 VGND VGND VPWR VPWR net3416 sky130_fd_sc_hd__buf_1
X_21185_ _01167_ _01186_ _01199_ _01200_ VGND VGND VPWR VPWR _01201_ sky130_fd_sc_hd__a22o_1
Xwire3427 net3428 VGND VGND VPWR VPWR net3427 sky130_fd_sc_hd__buf_1
Xwire3438 _07371_ VGND VGND VPWR VPWR net3438 sky130_fd_sc_hd__buf_1
XFILLER_0_99_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2704 _07320_ VGND VGND VPWR VPWR net2704 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2715 _07287_ VGND VGND VPWR VPWR net2715 sky130_fd_sc_hd__clkbuf_1
X_20136_ net3126 _11963_ VGND VGND VPWR VPWR _11964_ sky130_fd_sc_hd__and2b_1
Xwire2726 net2729 VGND VGND VPWR VPWR net2726 sky130_fd_sc_hd__buf_1
Xwire2737 net2738 VGND VGND VPWR VPWR net2737 sky130_fd_sc_hd__clkbuf_1
Xwire2748 _07207_ VGND VGND VPWR VPWR net2748 sky130_fd_sc_hd__buf_1
XFILLER_0_95_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2759 _07204_ VGND VGND VPWR VPWR net2759 sky130_fd_sc_hd__buf_1
X_24944_ _04723_ VGND VGND VPWR VPWR _00755_ sky130_fd_sc_hd__clkbuf_1
X_20067_ _11894_ _11895_ VGND VGND VPWR VPWR _11896_ sky130_fd_sc_hd__nand2_1
X_24875_ _04674_ net4646 net1996 VGND VGND VPWR VPWR _04675_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length7400 matmul0.matmul_stage_inst.e\[1\] VGND VGND VPWR VPWR net7400 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_174_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23826_ net4562 net4997 _03689_ _03690_ VGND VGND VPWR VPWR _03691_ sky130_fd_sc_hd__a31o_1
Xmax_length7422 matmul0.matmul_stage_inst.b\[9\] VGND VGND VPWR VPWR net7422 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23757_ net4665 net4875 VGND VGND VPWR VPWR _03623_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20969_ _00945_ _00946_ VGND VGND VPWR VPWR _00985_ sky130_fd_sc_hd__xnor2_1
X_13510_ net534 _05770_ _05771_ VGND VGND VPWR VPWR _05781_ sky130_fd_sc_hd__o21bai_1
X_22708_ pid_d.ki\[13\] net3705 _04886_ pid_d.kp\[13\] VGND VGND VPWR VPWR _02647_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14490_ net7336 net5286 VGND VGND VPWR VPWR _06674_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length6776 net6772 VGND VGND VPWR VPWR net6776 sky130_fd_sc_hd__clkbuf_1
X_23688_ net1165 _03554_ VGND VGND VPWR VPWR _03555_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_166_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length6798 net6799 VGND VGND VPWR VPWR net6798 sky130_fd_sc_hd__buf_1
XFILLER_0_83_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13441_ _05704_ _05713_ VGND VGND VPWR VPWR _05714_ sky130_fd_sc_hd__xnor2_1
X_25427_ clknet_leaf_98_clk _00310_ net8380 VGND VGND VPWR VPWR matmul0.sin\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_192_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22639_ net3767 VGND VGND VPWR VPWR _02604_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16160_ _08140_ net1256 _08225_ VGND VGND VPWR VPWR _08226_ sky130_fd_sc_hd__o21a_1
X_13372_ _05541_ _05542_ _05637_ VGND VGND VPWR VPWR _05645_ sky130_fd_sc_hd__a21o_1
X_25358_ clknet_leaf_56_clk _00241_ net8723 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult2\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire6020 net6023 VGND VGND VPWR VPWR net6020 sky130_fd_sc_hd__buf_1
XFILLER_0_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15111_ _07111_ _07184_ VGND VGND VPWR VPWR _07185_ sky130_fd_sc_hd__xnor2_1
X_24309_ _04045_ _04106_ _04168_ VGND VGND VPWR VPWR _04169_ sky130_fd_sc_hd__nor3_1
Xwire6042 net6041 VGND VGND VPWR VPWR net6042 sky130_fd_sc_hd__dlymetal6s2s_1
X_16091_ net572 _08157_ VGND VGND VPWR VPWR _08158_ sky130_fd_sc_hd__and2_1
Xwire6053 net6054 VGND VGND VPWR VPWR net6053 sky130_fd_sc_hd__clkbuf_1
X_25289_ clknet_leaf_89_clk _00172_ net8422 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.d\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire5330 net5331 VGND VGND VPWR VPWR net5330 sky130_fd_sc_hd__clkbuf_1
Xwire6075 net6076 VGND VGND VPWR VPWR net6075 sky130_fd_sc_hd__buf_1
Xwire5341 net5342 VGND VGND VPWR VPWR net5341 sky130_fd_sc_hd__clkbuf_1
Xwire6086 net6087 VGND VGND VPWR VPWR net6086 sky130_fd_sc_hd__buf_1
X_15042_ net4181 net4180 net3595 net3593 VGND VGND VPWR VPWR _07116_ sky130_fd_sc_hd__o22a_1
XFILLER_0_142_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5352 net5353 VGND VGND VPWR VPWR net5352 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout4556 pid_q.mult0.a\[11\] VGND VGND VPWR VPWR net4556 sky130_fd_sc_hd__buf_1
Xwire6097 net6098 VGND VGND VPWR VPWR net6097 sky130_fd_sc_hd__clkbuf_2
Xwire4640 net4639 VGND VGND VPWR VPWR net4640 sky130_fd_sc_hd__clkbuf_1
Xwire5385 net5386 VGND VGND VPWR VPWR net5385 sky130_fd_sc_hd__buf_1
XFILLER_0_103_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4651 net4652 VGND VGND VPWR VPWR net4651 sky130_fd_sc_hd__buf_1
Xwire5396 net5397 VGND VGND VPWR VPWR net5396 sky130_fd_sc_hd__buf_1
X_19850_ net6127 _11642_ VGND VGND VPWR VPWR _11683_ sky130_fd_sc_hd__nand2_1
Xwire4662 net4666 VGND VGND VPWR VPWR net4662 sky130_fd_sc_hd__buf_1
XFILLER_0_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4684 net4685 VGND VGND VPWR VPWR net4684 sky130_fd_sc_hd__buf_1
X_18801_ _10640_ _10643_ VGND VGND VPWR VPWR _10645_ sky130_fd_sc_hd__nand2_1
Xwire4695 net4692 VGND VGND VPWR VPWR net4695 sky130_fd_sc_hd__clkbuf_1
Xwire3950 _09876_ VGND VGND VPWR VPWR net3950 sky130_fd_sc_hd__clkbuf_1
Xwire3961 net3962 VGND VGND VPWR VPWR net3961 sky130_fd_sc_hd__buf_1
X_19781_ _11488_ _11609_ VGND VGND VPWR VPWR _11615_ sky130_fd_sc_hd__and2b_1
X_16993_ net6461 net4048 VGND VGND VPWR VPWR _08955_ sky130_fd_sc_hd__nand2_1
Xwire3972 _09689_ VGND VGND VPWR VPWR net3972 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_79_Left_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire3983 net3984 VGND VGND VPWR VPWR net3983 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3994 net3995 VGND VGND VPWR VPWR net3994 sky130_fd_sc_hd__buf_1
X_18732_ net3298 _10575_ _10576_ VGND VGND VPWR VPWR _10577_ sky130_fd_sc_hd__a21o_1
X_15944_ _07987_ _07995_ VGND VGND VPWR VPWR _08012_ sky130_fd_sc_hd__or2b_1
XFILLER_0_183_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15875_ net2714 net3422 _07694_ net2813 VGND VGND VPWR VPWR _07944_ sky130_fd_sc_hd__a22o_1
X_18663_ net422 net714 _10503_ _10509_ VGND VGND VPWR VPWR _10510_ sky130_fd_sc_hd__o31a_1
XFILLER_0_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17614_ net6734 svm0.tB\[2\] VGND VGND VPWR VPWR _09495_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14826_ matmul0.a\[2\] matmul0.matmul_stage_inst.e\[2\] net3610 VGND VGND VPWR VPWR
+ _06930_ sky130_fd_sc_hd__mux2_1
X_18594_ net6865 net2589 net6771 net2129 VGND VGND VPWR VPWR _10442_ sky130_fd_sc_hd__or4_1
XFILLER_0_153_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length8690 net8691 VGND VGND VPWR VPWR net8690 sky130_fd_sc_hd__buf_1
X_17545_ _09426_ svm0.tC\[13\] _09425_ net6698 VGND VGND VPWR VPWR _09427_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_157_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14757_ net7448 net7153 VGND VGND VPWR VPWR _06888_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13708_ net1562 _05976_ VGND VGND VPWR VPWR _05977_ sky130_fd_sc_hd__xnor2_1
X_17476_ svm0.delta\[6\] _09367_ VGND VGND VPWR VPWR _09368_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14688_ _06826_ _06835_ VGND VGND VPWR VPWR _06836_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_88_Left_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19215_ net3883 _11050_ _11051_ VGND VGND VPWR VPWR _11052_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13639_ net7638 net1982 net2360 VGND VGND VPWR VPWR _05909_ sky130_fd_sc_hd__and3_1
X_16427_ _08480_ _08488_ VGND VGND VPWR VPWR _08489_ sky130_fd_sc_hd__xor2_1
XFILLER_0_116_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19146_ net6299 net6327 VGND VGND VPWR VPWR _10983_ sky130_fd_sc_hd__nand2_2
X_16358_ _08415_ _08420_ VGND VGND VPWR VPWR _08421_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_26_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15309_ net3510 net3505 net4196 net4194 VGND VGND VPWR VPWR _07383_ sky130_fd_sc_hd__o22a_1
XFILLER_0_152_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6481 cordic0.gm0.iter\[2\] VGND VGND VPWR VPWR net6481 sky130_fd_sc_hd__buf_1
X_19077_ net6319 _10845_ _10913_ net6249 VGND VGND VPWR VPWR _10914_ sky130_fd_sc_hd__a211oi_1
X_16289_ _08310_ _08352_ VGND VGND VPWR VPWR _08353_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout6492 net6505 VGND VGND VPWR VPWR net6492 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18028_ net7013 net6936 VGND VGND VPWR VPWR _09879_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_97_Left_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19979_ net1406 _11809_ VGND VGND VPWR VPWR _11810_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_157_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22990_ matmul0.beta_pass\[14\] _08744_ net6575 VGND VGND VPWR VPWR _02863_ sky130_fd_sc_hd__mux2_1
X_21941_ _01847_ _01848_ _01846_ VGND VGND VPWR VPWR _01949_ sky130_fd_sc_hd__o21ba_1
X_24660_ net9228 net1378 _04512_ VGND VGND VPWR VPWR _00682_ sky130_fd_sc_hd__a21o_1
X_21872_ net2066 _01792_ VGND VGND VPWR VPWR _01881_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23611_ _03475_ _03476_ _03477_ VGND VGND VPWR VPWR _03479_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_167_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20823_ _12559_ net2484 VGND VGND VPWR VPWR _00839_ sky130_fd_sc_hd__nor2_1
X_24591_ pid_q.prev_error\[14\] pid_q.curr_error\[14\] VGND VGND VPWR VPWR _04447_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_38_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23542_ _03328_ net2426 _03409_ VGND VGND VPWR VPWR _03410_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8906 net8904 VGND VGND VPWR VPWR net8906 sky130_fd_sc_hd__buf_1
X_20754_ net5579 net5822 _12523_ _12524_ VGND VGND VPWR VPWR _12525_ sky130_fd_sc_hd__a31o_1
Xwire8917 net8918 VGND VGND VPWR VPWR net8917 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8928 net8929 VGND VGND VPWR VPWR net8928 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8939 net102 VGND VGND VPWR VPWR net8939 sky130_fd_sc_hd__clkbuf_1
X_23473_ _03283_ _03284_ _03285_ VGND VGND VPWR VPWR _03342_ sky130_fd_sc_hd__o21a_1
XFILLER_0_190_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20685_ net1403 _12460_ net8061 VGND VGND VPWR VPWR _12461_ sky130_fd_sc_hd__o21ai_1
Xwire607 net608 VGND VGND VPWR VPWR net607 sky130_fd_sc_hd__clkbuf_2
X_25212_ clknet_leaf_61_clk _00101_ net8717 VGND VGND VPWR VPWR svm0.vC\[0\] sky130_fd_sc_hd__dfrtp_1
Xwire618 _09125_ VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__clkbuf_2
Xwire629 net630 VGND VGND VPWR VPWR net629 sky130_fd_sc_hd__buf_1
X_22424_ net5708 _02349_ VGND VGND VPWR VPWR _02426_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25143_ clknet_leaf_48_clk _00032_ net8762 VGND VGND VPWR VPWR svm0.tC\[15\] sky130_fd_sc_hd__dfrtp_1
X_22355_ _02347_ _02357_ VGND VGND VPWR VPWR _02358_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_66_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21306_ net3119 _01319_ _01320_ _00862_ VGND VGND VPWR VPWR _01321_ sky130_fd_sc_hd__o22a_1
X_25074_ _04819_ _04820_ net1994 VGND VGND VPWR VPWR _04821_ sky130_fd_sc_hd__a21oi_1
X_22286_ _02210_ _02211_ _02289_ VGND VGND VPWR VPWR _02290_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_14_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24025_ _03699_ _03887_ VGND VGND VPWR VPWR _03888_ sky130_fd_sc_hd__xor2_2
Xwire3202 net3203 VGND VGND VPWR VPWR net3202 sky130_fd_sc_hd__buf_1
Xhold260 svm0.delta\[15\] VGND VGND VPWR VPWR net9213 sky130_fd_sc_hd__dlygate4sd3_1
X_21237_ _00935_ _01238_ _01239_ _01235_ VGND VGND VPWR VPWR _01252_ sky130_fd_sc_hd__o22a_1
XFILLER_0_130_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold271 pid_d.prev_int\[11\] VGND VGND VPWR VPWR net9224 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3213 _10811_ VGND VGND VPWR VPWR net3213 sky130_fd_sc_hd__buf_1
Xhold282 matmul0.beta_pass\[13\] VGND VGND VPWR VPWR net9235 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3224 _10391_ VGND VGND VPWR VPWR net3224 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3235 net3236 VGND VGND VPWR VPWR net3235 sky130_fd_sc_hd__clkbuf_2
Xwire2501 _11647_ VGND VGND VPWR VPWR net2501 sky130_fd_sc_hd__buf_1
Xwire3246 net3247 VGND VGND VPWR VPWR net3246 sky130_fd_sc_hd__clkbuf_1
Xwire2512 _11131_ VGND VGND VPWR VPWR net2512 sky130_fd_sc_hd__buf_1
Xwire3257 _09643_ VGND VGND VPWR VPWR net3257 sky130_fd_sc_hd__buf_1
X_21168_ net5882 _01182_ _01183_ VGND VGND VPWR VPWR _01184_ sky130_fd_sc_hd__mux2_1
Xwire2523 net2524 VGND VGND VPWR VPWR net2523 sky130_fd_sc_hd__clkbuf_2
Xwire3268 _09600_ VGND VGND VPWR VPWR net3268 sky130_fd_sc_hd__clkbuf_2
Xwire3279 _09258_ VGND VGND VPWR VPWR net3279 sky130_fd_sc_hd__buf_1
Xwire2534 net2535 VGND VGND VPWR VPWR net2534 sky130_fd_sc_hd__clkbuf_1
Xwire1800 _09190_ VGND VGND VPWR VPWR net1800 sky130_fd_sc_hd__clkbuf_2
Xwire2545 _10068_ VGND VGND VPWR VPWR net2545 sky130_fd_sc_hd__buf_1
Xwire1811 net1812 VGND VGND VPWR VPWR net1811 sky130_fd_sc_hd__clkbuf_1
Xwire2556 net2557 VGND VGND VPWR VPWR net2556 sky130_fd_sc_hd__buf_1
X_20119_ _11944_ _11945_ VGND VGND VPWR VPWR _11947_ sky130_fd_sc_hd__nand2_1
Xwire2567 net2570 VGND VGND VPWR VPWR net2567 sky130_fd_sc_hd__buf_1
X_13990_ _06253_ _06254_ VGND VGND VPWR VPWR _06255_ sky130_fd_sc_hd__xnor2_1
Xwire1822 net1823 VGND VGND VPWR VPWR net1822 sky130_fd_sc_hd__buf_1
X_21099_ _01099_ _01112_ _01114_ VGND VGND VPWR VPWR _01115_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_102_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1833 net1834 VGND VGND VPWR VPWR net1833 sky130_fd_sc_hd__buf_1
Xwire2578 _09272_ VGND VGND VPWR VPWR net2578 sky130_fd_sc_hd__buf_1
Xwire2589 _09158_ VGND VGND VPWR VPWR net2589 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1844 _07945_ VGND VGND VPWR VPWR net1844 sky130_fd_sc_hd__clkbuf_1
X_24927_ net8867 net141 VGND VGND VPWR VPWR _04712_ sky130_fd_sc_hd__and2b_1
X_12941_ _05212_ _05213_ VGND VGND VPWR VPWR _05214_ sky130_fd_sc_hd__xnor2_2
Xwire1855 net1856 VGND VGND VPWR VPWR net1855 sky130_fd_sc_hd__clkbuf_1
Xwire1866 net1867 VGND VGND VPWR VPWR net1866 sky130_fd_sc_hd__buf_1
Xwire1877 _07350_ VGND VGND VPWR VPWR net1877 sky130_fd_sc_hd__buf_1
XFILLER_0_88_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1888 _07220_ VGND VGND VPWR VPWR net1888 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15660_ _07730_ _07731_ VGND VGND VPWR VPWR _07732_ sky130_fd_sc_hd__nand2_1
Xwire1899 net1900 VGND VGND VPWR VPWR net1899 sky130_fd_sc_hd__clkbuf_1
X_24858_ _04662_ net4767 net2003 VGND VGND VPWR VPWR _04663_ sky130_fd_sc_hd__mux2_1
X_12872_ _05088_ _05143_ VGND VGND VPWR VPWR _05145_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14611_ net9097 net892 _06655_ _06779_ _06783_ VGND VGND VPWR VPWR _00116_ sky130_fd_sc_hd__a221o_1
XFILLER_0_139_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23809_ pid_q.curr_int\[5\] pid_q.prev_int\[5\] VGND VGND VPWR VPWR _03674_ sky130_fd_sc_hd__xor2_1
X_15591_ net1854 net1853 VGND VGND VPWR VPWR _07663_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_119_clk clknet_4_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_119_clk
+ sky130_fd_sc_hd__clkbuf_16
X_24789_ net5206 net1987 VGND VGND VPWR VPWR _04615_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length7274 matmul0.alpha_pass\[9\] VGND VGND VPWR VPWR net7274 sky130_fd_sc_hd__buf_1
X_17330_ net7890 _09206_ net7862 VGND VGND VPWR VPWR _09244_ sky130_fd_sc_hd__o21ai_1
Xmax_length6540 net6541 VGND VGND VPWR VPWR net6540 sky130_fd_sc_hd__buf_1
X_14542_ net4225 _06714_ _06716_ _06711_ _06720_ VGND VGND VPWR VPWR _06721_ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17261_ net3387 _09187_ _09186_ VGND VGND VPWR VPWR _09192_ sky130_fd_sc_hd__mux2_1
X_14473_ _06657_ _06658_ _06659_ VGND VGND VPWR VPWR _06660_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_165_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19000_ net6342 net6351 VGND VGND VPWR VPWR _10837_ sky130_fd_sc_hd__and2b_1
X_16212_ net3516 net3429 net3424 net3587 VGND VGND VPWR VPWR _08277_ sky130_fd_sc_hd__o211a_1
X_13424_ net843 net842 _05696_ VGND VGND VPWR VPWR _05697_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17192_ _09122_ _09123_ _09133_ net1076 VGND VGND VPWR VPWR _09142_ sky130_fd_sc_hd__o31a_1
XFILLER_0_11_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5021 pid_q.mult0.b\[5\] VGND VGND VPWR VPWR net5021 sky130_fd_sc_hd__buf_1
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16143_ _08207_ _08208_ VGND VGND VPWR VPWR _08209_ sky130_fd_sc_hd__nand2_1
X_13355_ _05511_ net1133 VGND VGND VPWR VPWR _05628_ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout5043 pid_q.mult0.b\[4\] VGND VGND VPWR VPWR net5043 sky130_fd_sc_hd__buf_1
XFILLER_0_178_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout4331 net4334 VGND VGND VPWR VPWR net4331 sky130_fd_sc_hd__clkbuf_2
X_16074_ net2662 _08028_ _08026_ VGND VGND VPWR VPWR _08141_ sky130_fd_sc_hd__o21ai_1
X_13286_ _05464_ _05465_ _05468_ _05467_ VGND VGND VPWR VPWR _05559_ sky130_fd_sc_hd__a211o_1
Xwire5160 net5161 VGND VGND VPWR VPWR net5160 sky130_fd_sc_hd__clkbuf_1
Xwire5171 pid_q.curr_int\[14\] VGND VGND VPWR VPWR net5171 sky130_fd_sc_hd__buf_1
X_19902_ _11661_ _11732_ _11733_ _11670_ VGND VGND VPWR VPWR _11734_ sky130_fd_sc_hd__o22a_1
X_15025_ net4171 net4167 VGND VGND VPWR VPWR _07099_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5193 net5194 VGND VGND VPWR VPWR net5193 sky130_fd_sc_hd__clkbuf_1
Xwire4481 pid_q.ki\[5\] VGND VGND VPWR VPWR net4481 sky130_fd_sc_hd__clkbuf_1
X_19833_ net567 VGND VGND VPWR VPWR _11667_ sky130_fd_sc_hd__buf_2
XFILLER_0_194_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3780 net3781 VGND VGND VPWR VPWR net3780 sky130_fd_sc_hd__buf_1
Xwire3791 net3792 VGND VGND VPWR VPWR net3791 sky130_fd_sc_hd__clkbuf_1
X_19764_ net958 net956 VGND VGND VPWR VPWR _11599_ sky130_fd_sc_hd__or2b_1
X_16976_ _08936_ _08938_ VGND VGND VPWR VPWR _08939_ sky130_fd_sc_hd__and2_1
X_18715_ _10552_ _10560_ VGND VGND VPWR VPWR _10561_ sky130_fd_sc_hd__xnor2_2
Xinput6 angle_in[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
X_15927_ _07987_ _07995_ VGND VGND VPWR VPWR _07996_ sky130_fd_sc_hd__xor2_1
XFILLER_0_127_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19695_ _11529_ _11530_ VGND VGND VPWR VPWR _11531_ sky130_fd_sc_hd__and2b_1
XFILLER_0_160_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18646_ _10464_ _10492_ VGND VGND VPWR VPWR _10493_ sky130_fd_sc_hd__xnor2_2
X_15858_ net2234 net2727 _07837_ VGND VGND VPWR VPWR _07927_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_143_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14809_ net9045 net3005 net2853 _06921_ VGND VGND VPWR VPWR _00176_ sky130_fd_sc_hd__o22a_1
X_18577_ net3308 _10171_ VGND VGND VPWR VPWR _10425_ sky130_fd_sc_hd__nand2_1
XFILLER_0_176_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15789_ _07857_ _07858_ VGND VGND VPWR VPWR _07859_ sky130_fd_sc_hd__or2b_1
XFILLER_0_52_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17528_ net4253 _09411_ net3388 VGND VGND VPWR VPWR _09412_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17459_ svm0.delta\[3\] _09347_ _09348_ svm0.counter\[3\] VGND VGND VPWR VPWR _09353_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_171_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20470_ _12259_ _08900_ net1810 VGND VGND VPWR VPWR _12261_ sky130_fd_sc_hd__and3b_1
XFILLER_0_144_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19129_ _10936_ _10965_ VGND VGND VPWR VPWR _10966_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_112_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22140_ _02135_ _02145_ VGND VGND VPWR VPWR _02146_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_164_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22071_ _01959_ net1713 _02077_ VGND VGND VPWR VPWR _02078_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_168_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21022_ net5622 net5868 VGND VGND VPWR VPWR _01038_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25830_ clknet_leaf_37_clk _00703_ net8680 VGND VGND VPWR VPWR pid_q.curr_error\[6\]
+ sky130_fd_sc_hd__dfrtp_2
Xwire1107 _07703_ VGND VGND VPWR VPWR net1107 sky130_fd_sc_hd__clkbuf_1
Xwire1118 _06857_ VGND VGND VPWR VPWR net1118 sky130_fd_sc_hd__clkbuf_1
Xwire1129 _05706_ VGND VGND VPWR VPWR net1129 sky130_fd_sc_hd__buf_1
X_25761_ clknet_leaf_95_clk _00634_ net8455 VGND VGND VPWR VPWR pid_d.out\[2\] sky130_fd_sc_hd__dfrtp_1
X_22973_ _02854_ VGND VGND VPWR VPWR _00653_ sky130_fd_sc_hd__clkbuf_1
X_24712_ net1621 _04547_ VGND VGND VPWR VPWR _04548_ sky130_fd_sc_hd__nand2_1
X_21924_ _01928_ _01931_ VGND VGND VPWR VPWR _01932_ sky130_fd_sc_hd__xnor2_1
X_25692_ clknet_leaf_6_clk _00565_ net8562 VGND VGND VPWR VPWR pid_d.curr_error\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_182_Right_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24643_ _04441_ net631 VGND VGND VPWR VPWR _04498_ sky130_fd_sc_hd__nor2_1
X_21855_ net5406 net5857 VGND VGND VPWR VPWR _01864_ sky130_fd_sc_hd__and2b_1
Xfanout8608 net8639 VGND VGND VPWR VPWR net8608 sky130_fd_sc_hd__clkbuf_2
Xmax_length5102 net5091 VGND VGND VPWR VPWR net5102 sky130_fd_sc_hd__buf_1
XFILLER_0_33_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20806_ _00820_ _00821_ VGND VGND VPWR VPWR _00822_ sky130_fd_sc_hd__xnor2_1
X_24574_ _04428_ _04429_ VGND VGND VPWR VPWR _04430_ sky130_fd_sc_hd__xor2_1
X_21786_ _01593_ VGND VGND VPWR VPWR _01796_ sky130_fd_sc_hd__buf_1
XFILLER_0_136_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8703 net8704 VGND VGND VPWR VPWR net8703 sky130_fd_sc_hd__buf_1
XFILLER_0_154_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout7918 net7929 VGND VGND VPWR VPWR net7918 sky130_fd_sc_hd__buf_1
XFILLER_0_108_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8714 net8715 VGND VGND VPWR VPWR net8714 sky130_fd_sc_hd__buf_1
X_23525_ _03391_ _03392_ VGND VGND VPWR VPWR _03393_ sky130_fd_sc_hd__xnor2_1
Xwire8725 net8726 VGND VGND VPWR VPWR net8725 sky130_fd_sc_hd__clkbuf_1
Xwire8736 net8737 VGND VGND VPWR VPWR net8736 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20737_ _12504_ _12507_ VGND VGND VPWR VPWR _12508_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire404 _06002_ VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__clkbuf_2
Xwire8758 net8759 VGND VGND VPWR VPWR net8758 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire415 net416 VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__clkbuf_1
X_23456_ _03323_ _03324_ VGND VGND VPWR VPWR _03325_ sky130_fd_sc_hd__xnor2_1
Xwire426 net427 VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__buf_1
XFILLER_0_190_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20668_ _12443_ _12444_ VGND VGND VPWR VPWR _12445_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire437 net438 VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__clkbuf_1
Xwire448 _06736_ VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__clkbuf_1
Xwire459 _04603_ VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__clkbuf_1
X_22407_ net549 VGND VGND VPWR VPWR _02409_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23387_ _03223_ net2428 _03221_ VGND VGND VPWR VPWR _03257_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_34_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20599_ net6239 _12371_ _12370_ VGND VGND VPWR VPWR _12381_ sky130_fd_sc_hd__a21o_1
XFILLER_0_150_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13140_ net7821 net2966 net2305 VGND VGND VPWR VPWR _05413_ sky130_fd_sc_hd__and3_1
X_25126_ pid_d.prev_int\[14\] _04849_ net2391 pid_d.curr_int\[14\] VGND VGND VPWR
+ VPWR _00807_ sky130_fd_sc_hd__a22o_1
X_22338_ _02304_ _02309_ _02340_ VGND VGND VPWR VPWR _02341_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_103_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13071_ net6677 net5204 net6673 VGND VGND VPWR VPWR _05344_ sky130_fd_sc_hd__and3b_1
X_25057_ net3737 net685 _04805_ VGND VGND VPWR VPWR _04806_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22269_ pid_d.curr_int\[12\] net4391 VGND VGND VPWR VPWR _02273_ sky130_fd_sc_hd__xor2_1
XFILLER_0_20_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3010 net3011 VGND VGND VPWR VPWR net3010 sky130_fd_sc_hd__buf_1
Xwire3021 net3027 VGND VGND VPWR VPWR net3021 sky130_fd_sc_hd__buf_1
X_24008_ _03703_ _03821_ VGND VGND VPWR VPWR _03871_ sky130_fd_sc_hd__or2b_1
Xwire3032 _04857_ VGND VGND VPWR VPWR net3032 sky130_fd_sc_hd__buf_1
Xwire3043 net3048 VGND VGND VPWR VPWR net3043 sky130_fd_sc_hd__clkbuf_1
Xwire3054 net3055 VGND VGND VPWR VPWR net3054 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2320 _04975_ VGND VGND VPWR VPWR net2320 sky130_fd_sc_hd__buf_1
Xwire3065 net3066 VGND VGND VPWR VPWR net3065 sky130_fd_sc_hd__buf_1
Xwire3076 net3077 VGND VGND VPWR VPWR net3076 sky130_fd_sc_hd__buf_1
Xwire2342 net2343 VGND VGND VPWR VPWR net2342 sky130_fd_sc_hd__buf_1
X_16830_ net6428 matmul0.sin\[3\] net3365 VGND VGND VPWR VPWR _08806_ sky130_fd_sc_hd__mux2_1
Xwire3087 net3088 VGND VGND VPWR VPWR net3087 sky130_fd_sc_hd__buf_1
Xwire3098 net3099 VGND VGND VPWR VPWR net3098 sky130_fd_sc_hd__buf_1
Xwire2353 _04917_ VGND VGND VPWR VPWR net2353 sky130_fd_sc_hd__buf_1
Xwire2364 _04907_ VGND VGND VPWR VPWR net2364 sky130_fd_sc_hd__buf_1
Xwire2375 net2376 VGND VGND VPWR VPWR net2375 sky130_fd_sc_hd__buf_1
Xwire1630 _04780_ VGND VGND VPWR VPWR net1630 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1641 _04554_ VGND VGND VPWR VPWR net1641 sky130_fd_sc_hd__clkbuf_1
Xwire2386 net2387 VGND VGND VPWR VPWR net2386 sky130_fd_sc_hd__clkbuf_1
X_13973_ net1965 net1583 _06235_ _06237_ net7633 VGND VGND VPWR VPWR _06238_ sky130_fd_sc_hd__a32o_1
Xwire1652 _04219_ VGND VGND VPWR VPWR net1652 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_73_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16761_ _08769_ VGND VGND VPWR VPWR _00280_ sky130_fd_sc_hd__clkbuf_1
Xwire2397 net2398 VGND VGND VPWR VPWR net2397 sky130_fd_sc_hd__clkbuf_2
Xwire1663 net1664 VGND VGND VPWR VPWR net1663 sky130_fd_sc_hd__clkbuf_1
Xwire1674 _03214_ VGND VGND VPWR VPWR net1674 sky130_fd_sc_hd__buf_1
XFILLER_0_38_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18500_ net6809 _09177_ VGND VGND VPWR VPWR _10349_ sky130_fd_sc_hd__nor2_2
Xwire1685 net1686 VGND VGND VPWR VPWR net1685 sky130_fd_sc_hd__clkbuf_1
X_12924_ _05194_ _05195_ _05108_ _05109_ VGND VGND VPWR VPWR _05197_ sky130_fd_sc_hd__o22a_1
X_15712_ _07778_ _07782_ VGND VGND VPWR VPWR _07783_ sky130_fd_sc_hd__xnor2_2
Xwire1696 _02662_ VGND VGND VPWR VPWR net1696 sky130_fd_sc_hd__buf_1
X_19480_ _10851_ _11264_ net3196 _11122_ VGND VGND VPWR VPWR _11317_ sky130_fd_sc_hd__a211o_1
X_16692_ matmul0.matmul_stage_inst.mult1\[10\] VGND VGND VPWR VPWR _08722_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18431_ _10277_ _10280_ VGND VGND VPWR VPWR _10281_ sky130_fd_sc_hd__xnor2_1
X_12855_ net3693 _05127_ VGND VGND VPWR VPWR _05128_ sky130_fd_sc_hd__nand2_1
X_15643_ _07714_ VGND VGND VPWR VPWR _07715_ sky130_fd_sc_hd__clkbuf_1
Xmax_length7071 net7072 VGND VGND VPWR VPWR net7071 sky130_fd_sc_hd__clkbuf_2
X_15574_ _07629_ _07630_ VGND VGND VPWR VPWR _07646_ sky130_fd_sc_hd__nor2_1
X_18362_ net6789 _10207_ VGND VGND VPWR VPWR _10213_ sky130_fd_sc_hd__nor2_1
XFILLER_0_185_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12786_ net7284 _04892_ _04894_ _05021_ VGND VGND VPWR VPWR _05059_ sky130_fd_sc_hd__a31oi_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17313_ net6711 _09226_ VGND VGND VPWR VPWR _09227_ sky130_fd_sc_hd__nand2_1
X_14525_ _06703_ _06704_ VGND VGND VPWR VPWR _06705_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18293_ net1215 net1447 VGND VGND VPWR VPWR _10144_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17244_ net2165 net325 net1800 net9155 VGND VGND VPWR VPWR _00342_ sky130_fd_sc_hd__a22o_1
X_14456_ _06541_ VGND VGND VPWR VPWR _06646_ sky130_fd_sc_hd__inv_2
X_13407_ _05482_ _05677_ _05678_ _05679_ VGND VGND VPWR VPWR _05680_ sky130_fd_sc_hd__a31o_1
XFILLER_0_114_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17175_ net6901 _09102_ net527 _09126_ VGND VGND VPWR VPWR _09127_ sky130_fd_sc_hd__a211o_1
X_14387_ _06593_ VGND VGND VPWR VPWR _00082_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire960 _11304_ VGND VGND VPWR VPWR net960 sky130_fd_sc_hd__clkbuf_1
Xwire971 _08993_ VGND VGND VPWR VPWR net971 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16126_ _08121_ _08122_ _08123_ VGND VGND VPWR VPWR _08192_ sky130_fd_sc_hd__a21o_1
Xwire982 _08266_ VGND VGND VPWR VPWR net982 sky130_fd_sc_hd__clkbuf_1
X_13338_ _05607_ _05610_ VGND VGND VPWR VPWR _05611_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire993 _06910_ VGND VGND VPWR VPWR net993 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16057_ _08122_ _08123_ VGND VGND VPWR VPWR _08124_ sky130_fd_sc_hd__xnor2_1
X_13269_ _05539_ _05540_ _05423_ VGND VGND VPWR VPWR _05542_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15008_ _07076_ _07079_ _07081_ VGND VGND VPWR VPWR _07082_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19816_ net6010 _11649_ VGND VGND VPWR VPWR _11650_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19747_ net6219 net6131 VGND VGND VPWR VPWR _11582_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_2_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16959_ net7129 _08920_ _08921_ net7147 VGND VGND VPWR VPWR _08922_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19678_ net6220 _11513_ net3162 VGND VGND VPWR VPWR _11514_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18629_ _10474_ _10475_ VGND VGND VPWR VPWR _10476_ sky130_fd_sc_hd__xor2_1
XFILLER_0_52_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21640_ _01554_ _01615_ VGND VGND VPWR VPWR _01651_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21571_ net1722 _01582_ VGND VGND VPWR VPWR _01583_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7309 net7310 VGND VGND VPWR VPWR net7309 sky130_fd_sc_hd__buf_1
X_23310_ _02965_ _02988_ _03178_ _03179_ VGND VGND VPWR VPWR _03180_ sky130_fd_sc_hd__a2bb2o_1
X_20522_ _12306_ _12307_ _12308_ net6324 VGND VGND VPWR VPWR _00503_ sky130_fd_sc_hd__o22a_1
X_24290_ net2024 net1653 VGND VGND VPWR VPWR _04150_ sky130_fd_sc_hd__xor2_2
XFILLER_0_28_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6608 matmul0.done_pass VGND VGND VPWR VPWR net6608 sky130_fd_sc_hd__buf_1
Xwire6619 net6620 VGND VGND VPWR VPWR net6619 sky130_fd_sc_hd__buf_1
X_23241_ net3060 _03110_ VGND VGND VPWR VPWR _03111_ sky130_fd_sc_hd__xnor2_1
X_20453_ _12244_ net809 VGND VGND VPWR VPWR _12246_ sky130_fd_sc_hd__xor2_1
XFILLER_0_104_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5907 net5908 VGND VGND VPWR VPWR net5907 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5918 net5919 VGND VGND VPWR VPWR net5918 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5929 net5930 VGND VGND VPWR VPWR net5929 sky130_fd_sc_hd__dlymetal6s2s_1
X_23172_ _03040_ _03041_ VGND VGND VPWR VPWR _03042_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20384_ net6374 _12159_ VGND VGND VPWR VPWR _12183_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_179_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22123_ net5708 net5464 VGND VGND VPWR VPWR _02129_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput151 net6683 VGND VGND VPWR VPWR pwmC_out sky130_fd_sc_hd__clkbuf_4
X_22054_ _02057_ _02059_ VGND VGND VPWR VPWR _02061_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21005_ _01011_ net1183 VGND VGND VPWR VPWR _01021_ sky130_fd_sc_hd__xnor2_1
X_25813_ clknet_leaf_36_clk _00686_ net8748 VGND VGND VPWR VPWR pid_q.prev_error\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_25744_ clknet_leaf_8_clk _00617_ net8554 VGND VGND VPWR VPWR pid_d.kp\[2\] sky130_fd_sc_hd__dfrtp_1
X_22956_ pid_d.out\[14\] pid_d.curr_int\[14\] VGND VGND VPWR VPWR _02844_ sky130_fd_sc_hd__nand2_1
XFILLER_0_186_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21907_ net9022 net3123 net2078 _01915_ VGND VGND VPWR VPWR _00526_ sky130_fd_sc_hd__a22o_1
X_25675_ clknet_leaf_4_clk _00548_ net8561 VGND VGND VPWR VPWR pid_d.prev_error\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_22887_ net5357 net3103 _02781_ net4338 VGND VGND VPWR VPWR _02782_ sky130_fd_sc_hd__a22o_1
X_24626_ net4823 net3745 net4807 _04475_ VGND VGND VPWR VPWR _04481_ sky130_fd_sc_hd__a211o_1
X_12640_ net2354 VGND VGND VPWR VPWR _04913_ sky130_fd_sc_hd__clkbuf_1
Xfanout8405 net8410 VGND VGND VPWR VPWR net8405 sky130_fd_sc_hd__clkbuf_2
X_21838_ net5801 net5408 VGND VGND VPWR VPWR _01847_ sky130_fd_sc_hd__nand2_1
XFILLER_0_183_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout8438 net8441 VGND VGND VPWR VPWR net8438 sky130_fd_sc_hd__buf_1
Xwire8500 net8499 VGND VGND VPWR VPWR net8500 sky130_fd_sc_hd__clkbuf_2
X_24557_ _04342_ _04353_ net1649 VGND VGND VPWR VPWR _04413_ sky130_fd_sc_hd__a21bo_1
X_12571_ net9150 _04854_ net1622 VGND VGND VPWR VPWR _00013_ sky130_fd_sc_hd__a21o_1
Xwire8511 net8512 VGND VGND VPWR VPWR net8511 sky130_fd_sc_hd__clkbuf_2
X_21769_ _01778_ VGND VGND VPWR VPWR _01779_ sky130_fd_sc_hd__buf_1
Xwire8522 net8523 VGND VGND VPWR VPWR net8522 sky130_fd_sc_hd__buf_1
XFILLER_0_194_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_50_clk clknet_4_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8533 net8534 VGND VGND VPWR VPWR net8533 sky130_fd_sc_hd__clkbuf_1
X_14310_ net6750 net6604 VGND VGND VPWR VPWR _06532_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length4231 _06708_ VGND VGND VPWR VPWR net4231 sky130_fd_sc_hd__clkbuf_1
Xwire8544 net8545 VGND VGND VPWR VPWR net8544 sky130_fd_sc_hd__clkbuf_1
X_23508_ _03370_ net1024 VGND VGND VPWR VPWR _03377_ sky130_fd_sc_hd__or2_1
Xwire7810 net7811 VGND VGND VPWR VPWR net7810 sky130_fd_sc_hd__buf_1
XFILLER_0_53_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7821 net7822 VGND VGND VPWR VPWR net7821 sky130_fd_sc_hd__buf_1
Xwire201 net202 VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_1
X_15290_ net1542 net1875 VGND VGND VPWR VPWR _07364_ sky130_fd_sc_hd__xnor2_1
X_24488_ net4848 net4505 VGND VGND VPWR VPWR _04345_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire212 net213 VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_1
Xwire223 net224 VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__buf_1
Xmax_length4264 _04973_ VGND VGND VPWR VPWR net4264 sky130_fd_sc_hd__clkbuf_1
Xwire7832 net7833 VGND VGND VPWR VPWR net7832 sky130_fd_sc_hd__buf_1
Xwire234 _04445_ VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__buf_1
Xwire8588 net8589 VGND VGND VPWR VPWR net8588 sky130_fd_sc_hd__buf_1
Xwire7854 net7855 VGND VGND VPWR VPWR net7854 sky130_fd_sc_hd__buf_1
Xwire8599 net8600 VGND VGND VPWR VPWR net8599 sky130_fd_sc_hd__clkbuf_1
X_14241_ net6456 net6446 net8319 VGND VGND VPWR VPWR _06497_ sky130_fd_sc_hd__or3b_1
Xwire245 _10766_ VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__buf_1
X_23439_ _03307_ net646 net640 VGND VGND VPWR VPWR _03309_ sky130_fd_sc_hd__and3_1
Xwire256 net257 VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__buf_1
Xwire7876 net7877 VGND VGND VPWR VPWR net7876 sky130_fd_sc_hd__buf_1
Xwire267 net268 VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__clkbuf_1
Xwire7887 net7880 VGND VGND VPWR VPWR net7887 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire278 net279 VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__clkbuf_1
Xwire289 _05856_ VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7898 net7888 VGND VGND VPWR VPWR net7898 sky130_fd_sc_hd__buf_1
X_14172_ net217 net403 _06368_ _06369_ VGND VGND VPWR VPWR _06432_ sky130_fd_sc_hd__a211o_1
Xmax_length3596 net3597 VGND VGND VPWR VPWR net3596 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13123_ _05382_ net849 VGND VGND VPWR VPWR _05396_ sky130_fd_sc_hd__xnor2_1
X_25109_ net8902 net4300 net4332 net3762 VGND VGND VPWR VPWR _04851_ sky130_fd_sc_hd__and4_1
X_18980_ net6356 net2529 VGND VGND VPWR VPWR _10817_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13054_ _05325_ net1155 _05326_ _05030_ VGND VGND VPWR VPWR _05327_ sky130_fd_sc_hd__o2bb2a_1
X_17931_ _09678_ _09780_ _09781_ VGND VGND VPWR VPWR _09782_ sky130_fd_sc_hd__o21ai_1
X_17862_ net3998 _09708_ _09710_ _09712_ VGND VGND VPWR VPWR _09713_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2150 _09577_ VGND VGND VPWR VPWR net2150 sky130_fd_sc_hd__clkbuf_1
Xwire2161 net2163 VGND VGND VPWR VPWR net2161 sky130_fd_sc_hd__buf_1
X_19601_ _11434_ _11435_ _11437_ VGND VGND VPWR VPWR _11438_ sky130_fd_sc_hd__and3_1
X_16813_ net8972 matmul0.cos\[9\] net3367 VGND VGND VPWR VPWR _08797_ sky130_fd_sc_hd__mux2_1
Xwire2172 _08989_ VGND VGND VPWR VPWR net2172 sky130_fd_sc_hd__buf_1
Xwire2183 net2184 VGND VGND VPWR VPWR net2183 sky130_fd_sc_hd__buf_1
X_17793_ net7108 net7136 VGND VGND VPWR VPWR _09644_ sky130_fd_sc_hd__nand2b_1
Xwire2194 _08818_ VGND VGND VPWR VPWR net2194 sky130_fd_sc_hd__clkbuf_1
Xwire1460 _09455_ VGND VGND VPWR VPWR net1460 sky130_fd_sc_hd__clkbuf_1
Xwire1471 net1472 VGND VGND VPWR VPWR net1471 sky130_fd_sc_hd__buf_1
X_19532_ _11300_ _11307_ _11306_ VGND VGND VPWR VPWR _11369_ sky130_fd_sc_hd__a21bo_1
X_16744_ matmul0.b_in\[8\] matmul0.b\[8\] net3381 VGND VGND VPWR VPWR _08761_ sky130_fd_sc_hd__mux2_1
X_13956_ _05191_ VGND VGND VPWR VPWR _06221_ sky130_fd_sc_hd__buf_2
Xwire1482 _08990_ VGND VGND VPWR VPWR net1482 sky130_fd_sc_hd__buf_1
XFILLER_0_191_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12907_ _05178_ _05179_ VGND VGND VPWR VPWR _05180_ sky130_fd_sc_hd__xor2_1
X_19463_ _11286_ _11299_ VGND VGND VPWR VPWR _11300_ sky130_fd_sc_hd__xnor2_1
X_13887_ _06081_ _06143_ VGND VGND VPWR VPWR _06153_ sky130_fd_sc_hd__or2_1
X_16675_ _08706_ _08707_ VGND VGND VPWR VPWR _08708_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_186_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18414_ net2135 VGND VGND VPWR VPWR _10264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12838_ net1956 VGND VGND VPWR VPWR _05111_ sky130_fd_sc_hd__clkbuf_2
X_15626_ net3597 net3591 net4083 net4081 VGND VGND VPWR VPWR _07698_ sky130_fd_sc_hd__o22a_1
X_19394_ net1061 _11230_ VGND VGND VPWR VPWR _11231_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_189_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18345_ _10192_ _10195_ VGND VGND VPWR VPWR _10196_ sky130_fd_sc_hd__and2_1
X_12769_ _05040_ _05041_ VGND VGND VPWR VPWR _05042_ sky130_fd_sc_hd__xor2_1
X_15557_ net2703 net3407 VGND VGND VPWR VPWR _07630_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_41_clk clknet_4_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_185_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14508_ _06685_ _06688_ VGND VGND VPWR VPWR _06690_ sky130_fd_sc_hd__or2_1
X_18276_ _10115_ _10116_ _10126_ VGND VGND VPWR VPWR _10127_ sky130_fd_sc_hd__nand3_1
X_15488_ _07561_ VGND VGND VPWR VPWR _00215_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput20 currA_in[12] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
X_17227_ net6791 net966 _09163_ _09165_ VGND VGND VPWR VPWR _09175_ sky130_fd_sc_hd__and4_1
X_14439_ _06633_ VGND VGND VPWR VPWR _00094_ sky130_fd_sc_hd__clkbuf_1
Xinput31 currA_in[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput42 currB_in[3] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_1
Xinput53 currT_in[13] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_1
Xinput64 currT_in[9] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_1
Xinput75 periodTop[4] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_1
Xwire790 _05205_ VGND VGND VPWR VPWR net790 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17158_ net4039 net4058 net3305 _09110_ VGND VGND VPWR VPWR _09111_ sky130_fd_sc_hd__a31o_1
Xinput86 pid_d_addr[14] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_1
Xinput97 pid_d_data[0] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16109_ _08170_ _08174_ VGND VGND VPWR VPWR _08175_ sky130_fd_sc_hd__xnor2_1
X_17089_ _09039_ net772 VGND VGND VPWR VPWR _09047_ sky130_fd_sc_hd__xor2_1
XFILLER_0_161_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22810_ net8895 _02713_ VGND VGND VPWR VPWR _02714_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23790_ _03652_ _03655_ VGND VGND VPWR VPWR _03656_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_165_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22741_ net3719 net108 VGND VGND VPWR VPWR _02672_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25460_ clknet_leaf_66_clk net8977 net8647 VGND VGND VPWR VPWR matmul0.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_22672_ _02622_ net5630 net2448 VGND VGND VPWR VPWR _02623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24411_ _04222_ _04225_ _04221_ VGND VGND VPWR VPWR _04269_ sky130_fd_sc_hd__a21o_1
X_21623_ net600 _01634_ VGND VGND VPWR VPWR _01635_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25391_ clknet_leaf_79_clk _00274_ net8493 VGND VGND VPWR VPWR matmul0.b\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_176_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_32_clk clknet_4_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_8_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24342_ net4522 net4873 VGND VGND VPWR VPWR _04201_ sky130_fd_sc_hd__nand2_1
X_21554_ _01562_ _01565_ VGND VGND VPWR VPWR _01566_ sky130_fd_sc_hd__xnor2_2
Xwire7117 net7114 VGND VGND VPWR VPWR net7117 sky130_fd_sc_hd__buf_1
XFILLER_0_30_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7128 net7125 VGND VGND VPWR VPWR net7128 sky130_fd_sc_hd__buf_1
Xwire6405 net6406 VGND VGND VPWR VPWR net6405 sky130_fd_sc_hd__clkbuf_1
X_20505_ net6350 _12282_ _12288_ _12289_ _12291_ VGND VGND VPWR VPWR _12292_ sky130_fd_sc_hd__o311a_1
X_24273_ net4536 net4862 VGND VGND VPWR VPWR _04133_ sky130_fd_sc_hd__nand2_1
Xwire6416 net6417 VGND VGND VPWR VPWR net6416 sky130_fd_sc_hd__buf_1
Xwire6427 cordic0.sin\[4\] VGND VGND VPWR VPWR net6427 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21485_ _01379_ _01384_ _01377_ VGND VGND VPWR VPWR _01498_ sky130_fd_sc_hd__o21a_1
Xwire6438 net6439 VGND VGND VPWR VPWR net6438 sky130_fd_sc_hd__clkbuf_1
Xwire5704 net5701 VGND VGND VPWR VPWR net5704 sky130_fd_sc_hd__buf_1
Xwire6449 net6447 VGND VGND VPWR VPWR net6449 sky130_fd_sc_hd__buf_1
X_23224_ net5063 net4696 VGND VGND VPWR VPWR _03094_ sky130_fd_sc_hd__nand2_1
Xwire5715 net5716 VGND VGND VPWR VPWR net5715 sky130_fd_sc_hd__buf_1
Xwire5726 net5727 VGND VGND VPWR VPWR net5726 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20436_ cordic0.slte0.opA\[12\] net2279 _12229_ VGND VGND VPWR VPWR _12231_ sky130_fd_sc_hd__or3_1
Xwire5737 net5738 VGND VGND VPWR VPWR net5737 sky130_fd_sc_hd__clkbuf_1
Xwire5748 net5749 VGND VGND VPWR VPWR net5748 sky130_fd_sc_hd__clkbuf_1
Xmax_length1446 _10261_ VGND VGND VPWR VPWR net1446 sky130_fd_sc_hd__buf_1
X_23155_ _03019_ _03024_ VGND VGND VPWR VPWR _03025_ sky130_fd_sc_hd__xnor2_1
X_20367_ _08836_ _12157_ net3314 VGND VGND VPWR VPWR _12167_ sky130_fd_sc_hd__mux2_1
Xmax_length1479 net1480 VGND VGND VPWR VPWR net1479 sky130_fd_sc_hd__buf_1
X_22106_ pid_d.curr_int\[10\] pid_d.prev_int\[10\] VGND VGND VPWR VPWR _02112_ sky130_fd_sc_hd__xor2_1
X_23086_ net5069 net4629 _02954_ _02955_ VGND VGND VPWR VPWR _02956_ sky130_fd_sc_hd__a31o_1
X_20298_ net1471 _12103_ net3317 VGND VGND VPWR VPWR _12104_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_99_clk clknet_4_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_99_clk sky130_fd_sc_hd__clkbuf_16
X_22037_ _01933_ _01935_ _01934_ VGND VGND VPWR VPWR _02044_ sky130_fd_sc_hd__o21a_1
XFILLER_0_101_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_42_Left_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13810_ net780 _05987_ _05988_ VGND VGND VPWR VPWR _06078_ sky130_fd_sc_hd__a21bo_1
X_14790_ _06818_ net7457 VGND VGND VPWR VPWR _06911_ sky130_fd_sc_hd__nand2_1
X_23988_ pid_q.curr_error\[5\] VGND VGND VPWR VPWR _03852_ sky130_fd_sc_hd__inv_2
X_13741_ net322 _06005_ _06008_ _06009_ VGND VGND VPWR VPWR _06010_ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22939_ pid_d.out\[14\] net3104 VGND VGND VPWR VPWR _02828_ sky130_fd_sc_hd__nor2_1
X_25727_ clknet_leaf_8_clk _00600_ net8553 VGND VGND VPWR VPWR pid_d.ki\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_196_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13672_ _05939_ _05940_ VGND VGND VPWR VPWR _05941_ sky130_fd_sc_hd__xor2_2
X_16460_ _08446_ net975 VGND VGND VPWR VPWR _08521_ sky130_fd_sc_hd__xnor2_1
X_25658_ clknet_leaf_3_clk _00531_ net8580 VGND VGND VPWR VPWR pid_d.curr_int\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12623_ net6664 net6678 net6673 VGND VGND VPWR VPWR _04896_ sky130_fd_sc_hd__nor3b_1
X_15411_ net4087 net4086 VGND VGND VPWR VPWR _07485_ sky130_fd_sc_hd__nor2_1
Xfanout7501 net7507 VGND VGND VPWR VPWR net7501 sky130_fd_sc_hd__buf_1
X_24609_ _04423_ _04463_ _04460_ VGND VGND VPWR VPWR _04464_ sky130_fd_sc_hd__o21a_1
X_16391_ _08448_ _08452_ VGND VGND VPWR VPWR _08453_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_39_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_51_Left_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25589_ clknet_leaf_99_clk _00462_ net8382 VGND VGND VPWR VPWR cordic0.cos\[9\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_23_clk clknet_4_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8330 net8331 VGND VGND VPWR VPWR net8330 sky130_fd_sc_hd__clkbuf_1
X_18130_ net7033 _09979_ _09980_ _09623_ net3976 VGND VGND VPWR VPWR _09981_ sky130_fd_sc_hd__o32a_1
X_15342_ net2236 net2796 net2756 net3497 VGND VGND VPWR VPWR _07416_ sky130_fd_sc_hd__a211o_1
XFILLER_0_93_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8352 net8348 VGND VGND VPWR VPWR net8352 sky130_fd_sc_hd__buf_1
XFILLER_0_81_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8363 net8364 VGND VGND VPWR VPWR net8363 sky130_fd_sc_hd__clkbuf_1
Xwire8374 net8375 VGND VGND VPWR VPWR net8374 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7640 net7634 VGND VGND VPWR VPWR net7640 sky130_fd_sc_hd__buf_1
X_18061_ net3330 _09911_ VGND VGND VPWR VPWR _09912_ sky130_fd_sc_hd__xnor2_1
X_15273_ net3559 net3482 VGND VGND VPWR VPWR _07347_ sky130_fd_sc_hd__nor2_1
Xwire7651 net7652 VGND VGND VPWR VPWR net7651 sky130_fd_sc_hd__clkbuf_1
Xwire8396 net8397 VGND VGND VPWR VPWR net8396 sky130_fd_sc_hd__buf_1
Xfanout6866 net6870 VGND VGND VPWR VPWR net6866 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14224_ net7629 net1304 _06470_ VGND VGND VPWR VPWR _06482_ sky130_fd_sc_hd__and3_1
X_17012_ net6465 net4052 VGND VGND VPWR VPWR _08973_ sky130_fd_sc_hd__or2_1
XFILLER_0_184_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6972 net6970 VGND VGND VPWR VPWR net6972 sky130_fd_sc_hd__buf_1
Xwire6983 net6981 VGND VGND VPWR VPWR net6983 sky130_fd_sc_hd__buf_1
X_14155_ net7662 _06374_ _06414_ VGND VGND VPWR VPWR _06416_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length2692 net2693 VGND VGND VPWR VPWR net2692 sky130_fd_sc_hd__buf_1
XFILLER_0_22_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13106_ _05370_ _05378_ VGND VGND VPWR VPWR _05379_ sky130_fd_sc_hd__xnor2_1
Xmax_length1980 _04913_ VGND VGND VPWR VPWR net1980 sky130_fd_sc_hd__clkbuf_1
X_14086_ _06346_ _06348_ VGND VGND VPWR VPWR _06349_ sky130_fd_sc_hd__nand2_2
Xmax_length1991 _04859_ VGND VGND VPWR VPWR net1991 sky130_fd_sc_hd__clkbuf_1
X_18963_ net6268 VGND VGND VPWR VPWR _10800_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_60_Left_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13037_ _05308_ _05309_ net684 VGND VGND VPWR VPWR _05310_ sky130_fd_sc_hd__a21bo_1
X_17914_ net3260 net3259 net2563 VGND VGND VPWR VPWR _09765_ sky130_fd_sc_hd__and3_1
X_18894_ _10680_ _10733_ _10734_ VGND VGND VPWR VPWR _10735_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17845_ net7094 net7068 VGND VGND VPWR VPWR _09696_ sky130_fd_sc_hd__nor2b_1
X_17776_ net7089 _09616_ _09621_ net7061 _09626_ VGND VGND VPWR VPWR _09627_ sky130_fd_sc_hd__o221a_1
X_14988_ net4206 net4202 VGND VGND VPWR VPWR _07062_ sky130_fd_sc_hd__nor2_1
Xwire1290 net1291 VGND VGND VPWR VPWR net1290 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19515_ _11342_ _11351_ VGND VGND VPWR VPWR _11352_ sky130_fd_sc_hd__xnor2_1
X_16727_ net7575 matmul0.b\[0\] net3702 VGND VGND VPWR VPWR _08752_ sky130_fd_sc_hd__mux2_1
X_13939_ _06172_ net677 VGND VGND VPWR VPWR _06205_ sky130_fd_sc_hd__xnor2_1
X_19446_ _11280_ _11281_ _11266_ VGND VGND VPWR VPWR _11283_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16658_ _08692_ _08688_ matmul0.matmul_stage_inst.mult2\[5\] VGND VGND VPWR VPWR
+ _08693_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_174_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15609_ matmul0.matmul_stage_inst.e\[15\] _07151_ _07152_ net7378 VGND VGND VPWR
+ VPWR _07681_ sky130_fd_sc_hd__a22oi_1
X_19377_ net3166 net6152 _11207_ VGND VGND VPWR VPWR _11214_ sky130_fd_sc_hd__or3b_1
XFILLER_0_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16589_ matmul0.matmul_stage_inst.mult2\[5\] net389 net2617 VGND VGND VPWR VPWR _08642_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_14_clk clknet_4_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_162_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18328_ _10172_ _10178_ VGND VGND VPWR VPWR _10179_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_84_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18259_ net3996 net3972 _10109_ VGND VGND VPWR VPWR _10110_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_163_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21270_ _00840_ _00841_ _00842_ VGND VGND VPWR VPWR _01285_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20221_ _12041_ cordic0.slte0.opB\[4\] net2937 VGND VGND VPWR VPWR _12042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20152_ net1055 _11953_ VGND VGND VPWR VPWR _11979_ sky130_fd_sc_hd__nand2_1
Xwire2908 net2909 VGND VGND VPWR VPWR net2908 sky130_fd_sc_hd__clkbuf_1
Xwire2919 net2920 VGND VGND VPWR VPWR net2919 sky130_fd_sc_hd__clkbuf_1
X_24960_ _04699_ net114 net3730 net2011 VGND VGND VPWR VPWR _04734_ sky130_fd_sc_hd__a2bb2o_1
X_20083_ _11911_ VGND VGND VPWR VPWR _11912_ sky130_fd_sc_hd__inv_2
XFILLER_0_176_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23911_ _03773_ _03774_ VGND VGND VPWR VPWR _03775_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24891_ _04685_ VGND VGND VPWR VPWR _00740_ sky130_fd_sc_hd__clkbuf_1
X_23842_ _03700_ _03706_ VGND VGND VPWR VPWR _03707_ sky130_fd_sc_hd__xor2_1
X_23773_ _03614_ _03638_ VGND VGND VPWR VPWR _03639_ sky130_fd_sc_hd__xnor2_1
Xmax_length7637 net7638 VGND VGND VPWR VPWR net7637 sky130_fd_sc_hd__buf_1
X_20985_ _00979_ _00999_ _01000_ VGND VGND VPWR VPWR _01001_ sky130_fd_sc_hd__o21a_2
XFILLER_0_79_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25512_ clknet_leaf_43_clk _00392_ net8778 VGND VGND VPWR VPWR svm0.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_22724_ _04865_ net4366 net4327 net3102 VGND VGND VPWR VPWR _02660_ sky130_fd_sc_hd__or4_1
Xmax_length6947 net6948 VGND VGND VPWR VPWR net6947 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25443_ clknet_leaf_113_clk _00326_ net8340 VGND VGND VPWR VPWR cordic0.vec\[1\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xmax_length6969 net6961 VGND VGND VPWR VPWR net6969 sky130_fd_sc_hd__clkbuf_1
X_22655_ _02180_ net3078 net941 _02612_ net8889 VGND VGND VPWR VPWR _00577_ sky130_fd_sc_hd__o311a_1
XFILLER_0_168_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21606_ net948 _01515_ net947 VGND VGND VPWR VPWR _01618_ sky130_fd_sc_hd__o21ba_1
X_25374_ clknet_leaf_57_clk _00257_ net8710 VGND VGND VPWR VPWR matmul0.alpha_pass\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22586_ net7317 _02554_ net7306 VGND VGND VPWR VPWR _02565_ sky130_fd_sc_hd__o21ai_1
Xfanout6118 net6124 VGND VGND VPWR VPWR net6118 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24325_ net7524 _04176_ net510 net7464 net460 VGND VGND VPWR VPWR _04185_ sky130_fd_sc_hd__a221o_1
Xfanout5406 net5421 VGND VGND VPWR VPWR net5406 sky130_fd_sc_hd__clkbuf_2
Xwire6202 net6203 VGND VGND VPWR VPWR net6202 sky130_fd_sc_hd__buf_1
X_21537_ net705 net703 _01328_ _01548_ net759 VGND VGND VPWR VPWR _01549_ sky130_fd_sc_hd__a2111o_1
Xwire6213 net6212 VGND VGND VPWR VPWR net6213 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6224 net6227 VGND VGND VPWR VPWR net6224 sky130_fd_sc_hd__buf_1
XFILLER_0_161_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6235 net6236 VGND VGND VPWR VPWR net6235 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24256_ pid_q.curr_int\[9\] net3758 _02870_ _04116_ VGND VGND VPWR VPWR _00674_ sky130_fd_sc_hd__a22o_1
Xwire5501 net5502 VGND VGND VPWR VPWR net5501 sky130_fd_sc_hd__buf_1
Xwire6246 net6243 VGND VGND VPWR VPWR net6246 sky130_fd_sc_hd__buf_1
Xwire6257 net6253 VGND VGND VPWR VPWR net6257 sky130_fd_sc_hd__buf_1
X_21468_ net1729 _01370_ _01359_ VGND VGND VPWR VPWR _01481_ sky130_fd_sc_hd__o21a_1
Xwire5534 net5539 VGND VGND VPWR VPWR net5534 sky130_fd_sc_hd__clkbuf_1
Xwire6279 net6280 VGND VGND VPWR VPWR net6279 sky130_fd_sc_hd__clkbuf_1
X_23207_ _03049_ _03050_ VGND VGND VPWR VPWR _03077_ sky130_fd_sc_hd__xor2_1
Xwire4800 net4805 VGND VGND VPWR VPWR net4800 sky130_fd_sc_hd__clkbuf_1
Xwire5545 net5546 VGND VGND VPWR VPWR net5545 sky130_fd_sc_hd__buf_1
Xwire4811 net4812 VGND VGND VPWR VPWR net4811 sky130_fd_sc_hd__buf_1
X_20419_ _12090_ net1500 VGND VGND VPWR VPWR _12215_ sky130_fd_sc_hd__or2_1
X_24187_ net739 _04046_ _04047_ VGND VGND VPWR VPWR _04048_ sky130_fd_sc_hd__o21ai_1
Xwire4822 net4821 VGND VGND VPWR VPWR net4822 sky130_fd_sc_hd__clkbuf_1
Xwire5567 net5563 VGND VGND VPWR VPWR net5567 sky130_fd_sc_hd__dlymetal6s2s_1
X_21399_ _01304_ _01309_ _01306_ net3789 VGND VGND VPWR VPWR _01413_ sky130_fd_sc_hd__a211o_1
Xwire4833 net4834 VGND VGND VPWR VPWR net4833 sky130_fd_sc_hd__clkbuf_1
Xwire5578 net5579 VGND VGND VPWR VPWR net5578 sky130_fd_sc_hd__buf_1
Xwire4844 net4848 VGND VGND VPWR VPWR net4844 sky130_fd_sc_hd__buf_1
Xwire5589 net5586 VGND VGND VPWR VPWR net5589 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23138_ _02984_ net1031 _02988_ _03006_ _03007_ VGND VGND VPWR VPWR _03008_ sky130_fd_sc_hd__a221o_1
Xwire4855 net4856 VGND VGND VPWR VPWR net4855 sky130_fd_sc_hd__buf_1
Xwire4866 net4867 VGND VGND VPWR VPWR net4866 sky130_fd_sc_hd__buf_1
Xmax_length1298 _06574_ VGND VGND VPWR VPWR net1298 sky130_fd_sc_hd__buf_1
Xwire4877 net4874 VGND VGND VPWR VPWR net4877 sky130_fd_sc_hd__clkbuf_1
Xwire4888 net4889 VGND VGND VPWR VPWR net4888 sky130_fd_sc_hd__buf_1
Xwire4899 net4900 VGND VGND VPWR VPWR net4899 sky130_fd_sc_hd__buf_1
X_23069_ _02876_ _02878_ _02938_ VGND VGND VPWR VPWR _02939_ sky130_fd_sc_hd__a21bo_1
X_15960_ net2646 net2637 VGND VGND VPWR VPWR _08028_ sky130_fd_sc_hd__nor2_2
XFILLER_0_41_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14911_ net4212 VGND VGND VPWR VPWR _06985_ sky130_fd_sc_hd__clkbuf_1
X_15891_ _07958_ _07959_ VGND VGND VPWR VPWR _07960_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17630_ svm0.tB\[11\] _09483_ VGND VGND VPWR VPWR _09511_ sky130_fd_sc_hd__or2_1
X_14842_ matmul0.a\[10\] matmul0.matmul_stage_inst.e\[10\] net3612 VGND VGND VPWR
+ VPWR _06938_ sky130_fd_sc_hd__mux2_1
X_17561_ _09393_ svm0.tC\[11\] _09442_ net6706 VGND VGND VPWR VPWR _09443_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_81_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14773_ net9003 net2857 net2866 _06899_ VGND VGND VPWR VPWR _00162_ sky130_fd_sc_hd__a22o_1
X_19300_ net6258 _10814_ VGND VGND VPWR VPWR _11137_ sky130_fd_sc_hd__xnor2_1
X_16512_ _08510_ _08519_ _08571_ VGND VGND VPWR VPWR _08572_ sky130_fd_sc_hd__a21o_1
XFILLER_0_184_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13724_ _05921_ _05924_ VGND VGND VPWR VPWR _05993_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17492_ net4027 net2567 _09379_ _09381_ VGND VGND VPWR VPWR _00399_ sky130_fd_sc_hd__a31o_1
XFILLER_0_168_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19231_ _11043_ _11039_ VGND VGND VPWR VPWR _11068_ sky130_fd_sc_hd__xnor2_1
X_16443_ net1084 _08502_ _08503_ VGND VGND VPWR VPWR _08504_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_195_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13655_ net7866 net1928 VGND VGND VPWR VPWR _05925_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8054 net8064 VGND VGND VPWR VPWR net8054 sky130_fd_sc_hd__buf_1
XFILLER_0_2_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12606_ net3699 VGND VGND VPWR VPWR _00008_ sky130_fd_sc_hd__buf_1
X_19162_ _10997_ _10998_ VGND VGND VPWR VPWR _10999_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13586_ net2371 VGND VGND VPWR VPWR _05857_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16374_ net1087 net1079 _08408_ VGND VGND VPWR VPWR _08436_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_183_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8160 net8161 VGND VGND VPWR VPWR net8160 sky130_fd_sc_hd__clkbuf_1
X_18113_ _09962_ _09963_ _09875_ VGND VGND VPWR VPWR _09964_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_182_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8171 net8172 VGND VGND VPWR VPWR net8171 sky130_fd_sc_hd__clkbuf_1
X_15325_ net2256 net2252 net1902 VGND VGND VPWR VPWR _07399_ sky130_fd_sc_hd__o21a_1
XFILLER_0_136_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8182 net8183 VGND VGND VPWR VPWR net8182 sky130_fd_sc_hd__clkbuf_1
X_19093_ net6292 net6244 VGND VGND VPWR VPWR _10930_ sky130_fd_sc_hd__nand2_1
Xfanout6641 net6645 VGND VGND VPWR VPWR net6641 sky130_fd_sc_hd__clkbuf_1
Xwire8193 net35 VGND VGND VPWR VPWR net8193 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6663 svm0.state\[2\] VGND VGND VPWR VPWR net6663 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18044_ net2551 _09894_ VGND VGND VPWR VPWR _09895_ sky130_fd_sc_hd__xnor2_2
Xwire7481 net7482 VGND VGND VPWR VPWR net7481 sky130_fd_sc_hd__buf_1
X_15256_ net990 _07326_ _07329_ VGND VGND VPWR VPWR _07330_ sky130_fd_sc_hd__o21ai_1
Xwire7492 net7493 VGND VGND VPWR VPWR net7492 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14207_ _06450_ _06452_ _06465_ _06403_ VGND VGND VPWR VPWR _06466_ sky130_fd_sc_hd__a2bb2o_1
X_15187_ _07255_ _07257_ _07260_ VGND VGND VPWR VPWR _07261_ sky130_fd_sc_hd__a21o_1
Xwire6791 net6788 VGND VGND VPWR VPWR net6791 sky130_fd_sc_hd__buf_1
X_14138_ net9198 net1308 net174 net2375 VGND VGND VPWR VPWR _00027_ sky130_fd_sc_hd__a22o_1
X_19995_ _11667_ _11739_ _11741_ VGND VGND VPWR VPWR _11826_ sky130_fd_sc_hd__o21a_1
XFILLER_0_190_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14069_ _06325_ _06331_ VGND VGND VPWR VPWR _06332_ sky130_fd_sc_hd__xnor2_2
X_18946_ net6375 net207 _10772_ VGND VGND VPWR VPWR _10784_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_3_clk clknet_4_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18877_ _10716_ _10717_ VGND VGND VPWR VPWR _10719_ sky130_fd_sc_hd__and2_1
X_17828_ net7122 net7139 VGND VGND VPWR VPWR _09679_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17759_ net6996 net3997 _09607_ _09608_ _09609_ VGND VGND VPWR VPWR _09610_ sky130_fd_sc_hd__a221o_1
XFILLER_0_178_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20770_ _12537_ _12538_ _12540_ VGND VGND VPWR VPWR _12541_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_18_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19429_ _11265_ VGND VGND VPWR VPWR _11266_ sky130_fd_sc_hd__inv_2
XFILLER_0_174_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22440_ net1169 _02344_ _02441_ VGND VGND VPWR VPWR _02442_ sky130_fd_sc_hd__o21a_1
XFILLER_0_162_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22371_ net5817 _02372_ _02373_ net2051 VGND VGND VPWR VPWR _02374_ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24110_ _03879_ _03881_ _03880_ VGND VGND VPWR VPWR _03972_ sky130_fd_sc_hd__o21a_1
XFILLER_0_26_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_107_Left_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21322_ net9009 net3122 net2077 _01336_ VGND VGND VPWR VPWR _00520_ sky130_fd_sc_hd__a22o_1
X_25090_ net4401 _04787_ _04832_ VGND VGND VPWR VPWR _04835_ sky130_fd_sc_hd__or3_1
XFILLER_0_130_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24041_ net4652 net4801 _03902_ VGND VGND VPWR VPWR _03904_ sky130_fd_sc_hd__a21oi_1
Xwire4107 _07131_ VGND VGND VPWR VPWR net4107 sky130_fd_sc_hd__clkbuf_1
X_21253_ _01264_ _01267_ VGND VGND VPWR VPWR _01268_ sky130_fd_sc_hd__xnor2_2
Xwire4118 _07089_ VGND VGND VPWR VPWR net4118 sky130_fd_sc_hd__buf_1
Xwire4129 net4130 VGND VGND VPWR VPWR net4129 sky130_fd_sc_hd__buf_1
XFILLER_0_187_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3406 _07574_ VGND VGND VPWR VPWR net3406 sky130_fd_sc_hd__buf_1
X_20204_ net243 _12028_ net3126 VGND VGND VPWR VPWR _12029_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_130_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21184_ net5638 net5878 _01172_ _01180_ VGND VGND VPWR VPWR _01200_ sky130_fd_sc_hd__a211o_1
Xwire3417 net3418 VGND VGND VPWR VPWR net3417 sky130_fd_sc_hd__buf_1
XFILLER_0_187_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3428 net3430 VGND VGND VPWR VPWR net3428 sky130_fd_sc_hd__buf_1
XFILLER_0_96_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2705 net2706 VGND VGND VPWR VPWR net2705 sky130_fd_sc_hd__buf_1
XFILLER_0_25_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2716 net2718 VGND VGND VPWR VPWR net2716 sky130_fd_sc_hd__clkbuf_1
X_20135_ _11914_ _11962_ VGND VGND VPWR VPWR _11963_ sky130_fd_sc_hd__or2_1
Xwire2727 net2728 VGND VGND VPWR VPWR net2727 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2738 net2739 VGND VGND VPWR VPWR net2738 sky130_fd_sc_hd__clkbuf_1
Xwire2749 _07205_ VGND VGND VPWR VPWR net2749 sky130_fd_sc_hd__clkbuf_1
X_24943_ pid_q.ki\[10\] _04722_ net1636 VGND VGND VPWR VPWR _04723_ sky130_fd_sc_hd__mux2_1
X_20066_ _11892_ net2493 VGND VGND VPWR VPWR _11895_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_116_Left_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24874_ pid_q.ki\[6\] net2397 net3009 pid_q.kp\[6\] VGND VGND VPWR VPWR _04674_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23825_ _03589_ _03591_ VGND VGND VPWR VPWR _03690_ sky130_fd_sc_hd__nor2_1
Xmax_length6700 net6697 VGND VGND VPWR VPWR net6700 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length7445 net7446 VGND VGND VPWR VPWR net7445 sky130_fd_sc_hd__clkbuf_1
Xmax_length6711 net6712 VGND VGND VPWR VPWR net6711 sky130_fd_sc_hd__clkbuf_1
X_23756_ _03489_ _03491_ _03621_ VGND VGND VPWR VPWR _03622_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_166_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20968_ net5621 net5821 VGND VGND VPWR VPWR _00984_ sky130_fd_sc_hd__nand2_1
Xmax_length7478 pid_q.state\[4\] VGND VGND VPWR VPWR net7478 sky130_fd_sc_hd__clkbuf_1
Xmax_length6744 svm0.delta\[1\] VGND VGND VPWR VPWR net6744 sky130_fd_sc_hd__buf_1
Xmax_length7489 net7483 VGND VGND VPWR VPWR net7489 sky130_fd_sc_hd__buf_1
XFILLER_0_166_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22707_ _02646_ VGND VGND VPWR VPWR _00595_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23687_ _03552_ _03553_ VGND VGND VPWR VPWR _03554_ sky130_fd_sc_hd__and2b_1
XFILLER_0_138_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20899_ _00906_ _00910_ _00891_ VGND VGND VPWR VPWR _00915_ sky130_fd_sc_hd__and3_1
X_13440_ net1129 net1128 VGND VGND VPWR VPWR _05713_ sky130_fd_sc_hd__xor2_1
X_22638_ net3821 _02600_ net2455 net2070 net3717 VGND VGND VPWR VPWR _00569_ sky130_fd_sc_hd__a221oi_1
X_25426_ clknet_leaf_91_clk _00309_ net8427 VGND VGND VPWR VPWR matmul0.cos\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13371_ net1130 _05643_ VGND VGND VPWR VPWR _05644_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_125_Left_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25357_ clknet_leaf_84_clk _00240_ net8723 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult2\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_22569_ net7369 net7352 net7343 VGND VGND VPWR VPWR _02551_ sky130_fd_sc_hd__or3_1
XFILLER_0_1_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire6010 net6007 VGND VGND VPWR VPWR net6010 sky130_fd_sc_hd__buf_1
XFILLER_0_133_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6021 net6022 VGND VGND VPWR VPWR net6021 sky130_fd_sc_hd__clkbuf_2
X_15110_ _07120_ _07115_ VGND VGND VPWR VPWR _07184_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24308_ net634 net633 VGND VGND VPWR VPWR _04168_ sky130_fd_sc_hd__xnor2_2
X_16090_ _08150_ _08156_ VGND VGND VPWR VPWR _08157_ sky130_fd_sc_hd__xnor2_1
Xwire6032 net6033 VGND VGND VPWR VPWR net6032 sky130_fd_sc_hd__buf_1
Xwire6043 net6041 VGND VGND VPWR VPWR net6043 sky130_fd_sc_hd__buf_1
XFILLER_0_50_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25288_ clknet_leaf_89_clk _00171_ net8422 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.a\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire5320 net5321 VGND VGND VPWR VPWR net5320 sky130_fd_sc_hd__clkbuf_1
Xwire6065 net6066 VGND VGND VPWR VPWR net6065 sky130_fd_sc_hd__buf_1
X_15041_ _07112_ _07114_ VGND VGND VPWR VPWR _07115_ sky130_fd_sc_hd__xnor2_1
X_24239_ _04012_ _04098_ _04099_ VGND VGND VPWR VPWR _04100_ sky130_fd_sc_hd__o21a_1
Xwire5331 net5332 VGND VGND VPWR VPWR net5331 sky130_fd_sc_hd__clkbuf_1
Xwire6076 cordic0.vec\[0\]\[14\] VGND VGND VPWR VPWR net6076 sky130_fd_sc_hd__buf_1
XFILLER_0_160_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5342 net5343 VGND VGND VPWR VPWR net5342 sky130_fd_sc_hd__clkbuf_1
Xwire6087 net6084 VGND VGND VPWR VPWR net6087 sky130_fd_sc_hd__buf_1
Xwire5353 pid_d.out\[9\] VGND VGND VPWR VPWR net5353 sky130_fd_sc_hd__clkbuf_1
Xwire6098 net6099 VGND VGND VPWR VPWR net6098 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_142_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5364 pid_d.out\[5\] VGND VGND VPWR VPWR net5364 sky130_fd_sc_hd__buf_1
Xwire5375 net5377 VGND VGND VPWR VPWR net5375 sky130_fd_sc_hd__buf_1
Xwire4641 net4642 VGND VGND VPWR VPWR net4641 sky130_fd_sc_hd__buf_1
Xwire5386 net5381 VGND VGND VPWR VPWR net5386 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4652 net4653 VGND VGND VPWR VPWR net4652 sky130_fd_sc_hd__buf_1
Xwire5397 net5391 VGND VGND VPWR VPWR net5397 sky130_fd_sc_hd__buf_1
XFILLER_0_102_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4663 net4665 VGND VGND VPWR VPWR net4663 sky130_fd_sc_hd__clkbuf_1
Xwire4674 net4675 VGND VGND VPWR VPWR net4674 sky130_fd_sc_hd__buf_1
X_18800_ _10640_ _10643_ VGND VGND VPWR VPWR _10644_ sky130_fd_sc_hd__nor2_1
Xwire4685 net4687 VGND VGND VPWR VPWR net4685 sky130_fd_sc_hd__buf_1
Xwire3940 _09934_ VGND VGND VPWR VPWR net3940 sky130_fd_sc_hd__clkbuf_1
X_19780_ _11542_ net604 VGND VGND VPWR VPWR _11614_ sky130_fd_sc_hd__or2_1
Xwire4696 net4697 VGND VGND VPWR VPWR net4696 sky130_fd_sc_hd__clkbuf_1
X_16992_ net5995 VGND VGND VPWR VPWR _08954_ sky130_fd_sc_hd__inv_2
Xwire3962 _09795_ VGND VGND VPWR VPWR net3962 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_196_Right_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire3973 _09685_ VGND VGND VPWR VPWR net3973 sky130_fd_sc_hd__clkbuf_1
Xwire3984 _09663_ VGND VGND VPWR VPWR net3984 sky130_fd_sc_hd__clkbuf_1
X_18731_ _10533_ _10534_ _10573_ net6896 VGND VGND VPWR VPWR _10576_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_134_Left_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire3995 _09624_ VGND VGND VPWR VPWR net3995 sky130_fd_sc_hd__buf_1
X_15943_ _08011_ VGND VGND VPWR VPWR _00220_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18662_ net6379 _10506_ _10508_ VGND VGND VPWR VPWR _10509_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15874_ net2714 net2812 net3422 _07694_ VGND VGND VPWR VPWR _07943_ sky130_fd_sc_hd__and4_1
X_17613_ net4023 svm0.tB\[5\] svm0.tB\[4\] net4009 VGND VGND VPWR VPWR _09494_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14825_ _06929_ VGND VGND VPWR VPWR _00184_ sky130_fd_sc_hd__clkbuf_1
X_18593_ net1762 _10440_ VGND VGND VPWR VPWR _10441_ sky130_fd_sc_hd__xnor2_2
X_17544_ net6692 VGND VGND VPWR VPWR _09426_ sky130_fd_sc_hd__inv_2
X_14756_ _06842_ _06886_ VGND VGND VPWR VPWR _06887_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13707_ _05974_ _05975_ VGND VGND VPWR VPWR _05976_ sky130_fd_sc_hd__xor2_1
X_17475_ net6729 _09366_ _09362_ VGND VGND VPWR VPWR _09367_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_6_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14687_ matmul0.sin\[4\] _06832_ VGND VGND VPWR VPWR _06835_ sky130_fd_sc_hd__nor2_1
X_19214_ net6287 net6337 VGND VGND VPWR VPWR _11051_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_143_Left_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16426_ _08428_ _08481_ _08482_ _08427_ _08487_ VGND VGND VPWR VPWR _08488_ sky130_fd_sc_hd__o221a_1
XFILLER_0_172_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13638_ net7616 net1337 VGND VGND VPWR VPWR _05908_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_183_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19145_ _10974_ _10981_ VGND VGND VPWR VPWR _10982_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_54_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16357_ _08418_ net1247 VGND VGND VPWR VPWR _08420_ sky130_fd_sc_hd__xor2_1
X_13569_ net7895 net1928 _05839_ VGND VGND VPWR VPWR _05840_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6460 net6465 VGND VGND VPWR VPWR net6460 sky130_fd_sc_hd__clkbuf_2
X_15308_ net4192 net4186 net4176 net4174 VGND VGND VPWR VPWR _07382_ sky130_fd_sc_hd__o22a_1
X_19076_ net3211 _10912_ VGND VGND VPWR VPWR _10913_ sky130_fd_sc_hd__nor2_1
X_16288_ _08318_ _08351_ VGND VGND VPWR VPWR _08352_ sky130_fd_sc_hd__xor2_1
XFILLER_0_87_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18027_ net3949 _09877_ VGND VGND VPWR VPWR _09878_ sky130_fd_sc_hd__xnor2_2
X_15239_ _07310_ _07312_ VGND VGND VPWR VPWR _07313_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5792 net5797 VGND VGND VPWR VPWR net5792 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_50_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19978_ net2093 _11808_ VGND VGND VPWR VPWR _11809_ sky130_fd_sc_hd__xor2_1
XFILLER_0_157_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_163_Right_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18929_ net1437 _10768_ VGND VGND VPWR VPWR _10769_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21940_ _01837_ _01839_ _01947_ VGND VGND VPWR VPWR _01948_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_55_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21871_ net2066 _01792_ VGND VGND VPWR VPWR _01880_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23610_ _03475_ _03476_ _03477_ VGND VGND VPWR VPWR _03478_ sky130_fd_sc_hd__and3_1
X_20822_ net1737 _00837_ VGND VGND VPWR VPWR _00838_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_173_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24590_ pid_q.prev_error\[14\] pid_q.curr_error\[14\] VGND VGND VPWR VPWR _04446_
+ sky130_fd_sc_hd__and2_1
Xmax_length6029 net6030 VGND VGND VPWR VPWR net6029 sky130_fd_sc_hd__buf_1
X_23541_ _03328_ net2426 _03326_ VGND VGND VPWR VPWR _03409_ sky130_fd_sc_hd__o21a_1
XFILLER_0_187_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20753_ _12521_ _12522_ VGND VGND VPWR VPWR _12524_ sky130_fd_sc_hd__nor2_1
Xwire8907 net8908 VGND VGND VPWR VPWR net8907 sky130_fd_sc_hd__buf_1
Xmax_length5339 pid_d.out\[12\] VGND VGND VPWR VPWR net5339 sky130_fd_sc_hd__buf_1
Xwire8918 net8919 VGND VGND VPWR VPWR net8918 sky130_fd_sc_hd__clkbuf_1
Xwire8929 net8930 VGND VGND VPWR VPWR net8929 sky130_fd_sc_hd__clkbuf_1
X_23472_ _03337_ _03340_ VGND VGND VPWR VPWR _03341_ sky130_fd_sc_hd__xnor2_2
X_20684_ _12458_ _12459_ VGND VGND VPWR VPWR _12460_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25211_ clknet_leaf_64_clk _00100_ net8661 VGND VGND VPWR VPWR matmul0.op_in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire608 net609 VGND VGND VPWR VPWR net608 sky130_fd_sc_hd__clkbuf_1
X_22423_ net5708 _02349_ VGND VGND VPWR VPWR _02425_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire619 net620 VGND VGND VPWR VPWR net619 sky130_fd_sc_hd__buf_1
XFILLER_0_163_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25142_ clknet_leaf_50_clk _00031_ net8757 VGND VGND VPWR VPWR svm0.tC\[14\] sky130_fd_sc_hd__dfrtp_1
X_22354_ _02351_ _02356_ VGND VGND VPWR VPWR _02357_ sky130_fd_sc_hd__xor2_1
XFILLER_0_115_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21305_ net3796 net3119 _00864_ VGND VGND VPWR VPWR _01320_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_131_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25073_ _04817_ _04818_ VGND VGND VPWR VPWR _04820_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22285_ _02210_ _02211_ _02212_ VGND VGND VPWR VPWR _02289_ sky130_fd_sc_hd__o21a_1
XFILLER_0_142_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24024_ net4486 _03886_ VGND VGND VPWR VPWR _03887_ sky130_fd_sc_hd__nand2_2
Xhold250 _00424_ VGND VGND VPWR VPWR net9203 sky130_fd_sc_hd__dlygate4sd3_1
X_21236_ net761 net760 _01220_ _01239_ VGND VGND VPWR VPWR _01251_ sky130_fd_sc_hd__a211o_1
Xhold261 svm0.tB\[15\] VGND VGND VPWR VPWR net9214 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3214 _10805_ VGND VGND VPWR VPWR net3214 sky130_fd_sc_hd__clkbuf_2
Xhold272 matmul0.b\[11\] VGND VGND VPWR VPWR net9225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 pid_d.prev_int\[5\] VGND VGND VPWR VPWR net9236 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3236 _09880_ VGND VGND VPWR VPWR net3236 sky130_fd_sc_hd__clkbuf_1
X_21167_ _01168_ _01169_ net3816 VGND VGND VPWR VPWR _01183_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2502 net2503 VGND VGND VPWR VPWR net2502 sky130_fd_sc_hd__clkbuf_2
Xwire3247 _09675_ VGND VGND VPWR VPWR net3247 sky130_fd_sc_hd__buf_1
Xwire2513 net2515 VGND VGND VPWR VPWR net2513 sky130_fd_sc_hd__buf_1
Xwire3258 _09643_ VGND VGND VPWR VPWR net3258 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3269 _09575_ VGND VGND VPWR VPWR net3269 sky130_fd_sc_hd__buf_1
Xwire2524 net2525 VGND VGND VPWR VPWR net2524 sky130_fd_sc_hd__clkbuf_1
Xwire2535 net2536 VGND VGND VPWR VPWR net2535 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1801 _09099_ VGND VGND VPWR VPWR net1801 sky130_fd_sc_hd__clkbuf_2
X_20118_ _11944_ _11945_ VGND VGND VPWR VPWR _11946_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_130_Right_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2546 _10067_ VGND VGND VPWR VPWR net2546 sky130_fd_sc_hd__buf_1
Xwire1812 net1813 VGND VGND VPWR VPWR net1812 sky130_fd_sc_hd__clkbuf_1
Xwire2557 net2558 VGND VGND VPWR VPWR net2557 sky130_fd_sc_hd__clkbuf_2
X_21098_ _01031_ _01113_ VGND VGND VPWR VPWR _01114_ sky130_fd_sc_hd__xnor2_1
Xwire2568 net2569 VGND VGND VPWR VPWR net2568 sky130_fd_sc_hd__buf_1
Xwire1823 net1824 VGND VGND VPWR VPWR net1823 sky130_fd_sc_hd__clkbuf_1
Xwire2579 _09272_ VGND VGND VPWR VPWR net2579 sky130_fd_sc_hd__buf_1
Xwire1834 net1835 VGND VGND VPWR VPWR net1834 sky130_fd_sc_hd__clkbuf_1
Xwire1845 _07942_ VGND VGND VPWR VPWR net1845 sky130_fd_sc_hd__buf_1
X_24926_ _04711_ VGND VGND VPWR VPWR _00749_ sky130_fd_sc_hd__clkbuf_1
X_12940_ _05005_ _05006_ VGND VGND VPWR VPWR _05213_ sky130_fd_sc_hd__xor2_1
X_20049_ _11848_ _11870_ _11877_ VGND VGND VPWR VPWR _11878_ sky130_fd_sc_hd__a21o_1
Xwire1856 _07619_ VGND VGND VPWR VPWR net1856 sky130_fd_sc_hd__clkbuf_1
Xwire1867 _07396_ VGND VGND VPWR VPWR net1867 sky130_fd_sc_hd__clkbuf_1
Xwire1878 _07308_ VGND VGND VPWR VPWR net1878 sky130_fd_sc_hd__clkbuf_2
Xwire1889 net1890 VGND VGND VPWR VPWR net1889 sky130_fd_sc_hd__buf_1
XFILLER_0_73_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24857_ pid_q.ki\[1\] net3022 net3007 pid_q.kp\[1\] VGND VGND VPWR VPWR _04662_ sky130_fd_sc_hd__a22o_1
X_12871_ _05088_ _05143_ VGND VGND VPWR VPWR _05144_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14610_ net2882 _06780_ _06781_ _06782_ net2887 VGND VGND VPWR VPWR _06783_ sky130_fd_sc_hd__o221a_1
X_23808_ _03670_ _03580_ _03672_ VGND VGND VPWR VPWR _03673_ sky130_fd_sc_hd__a21o_1
XFILLER_0_157_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15590_ net1859 _07582_ _07661_ VGND VGND VPWR VPWR _07662_ sky130_fd_sc_hd__o21a_1
X_24788_ net7967 VGND VGND VPWR VPWR _04614_ sky130_fd_sc_hd__inv_2
X_14541_ net7278 net5247 _06717_ _06718_ net2885 VGND VGND VPWR VPWR _06720_ sky130_fd_sc_hd__a311o_1
X_23739_ net4504 VGND VGND VPWR VPWR _03605_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6574 net6575 VGND VGND VPWR VPWR net6574 sky130_fd_sc_hd__buf_1
XFILLER_0_166_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17260_ net2981 VGND VGND VPWR VPWR _09191_ sky130_fd_sc_hd__buf_1
X_14472_ net7365 net5311 VGND VGND VPWR VPWR _06659_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length5873 net5874 VGND VGND VPWR VPWR net5873 sky130_fd_sc_hd__buf_1
X_16211_ _08187_ _08188_ _08275_ VGND VGND VPWR VPWR _08276_ sky130_fd_sc_hd__o21a_1
XFILLER_0_180_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13423_ net843 net842 _05629_ VGND VGND VPWR VPWR _05696_ sky130_fd_sc_hd__o21ba_1
X_25409_ clknet_leaf_80_clk _00292_ net8489 VGND VGND VPWR VPWR matmul0.a\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17191_ _09141_ VGND VGND VPWR VPWR _00338_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5011 net5027 VGND VGND VPWR VPWR net5011 sky130_fd_sc_hd__buf_1
XFILLER_0_125_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13354_ _05511_ net1133 VGND VGND VPWR VPWR _05627_ sky130_fd_sc_hd__nand2_1
X_16142_ _08186_ _08206_ VGND VGND VPWR VPWR _08208_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13285_ _05554_ net1132 VGND VGND VPWR VPWR _05558_ sky130_fd_sc_hd__xnor2_2
X_16073_ _08034_ net1261 _08139_ VGND VGND VPWR VPWR _08140_ sky130_fd_sc_hd__o21a_1
Xwire5150 net5151 VGND VGND VPWR VPWR net5150 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5161 net5165 VGND VGND VPWR VPWR net5161 sky130_fd_sc_hd__buf_1
X_19901_ _11661_ _11715_ VGND VGND VPWR VPWR _11733_ sky130_fd_sc_hd__nand2_1
X_15024_ net4190 net4184 _07026_ _07028_ VGND VGND VPWR VPWR _07098_ sky130_fd_sc_hd__o22a_1
Xwire5172 net5173 VGND VGND VPWR VPWR net5172 sky130_fd_sc_hd__clkbuf_2
Xwire5183 net5184 VGND VGND VPWR VPWR net5183 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire5194 net5195 VGND VGND VPWR VPWR net5194 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4460 net4461 VGND VGND VPWR VPWR net4460 sky130_fd_sc_hd__clkbuf_1
X_19832_ net604 _11663_ _11665_ VGND VGND VPWR VPWR _11666_ sky130_fd_sc_hd__a21oi_1
Xwire4471 net4472 VGND VGND VPWR VPWR net4471 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4493 net4494 VGND VGND VPWR VPWR net4493 sky130_fd_sc_hd__buf_1
XFILLER_0_78_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3770 net3771 VGND VGND VPWR VPWR net3770 sky130_fd_sc_hd__buf_1
X_19763_ _11594_ _11596_ VGND VGND VPWR VPWR _11598_ sky130_fd_sc_hd__nand2_1
Xwire3781 net3782 VGND VGND VPWR VPWR net3781 sky130_fd_sc_hd__clkbuf_1
X_16975_ net5989 net1825 _08937_ _08924_ VGND VGND VPWR VPWR _08938_ sky130_fd_sc_hd__a211o_1
Xwire3792 net3793 VGND VGND VPWR VPWR net3792 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18714_ _10558_ _10559_ VGND VGND VPWR VPWR _10560_ sky130_fd_sc_hd__nor2_1
X_15926_ _07988_ _07994_ VGND VGND VPWR VPWR _07995_ sky130_fd_sc_hd__xnor2_1
X_19694_ net1058 _11528_ VGND VGND VPWR VPWR _11530_ sky130_fd_sc_hd__nand2_1
Xinput7 angle_in[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
X_18645_ _10485_ _10491_ VGND VGND VPWR VPWR _10492_ sky130_fd_sc_hd__xnor2_1
X_15857_ net827 _07888_ _07925_ VGND VGND VPWR VPWR _07926_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14808_ net7442 net7172 net3628 VGND VGND VPWR VPWR _06921_ sky130_fd_sc_hd__a21o_1
X_18576_ net3308 _10171_ VGND VGND VPWR VPWR _10424_ sky130_fd_sc_hd__or2_1
X_15788_ net1264 _07856_ VGND VGND VPWR VPWR _07858_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17527_ svm0.delta\[14\] _09410_ VGND VGND VPWR VPWR _09411_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14739_ _06832_ VGND VGND VPWR VPWR _06873_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17458_ svm0.counter\[3\] _09351_ _09352_ _09350_ VGND VGND VPWR VPWR _00394_ sky130_fd_sc_hd__a22o_1
XFILLER_0_184_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16409_ _08469_ _08468_ VGND VGND VPWR VPWR _08471_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17389_ net2572 _09296_ VGND VGND VPWR VPWR _09297_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19128_ _10960_ _10964_ VGND VGND VPWR VPWR _10965_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_131_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6290 net6305 VGND VGND VPWR VPWR net6290 sky130_fd_sc_hd__dlymetal6s2s_1
X_19059_ net3208 _10895_ VGND VGND VPWR VPWR _10896_ sky130_fd_sc_hd__xnor2_1
X_22070_ _01959_ net1713 _02075_ _02076_ VGND VGND VPWR VPWR _02077_ sky130_fd_sc_hd__o22a_1
XFILLER_0_168_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21021_ net5631 net5831 VGND VGND VPWR VPWR _01037_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1108 _07660_ VGND VGND VPWR VPWR net1108 sky130_fd_sc_hd__buf_1
XFILLER_0_96_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25760_ clknet_leaf_95_clk _00633_ net8455 VGND VGND VPWR VPWR pid_d.out\[1\] sky130_fd_sc_hd__dfrtp_1
X_22972_ net9238 net1240 net6570 VGND VGND VPWR VPWR _02854_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24711_ net5290 _04546_ VGND VGND VPWR VPWR _04547_ sky130_fd_sc_hd__xnor2_1
X_21923_ _01929_ _01930_ VGND VGND VPWR VPWR _01931_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_179_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25691_ clknet_leaf_3_clk _00564_ net8569 VGND VGND VPWR VPWR pid_d.curr_error\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24642_ _04467_ _04496_ VGND VGND VPWR VPWR _04497_ sky130_fd_sc_hd__xnor2_1
X_21854_ net5809 VGND VGND VPWR VPWR _01863_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20805_ net5960 net5414 VGND VGND VPWR VPWR _00821_ sky130_fd_sc_hd__nand2_1
X_24573_ net4919 net4894 net4871 _04351_ VGND VGND VPWR VPWR _04429_ sky130_fd_sc_hd__a31o_1
X_21785_ _01698_ _01704_ _01703_ VGND VGND VPWR VPWR _01795_ sky130_fd_sc_hd__a21o_1
XFILLER_0_93_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8704 net8705 VGND VGND VPWR VPWR net8704 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23524_ net5180 pid_q.prev_int\[2\] VGND VGND VPWR VPWR _03392_ sky130_fd_sc_hd__xnor2_1
Xwire8715 net8716 VGND VGND VPWR VPWR net8715 sky130_fd_sc_hd__dlymetal6s2s_1
X_20736_ _12505_ _12506_ VGND VGND VPWR VPWR _12507_ sky130_fd_sc_hd__xor2_1
Xwire8726 net8722 VGND VGND VPWR VPWR net8726 sky130_fd_sc_hd__buf_1
Xwire8737 net8738 VGND VGND VPWR VPWR net8737 sky130_fd_sc_hd__clkbuf_1
Xmax_length4424 pid_q.out\[10\] VGND VGND VPWR VPWR net4424 sky130_fd_sc_hd__buf_1
Xwire8748 net8750 VGND VGND VPWR VPWR net8748 sky130_fd_sc_hd__buf_1
Xmax_length4435 pid_q.out\[8\] VGND VGND VPWR VPWR net4435 sky130_fd_sc_hd__clkbuf_1
Xwire8759 net8756 VGND VGND VPWR VPWR net8759 sky130_fd_sc_hd__dlymetal6s2s_1
X_23455_ net4563 net5080 VGND VGND VPWR VPWR _03324_ sky130_fd_sc_hd__nand2_1
XFILLER_0_162_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4457 pid_q.out\[4\] VGND VGND VPWR VPWR net4457 sky130_fd_sc_hd__buf_1
Xwire405 net406 VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20667_ net1394 _12429_ net1077 VGND VGND VPWR VPWR _12444_ sky130_fd_sc_hd__o21a_1
Xwire416 net417 VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__buf_1
XFILLER_0_135_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire427 net428 VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__clkbuf_1
Xwire438 net439 VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__clkbuf_1
Xwire449 net450 VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__clkbuf_2
X_22406_ net4382 _02399_ _02400_ net206 VGND VGND VPWR VPWR _02408_ sky130_fd_sc_hd__a31o_1
Xmax_length3756 _02925_ VGND VGND VPWR VPWR net3756 sky130_fd_sc_hd__clkbuf_1
X_23386_ _03193_ _03190_ _03255_ VGND VGND VPWR VPWR _03256_ sky130_fd_sc_hd__o21a_1
XFILLER_0_162_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20598_ _12375_ _12379_ VGND VGND VPWR VPWR _12380_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22337_ _02304_ _02309_ _02311_ VGND VGND VPWR VPWR _02340_ sky130_fd_sc_hd__a21o_1
X_25125_ net9109 _04849_ net2391 pid_d.curr_int\[13\] VGND VGND VPWR VPWR _00806_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13070_ net6673 net6677 net7232 VGND VGND VPWR VPWR _05343_ sky130_fd_sc_hd__and3b_1
X_25056_ net3737 net685 pid_q.out\[8\] VGND VGND VPWR VPWR _04805_ sky130_fd_sc_hd__o21ba_1
X_22268_ _02269_ _02185_ _02271_ VGND VGND VPWR VPWR _02272_ sky130_fd_sc_hd__a21o_1
XFILLER_0_103_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24007_ net3749 _03821_ net5149 VGND VGND VPWR VPWR _03870_ sky130_fd_sc_hd__o21ai_1
Xwire3011 net3012 VGND VGND VPWR VPWR net3011 sky130_fd_sc_hd__clkbuf_1
Xwire3022 net3023 VGND VGND VPWR VPWR net3022 sky130_fd_sc_hd__buf_1
XFILLER_0_104_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21219_ net808 _01078_ _01027_ _01234_ VGND VGND VPWR VPWR _01235_ sky130_fd_sc_hd__o22a_1
Xwire3033 _04849_ VGND VGND VPWR VPWR net3033 sky130_fd_sc_hd__buf_1
Xwire3044 net3045 VGND VGND VPWR VPWR net3044 sky130_fd_sc_hd__buf_1
X_22199_ net1036 _02202_ _02203_ VGND VGND VPWR VPWR _02204_ sky130_fd_sc_hd__o21a_1
Xwire2310 _05129_ VGND VGND VPWR VPWR net2310 sky130_fd_sc_hd__buf_1
XFILLER_0_40_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2321 net2322 VGND VGND VPWR VPWR net2321 sky130_fd_sc_hd__buf_1
Xwire3066 net3067 VGND VGND VPWR VPWR net3066 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2332 net2333 VGND VGND VPWR VPWR net2332 sky130_fd_sc_hd__buf_1
Xwire3077 net3078 VGND VGND VPWR VPWR net3077 sky130_fd_sc_hd__clkbuf_2
Xwire2343 _04925_ VGND VGND VPWR VPWR net2343 sky130_fd_sc_hd__clkbuf_1
Xwire3088 _02561_ VGND VGND VPWR VPWR net3088 sky130_fd_sc_hd__buf_1
Xwire2354 net2355 VGND VGND VPWR VPWR net2354 sky130_fd_sc_hd__buf_1
Xwire3099 net3100 VGND VGND VPWR VPWR net3099 sky130_fd_sc_hd__clkbuf_1
Xwire2365 net2366 VGND VGND VPWR VPWR net2365 sky130_fd_sc_hd__buf_1
Xwire2376 net2377 VGND VGND VPWR VPWR net2376 sky130_fd_sc_hd__buf_1
Xwire1631 net1632 VGND VGND VPWR VPWR net1631 sky130_fd_sc_hd__buf_1
X_16760_ matmul0.a_in\[0\] matmul0.a\[0\] net3382 VGND VGND VPWR VPWR _08769_ sky130_fd_sc_hd__mux2_1
X_13972_ net1583 _06236_ net7601 VGND VGND VPWR VPWR _06237_ sky130_fd_sc_hd__mux2_1
Xwire1642 _04542_ VGND VGND VPWR VPWR net1642 sky130_fd_sc_hd__buf_1
Xwire2387 net2388 VGND VGND VPWR VPWR net2387 sky130_fd_sc_hd__clkbuf_1
Xwire2398 _04664_ VGND VGND VPWR VPWR net2398 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1653 _04149_ VGND VGND VPWR VPWR net1653 sky130_fd_sc_hd__buf_1
XFILLER_0_189_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1664 net1665 VGND VGND VPWR VPWR net1664 sky130_fd_sc_hd__clkbuf_1
Xwire1675 _03185_ VGND VGND VPWR VPWR net1675 sky130_fd_sc_hd__clkbuf_2
X_15711_ _07779_ _07781_ VGND VGND VPWR VPWR _07782_ sky130_fd_sc_hd__xor2_1
XFILLER_0_88_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24909_ _04695_ _04696_ _04697_ _04698_ VGND VGND VPWR VPWR _04699_ sky130_fd_sc_hd__or4_1
X_12923_ _05194_ _05195_ _05108_ _05109_ VGND VGND VPWR VPWR _05196_ sky130_fd_sc_hd__or4_1
XFILLER_0_77_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1686 net1687 VGND VGND VPWR VPWR net1686 sky130_fd_sc_hd__clkbuf_1
X_16691_ _08721_ VGND VGND VPWR VPWR _00258_ sky130_fd_sc_hd__clkbuf_1
X_25889_ clknet_leaf_17_clk _00762_ net8628 VGND VGND VPWR VPWR pid_q.kp\[1\] sky130_fd_sc_hd__dfrtp_1
Xwire1697 net1698 VGND VGND VPWR VPWR net1697 sky130_fd_sc_hd__clkbuf_1
X_18430_ _10278_ _10279_ VGND VGND VPWR VPWR _10280_ sky130_fd_sc_hd__nor2_1
X_15642_ _07572_ _07573_ VGND VGND VPWR VPWR _07714_ sky130_fd_sc_hd__or2_1
X_12854_ net6749 net6599 net5236 VGND VGND VPWR VPWR _05127_ sky130_fd_sc_hd__and3_1
XFILLER_0_84_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18361_ net6789 _10171_ VGND VGND VPWR VPWR _10212_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_186_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15573_ _07627_ _07643_ _07644_ VGND VGND VPWR VPWR _07645_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_69_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12785_ net7875 net1602 VGND VGND VPWR VPWR _05058_ sky130_fd_sc_hd__xnor2_1
X_17312_ _09221_ _09222_ _09224_ VGND VGND VPWR VPWR _09226_ sky130_fd_sc_hd__mux2_1
X_14524_ net7278 net5246 VGND VGND VPWR VPWR _06704_ sky130_fd_sc_hd__xnor2_1
X_18292_ net963 _09835_ _09829_ VGND VGND VPWR VPWR _10143_ sky130_fd_sc_hd__and3b_1
XFILLER_0_44_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17243_ net2161 VGND VGND VPWR VPWR _09190_ sky130_fd_sc_hd__buf_1
X_14455_ _06645_ VGND VGND VPWR VPWR _00098_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13406_ _05654_ _05570_ VGND VGND VPWR VPWR _05679_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17174_ net6891 net670 VGND VGND VPWR VPWR _09126_ sky130_fd_sc_hd__and2_1
X_14386_ _06592_ net7580 net899 VGND VGND VPWR VPWR _06593_ sky130_fd_sc_hd__mux2_1
Xwire950 _12135_ VGND VGND VPWR VPWR net950 sky130_fd_sc_hd__clkbuf_2
Xwire961 _10382_ VGND VGND VPWR VPWR net961 sky130_fd_sc_hd__buf_1
Xwire972 net973 VGND VGND VPWR VPWR net972 sky130_fd_sc_hd__buf_1
Xwire983 _08204_ VGND VGND VPWR VPWR net983 sky130_fd_sc_hd__buf_1
X_16125_ _08187_ _08190_ VGND VGND VPWR VPWR _08191_ sky130_fd_sc_hd__xnor2_1
X_13337_ net7815 net1942 net2291 VGND VGND VPWR VPWR _05610_ sky130_fd_sc_hd__and3_1
Xwire994 net995 VGND VGND VPWR VPWR net994 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16056_ net2753 net2627 VGND VGND VPWR VPWR _08123_ sky130_fd_sc_hd__nor2_1
X_13268_ _05539_ _05540_ VGND VGND VPWR VPWR _05541_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15007_ net2827 _07015_ net3555 net2834 VGND VGND VPWR VPWR _07081_ sky130_fd_sc_hd__a211o_1
X_13199_ net919 _05360_ VGND VGND VPWR VPWR _05472_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19815_ net6034 _11648_ net3128 VGND VGND VPWR VPWR _11649_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16958_ net2177 net1825 VGND VGND VPWR VPWR _08921_ sky130_fd_sc_hd__xnor2_1
X_19746_ net3175 _10972_ _11521_ net6175 VGND VGND VPWR VPWR _11581_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15909_ _07871_ _07876_ _07869_ VGND VGND VPWR VPWR _07978_ sky130_fd_sc_hd__a21o_1
XFILLER_0_189_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19677_ net6220 net6286 VGND VGND VPWR VPWR _11513_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16889_ cordic0.slte0.opA\[14\] net6393 VGND VGND VPWR VPWR _08853_ sky130_fd_sc_hd__or2b_1
X_18628_ net6976 net6874 VGND VGND VPWR VPWR _10475_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_154_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_188_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18559_ net607 _10406_ VGND VGND VPWR VPWR _10407_ sky130_fd_sc_hd__nand2_1
X_21570_ _01570_ _01581_ VGND VGND VPWR VPWR _01582_ sky130_fd_sc_hd__xor2_1
XFILLER_0_145_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20521_ net1470 _12306_ _08909_ VGND VGND VPWR VPWR _12308_ sky130_fd_sc_hd__a21oi_1
Xmax_length3008 _00008_ VGND VGND VPWR VPWR net3008 sky130_fd_sc_hd__buf_1
XFILLER_0_144_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23240_ _03093_ _03095_ _03109_ VGND VGND VPWR VPWR _03110_ sky130_fd_sc_hd__a21o_1
X_20452_ net6515 net1501 net2586 _12136_ VGND VGND VPWR VPWR _12245_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_7_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5919 net5920 VGND VGND VPWR VPWR net5919 sky130_fd_sc_hd__clkbuf_1
X_23171_ net5116 net4719 _03039_ net4698 net5139 VGND VGND VPWR VPWR _03041_ sky130_fd_sc_hd__a32o_1
XFILLER_0_162_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length1617 _04920_ VGND VGND VPWR VPWR net1617 sky130_fd_sc_hd__buf_1
X_20383_ net6458 net4055 _12177_ _12180_ _12181_ VGND VGND VPWR VPWR _12182_ sky130_fd_sc_hd__o32a_1
XFILLER_0_113_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22122_ _02025_ _02027_ _02127_ VGND VGND VPWR VPWR _02128_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_30_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput152 net8075 VGND VGND VPWR VPWR ready sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22053_ _02057_ _02059_ VGND VGND VPWR VPWR _02060_ sky130_fd_sc_hd__and2_1
X_21004_ _00912_ _01019_ VGND VGND VPWR VPWR _01020_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_195_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25812_ clknet_leaf_36_clk _00685_ net8748 VGND VGND VPWR VPWR pid_q.prev_error\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25743_ clknet_leaf_8_clk _00616_ net8553 VGND VGND VPWR VPWR pid_d.kp\[1\] sky130_fd_sc_hd__dfrtp_1
X_22955_ net5314 net5974 VGND VGND VPWR VPWR _02843_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21906_ net4385 net803 net413 net4319 net699 VGND VGND VPWR VPWR _01915_ sky130_fd_sc_hd__a221o_1
X_25674_ clknet_leaf_4_clk _00547_ net8563 VGND VGND VPWR VPWR pid_d.prev_error\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22886_ net5357 _02777_ _02780_ VGND VGND VPWR VPWR _02781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24625_ _04296_ net4842 net4823 _04478_ VGND VGND VPWR VPWR _04480_ sky130_fd_sc_hd__a211o_1
X_21837_ net5764 net5461 VGND VGND VPWR VPWR _01846_ sky130_fd_sc_hd__and2_1
XFILLER_0_195_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout7705 net7712 VGND VGND VPWR VPWR net7705 sky130_fd_sc_hd__buf_1
X_12570_ net1987 VGND VGND VPWR VPWR _04860_ sky130_fd_sc_hd__buf_1
X_24556_ _04355_ _04364_ _04411_ VGND VGND VPWR VPWR _04412_ sky130_fd_sc_hd__a21oi_1
X_21768_ net5384 _01592_ VGND VGND VPWR VPWR _01778_ sky130_fd_sc_hd__and2_1
Xwire8512 net8517 VGND VGND VPWR VPWR net8512 sky130_fd_sc_hd__clkbuf_1
Xwire8523 net8524 VGND VGND VPWR VPWR net8523 sky130_fd_sc_hd__buf_1
XFILLER_0_110_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8534 net8535 VGND VGND VPWR VPWR net8534 sky130_fd_sc_hd__clkbuf_1
X_23507_ _03370_ net1024 VGND VGND VPWR VPWR _03376_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20719_ _12488_ _12490_ VGND VGND VPWR VPWR _12491_ sky130_fd_sc_hd__xnor2_1
Xwire8545 net8537 VGND VGND VPWR VPWR net8545 sky130_fd_sc_hd__clkbuf_1
Xwire7811 net7805 VGND VGND VPWR VPWR net7811 sky130_fd_sc_hd__buf_1
Xwire202 net203 VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_1
Xwire8556 net8557 VGND VGND VPWR VPWR net8556 sky130_fd_sc_hd__clkbuf_1
X_24487_ net4545 net4809 VGND VGND VPWR VPWR _04344_ sky130_fd_sc_hd__nand2_1
Xwire7822 net7823 VGND VGND VPWR VPWR net7822 sky130_fd_sc_hd__buf_1
X_21699_ net5891 net3107 net5384 VGND VGND VPWR VPWR _01710_ sky130_fd_sc_hd__o21ai_1
Xwire213 net214 VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_1
Xwire7833 net7834 VGND VGND VPWR VPWR net7833 sky130_fd_sc_hd__buf_1
Xwire8578 net8580 VGND VGND VPWR VPWR net8578 sky130_fd_sc_hd__buf_1
XFILLER_0_80_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire224 net225 VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__buf_1
Xmax_length4276 _04898_ VGND VGND VPWR VPWR net4276 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3531 net3532 VGND VGND VPWR VPWR net3531 sky130_fd_sc_hd__buf_1
XFILLER_0_68_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8589 net8585 VGND VGND VPWR VPWR net8589 sky130_fd_sc_hd__buf_1
Xwire235 net236 VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__clkbuf_1
X_14240_ net6456 net6649 net6446 VGND VGND VPWR VPWR _06496_ sky130_fd_sc_hd__o21a_1
X_23438_ net646 net640 _03307_ VGND VGND VPWR VPWR _03308_ sky130_fd_sc_hd__a21oi_1
Xwire7855 net7851 VGND VGND VPWR VPWR net7855 sky130_fd_sc_hd__buf_1
Xwire246 _10511_ VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__clkbuf_1
Xwire257 _06086_ VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__buf_1
Xwire7866 net7867 VGND VGND VPWR VPWR net7866 sky130_fd_sc_hd__buf_1
Xwire7877 net7873 VGND VGND VPWR VPWR net7877 sky130_fd_sc_hd__buf_1
Xmax_length3564 _07035_ VGND VGND VPWR VPWR net3564 sky130_fd_sc_hd__clkbuf_1
Xmax_length3575 net3576 VGND VGND VPWR VPWR net3575 sky130_fd_sc_hd__clkbuf_1
X_14171_ net9222 net1308 net157 net2375 VGND VGND VPWR VPWR _00028_ sky130_fd_sc_hd__a22o_1
Xwire279 net280 VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__clkbuf_1
X_23369_ _03232_ _03234_ _03231_ VGND VGND VPWR VPWR _03239_ sky130_fd_sc_hd__o21ba_1
Xmax_length2852 _06988_ VGND VGND VPWR VPWR net2852 sky130_fd_sc_hd__buf_1
XFILLER_0_132_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2874 net2875 VGND VGND VPWR VPWR net2874 sky130_fd_sc_hd__buf_1
X_13122_ net1585 _05394_ VGND VGND VPWR VPWR _05395_ sky130_fd_sc_hd__xnor2_1
X_25108_ net3033 VGND VGND VPWR VPWR _04850_ sky130_fd_sc_hd__buf_1
XFILLER_0_104_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13053_ _05323_ _05321_ _05322_ VGND VGND VPWR VPWR _05326_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17930_ net2145 net2143 VGND VGND VPWR VPWR _09781_ sky130_fd_sc_hd__nand2_1
X_25039_ net3738 _04790_ VGND VGND VPWR VPWR _04791_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17861_ net7069 _09709_ _09711_ net7105 net3258 VGND VGND VPWR VPWR _09712_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_84_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2140 _09815_ VGND VGND VPWR VPWR net2140 sky130_fd_sc_hd__clkbuf_1
Xwire2151 net2152 VGND VGND VPWR VPWR net2151 sky130_fd_sc_hd__clkbuf_1
X_19600_ net6029 _11387_ _11388_ net3864 VGND VGND VPWR VPWR _11437_ sky130_fd_sc_hd__o22a_1
X_16812_ _08796_ VGND VGND VPWR VPWR _00304_ sky130_fd_sc_hd__clkbuf_1
Xwire2162 net2163 VGND VGND VPWR VPWR net2162 sky130_fd_sc_hd__buf_1
XFILLER_0_108_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2173 _08951_ VGND VGND VPWR VPWR net2173 sky130_fd_sc_hd__buf_1
X_17792_ _09642_ VGND VGND VPWR VPWR _09643_ sky130_fd_sc_hd__buf_1
XFILLER_0_17_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2184 net2185 VGND VGND VPWR VPWR net2184 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1450 _09598_ VGND VGND VPWR VPWR net1450 sky130_fd_sc_hd__dlymetal6s2s_1
X_19531_ _11023_ net713 net712 net709 VGND VGND VPWR VPWR _11368_ sky130_fd_sc_hd__a31o_1
Xwire2195 net2196 VGND VGND VPWR VPWR net2195 sky130_fd_sc_hd__clkbuf_1
Xwire1461 _09304_ VGND VGND VPWR VPWR net1461 sky130_fd_sc_hd__buf_1
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16743_ _08760_ VGND VGND VPWR VPWR _00271_ sky130_fd_sc_hd__clkbuf_1
X_13955_ _06117_ net1597 VGND VGND VPWR VPWR _06220_ sky130_fd_sc_hd__nor2_1
Xwire1472 net1473 VGND VGND VPWR VPWR net1472 sky130_fd_sc_hd__clkbuf_1
Xwire1494 net1495 VGND VGND VPWR VPWR net1494 sky130_fd_sc_hd__buf_1
X_12906_ net7758 _04913_ net2315 VGND VGND VPWR VPWR _05179_ sky130_fd_sc_hd__and3_1
X_19462_ _11288_ _11298_ VGND VGND VPWR VPWR _11299_ sky130_fd_sc_hd__xor2_1
X_16674_ matmul0.matmul_stage_inst.mult2\[8\] matmul0.matmul_stage_inst.mult1\[8\]
+ VGND VGND VPWR VPWR _08707_ sky130_fd_sc_hd__xor2_1
X_13886_ net9180 net1126 net191 net1926 VGND VGND VPWR VPWR _00022_ sky130_fd_sc_hd__a22o_1
XFILLER_0_158_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18413_ net4245 net2932 VGND VGND VPWR VPWR _10263_ sky130_fd_sc_hd__nor2_1
XFILLER_0_185_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15625_ net2813 _07511_ VGND VGND VPWR VPWR _07697_ sky130_fd_sc_hd__nand2_1
X_12837_ net2975 _05059_ VGND VGND VPWR VPWR _05110_ sky130_fd_sc_hd__and2_1
X_19393_ net1192 _11229_ VGND VGND VPWR VPWR _11230_ sky130_fd_sc_hd__xor2_1
XFILLER_0_186_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18344_ _10193_ _10131_ _10194_ VGND VGND VPWR VPWR _10195_ sky130_fd_sc_hd__o21a_1
XFILLER_0_127_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15556_ net1273 _07496_ _07628_ VGND VGND VPWR VPWR _07629_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12768_ net7737 net2978 net2336 VGND VGND VPWR VPWR _05041_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14507_ _06685_ _06688_ VGND VGND VPWR VPWR _06689_ sky130_fd_sc_hd__nand2_1
XFILLER_0_182_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18275_ net1776 _10125_ VGND VGND VPWR VPWR _10126_ sky130_fd_sc_hd__xnor2_1
X_15487_ matmul0.matmul_stage_inst.mult1\[0\] net494 net2678 VGND VGND VPWR VPWR _07561_
+ sky130_fd_sc_hd__mux2_1
X_12699_ _04941_ _04971_ VGND VGND VPWR VPWR _04972_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17226_ net6791 _09172_ _09173_ _09162_ VGND VGND VPWR VPWR _09174_ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14438_ _06632_ matmul0.b_in\[11\] net896 VGND VGND VPWR VPWR _06633_ sky130_fd_sc_hd__mux2_1
Xinput10 angle_in[3] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_1
XFILLER_0_4_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput21 currA_in[13] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput32 currA_in[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput43 currB_in[4] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_1
Xinput54 currT_in[14] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17157_ net4039 _09097_ VGND VGND VPWR VPWR _09110_ sky130_fd_sc_hd__nor2_1
Xwire780 _05985_ VGND VGND VPWR VPWR net780 sky130_fd_sc_hd__clkbuf_2
Xinput65 periodTop[0] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_1
X_14369_ net7247 net1296 net2893 net5341 _06579_ VGND VGND VPWR VPWR _06580_ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput76 periodTop[5] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_1
Xwire791 _05141_ VGND VGND VPWR VPWR net791 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput87 pid_d_addr[15] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_1
Xinput98 pid_d_data[10] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16108_ net4074 _08171_ _08172_ net2816 _08173_ VGND VGND VPWR VPWR _08174_ sky130_fd_sc_hd__o221a_1
X_17088_ net7008 _09012_ _09044_ _09045_ VGND VGND VPWR VPWR _09046_ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16039_ net2712 _08053_ VGND VGND VPWR VPWR _08106_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19729_ net6066 _11562_ _11563_ VGND VGND VPWR VPWR _11564_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length7819 net7812 VGND VGND VPWR VPWR net7819 sky130_fd_sc_hd__buf_1
X_22740_ _02671_ VGND VGND VPWR VPWR _00603_ sky130_fd_sc_hd__clkbuf_1
X_22671_ pid_d.ki\[1\] net3010 net2994 pid_d.kp\[1\] VGND VGND VPWR VPWR _02622_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24410_ _04238_ _04244_ _04243_ VGND VGND VPWR VPWR _04268_ sky130_fd_sc_hd__a21oi_2
X_21622_ _01631_ _01633_ VGND VGND VPWR VPWR _01634_ sky130_fd_sc_hd__nand2_1
XFILLER_0_181_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25390_ clknet_leaf_83_clk _00273_ net8493 VGND VGND VPWR VPWR matmul0.b\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_191_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24341_ net4917 net4485 VGND VGND VPWR VPWR _04200_ sky130_fd_sc_hd__nand2_1
X_21553_ _01563_ _01564_ VGND VGND VPWR VPWR _01565_ sky130_fd_sc_hd__xor2_1
XFILLER_0_7_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7107 net7108 VGND VGND VPWR VPWR net7107 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_74_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7129 net7125 VGND VGND VPWR VPWR net7129 sky130_fd_sc_hd__buf_1
X_20504_ net1484 net2088 _12287_ _12290_ VGND VGND VPWR VPWR _12291_ sky130_fd_sc_hd__a211o_1
X_24272_ net4522 net4885 VGND VGND VPWR VPWR _04132_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6406 cordic0.slte0.opB\[9\] VGND VGND VPWR VPWR net6406 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21484_ _01366_ _01368_ _01496_ VGND VGND VPWR VPWR _01497_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_117_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6428 net6429 VGND VGND VPWR VPWR net6428 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23223_ net5012 net4738 VGND VGND VPWR VPWR _03093_ sky130_fd_sc_hd__nand2_2
XFILLER_0_16_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire6439 net6440 VGND VGND VPWR VPWR net6439 sky130_fd_sc_hd__clkbuf_1
X_20435_ net1487 _12229_ net3315 VGND VGND VPWR VPWR _12230_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5716 net5717 VGND VGND VPWR VPWR net5716 sky130_fd_sc_hd__buf_1
Xmax_length1403 _12142_ VGND VGND VPWR VPWR net1403 sky130_fd_sc_hd__buf_1
Xmax_length2159 net2160 VGND VGND VPWR VPWR net2159 sky130_fd_sc_hd__buf_1
Xwire5727 net5728 VGND VGND VPWR VPWR net5727 sky130_fd_sc_hd__clkbuf_1
Xwire5738 pid_d.mult0.b\[11\] VGND VGND VPWR VPWR net5738 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5749 net5744 VGND VGND VPWR VPWR net5749 sky130_fd_sc_hd__dlymetal6s2s_1
X_23154_ _03020_ _03023_ VGND VGND VPWR VPWR _03024_ sky130_fd_sc_hd__xnor2_2
X_20366_ _12164_ _12165_ net4055 VGND VGND VPWR VPWR _12166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length1469 _09068_ VGND VGND VPWR VPWR net1469 sky130_fd_sc_hd__clkbuf_1
X_22105_ _02108_ _02019_ _02110_ VGND VGND VPWR VPWR _02111_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23085_ _02871_ _02873_ VGND VGND VPWR VPWR _02955_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20297_ _12101_ _12102_ VGND VGND VPWR VPWR _12103_ sky130_fd_sc_hd__or2b_1
XFILLER_0_98_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22036_ _02039_ _02042_ VGND VGND VPWR VPWR _02043_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_98_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23987_ _03778_ _03850_ VGND VGND VPWR VPWR _03851_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13740_ _06004_ _06006_ _05872_ VGND VGND VPWR VPWR _06009_ sky130_fd_sc_hd__mux2_1
X_25726_ clknet_leaf_8_clk _00599_ net8553 VGND VGND VPWR VPWR pid_d.ki\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22938_ net205 net2030 VGND VGND VPWR VPWR _02827_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_196_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13671_ net7717 net1943 net2292 VGND VGND VPWR VPWR _05940_ sky130_fd_sc_hd__and3_2
X_25657_ clknet_leaf_25_clk _00530_ net8577 VGND VGND VPWR VPWR pid_d.curr_int\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_22869_ net4337 _02764_ _02765_ net472 net4359 VGND VGND VPWR VPWR _02766_ sky130_fd_sc_hd__a32o_1
XFILLER_0_183_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15410_ net6541 net6594 matmul0.matmul_stage_inst.e\[13\] VGND VGND VPWR VPWR _07484_
+ sky130_fd_sc_hd__o21a_1
X_24608_ _04409_ _04438_ _04408_ VGND VGND VPWR VPWR _04463_ sky130_fd_sc_hd__a21oi_1
X_12622_ net7314 _04892_ net3695 VGND VGND VPWR VPWR _04895_ sky130_fd_sc_hd__nand3_1
X_16390_ _08449_ _08451_ VGND VGND VPWR VPWR _08452_ sky130_fd_sc_hd__xnor2_1
X_25588_ clknet_leaf_99_clk _00461_ net8381 VGND VGND VPWR VPWR cordic0.cos\[8\] sky130_fd_sc_hd__dfrtp_1
Xwire8320 net8321 VGND VGND VPWR VPWR net8320 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8331 net8332 VGND VGND VPWR VPWR net8331 sky130_fd_sc_hd__buf_1
X_15341_ _07413_ _07414_ VGND VGND VPWR VPWR _07415_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_136_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24539_ _04373_ _04376_ _04394_ _04268_ _04266_ VGND VGND VPWR VPWR _04395_ sky130_fd_sc_hd__a221o_1
XFILLER_0_108_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4040 net4042 VGND VGND VPWR VPWR net4040 sky130_fd_sc_hd__buf_1
XFILLER_0_38_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4051 _08945_ VGND VGND VPWR VPWR net4051 sky130_fd_sc_hd__clkbuf_1
Xfanout6812 net6816 VGND VGND VPWR VPWR net6812 sky130_fd_sc_hd__buf_1
Xwire8364 net8365 VGND VGND VPWR VPWR net8364 sky130_fd_sc_hd__buf_1
Xwire7630 net7631 VGND VGND VPWR VPWR net7630 sky130_fd_sc_hd__buf_1
Xwire8375 net8376 VGND VGND VPWR VPWR net8375 sky130_fd_sc_hd__buf_1
X_18060_ _09909_ _09910_ VGND VGND VPWR VPWR _09911_ sky130_fd_sc_hd__xor2_1
Xfanout6834 net6849 VGND VGND VPWR VPWR net6834 sky130_fd_sc_hd__buf_1
XFILLER_0_0_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15272_ _07149_ net2768 VGND VGND VPWR VPWR _07346_ sky130_fd_sc_hd__nor2_1
Xwire8386 net8385 VGND VGND VPWR VPWR net8386 sky130_fd_sc_hd__buf_1
Xwire7652 net7653 VGND VGND VPWR VPWR net7652 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7663 net7664 VGND VGND VPWR VPWR net7663 sky130_fd_sc_hd__buf_1
XFILLER_0_124_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17011_ net3335 net3363 net4057 _08970_ _08971_ VGND VGND VPWR VPWR _08972_ sky130_fd_sc_hd__a221o_1
X_14223_ _06477_ _06480_ _06476_ VGND VGND VPWR VPWR _06481_ sky130_fd_sc_hd__a21oi_1
Xwire7674 net7670 VGND VGND VPWR VPWR net7674 sky130_fd_sc_hd__buf_1
Xfanout6878 net6880 VGND VGND VPWR VPWR net6878 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire7685 net7684 VGND VGND VPWR VPWR net7685 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire6940 net6941 VGND VGND VPWR VPWR net6940 sky130_fd_sc_hd__buf_1
XFILLER_0_46_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3372 net3373 VGND VGND VPWR VPWR net3372 sky130_fd_sc_hd__buf_1
Xwire7696 net7697 VGND VGND VPWR VPWR net7696 sky130_fd_sc_hd__clkbuf_1
Xwire6951 net6945 VGND VGND VPWR VPWR net6951 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire6962 net6961 VGND VGND VPWR VPWR net6962 sky130_fd_sc_hd__buf_1
XFILLER_0_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14154_ net7662 _06374_ _06414_ VGND VGND VPWR VPWR _06415_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6995 net6996 VGND VGND VPWR VPWR net6995 sky130_fd_sc_hd__buf_1
X_13105_ _05372_ net1138 VGND VGND VPWR VPWR _05378_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14085_ _06298_ _06303_ _06347_ VGND VGND VPWR VPWR _06348_ sky130_fd_sc_hd__o21a_1
X_18962_ _10797_ _10798_ VGND VGND VPWR VPWR _10799_ sky130_fd_sc_hd__xnor2_1
X_13036_ _05307_ net735 VGND VGND VPWR VPWR _05309_ sky130_fd_sc_hd__or2_1
X_17913_ net1781 _09763_ _09667_ VGND VGND VPWR VPWR _09764_ sky130_fd_sc_hd__a21oi_1
X_18893_ _10705_ net1194 VGND VGND VPWR VPWR _10734_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17844_ net7132 _09694_ VGND VGND VPWR VPWR _09695_ sky130_fd_sc_hd__nand2_1
X_17775_ net7061 _09625_ VGND VGND VPWR VPWR _09626_ sky130_fd_sc_hd__nand2_1
XFILLER_0_191_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14987_ net4195 net4193 VGND VGND VPWR VPWR _07061_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1280 net1281 VGND VGND VPWR VPWR net1280 sky130_fd_sc_hd__clkbuf_2
X_16726_ _08751_ VGND VGND VPWR VPWR _00263_ sky130_fd_sc_hd__clkbuf_1
X_19514_ _11346_ _11350_ VGND VGND VPWR VPWR _11351_ sky130_fd_sc_hd__xnor2_1
Xwire1291 _06852_ VGND VGND VPWR VPWR net1291 sky130_fd_sc_hd__clkbuf_1
X_13938_ net836 _06203_ VGND VGND VPWR VPWR _06204_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19445_ _11266_ _11280_ _11281_ VGND VGND VPWR VPWR _11282_ sky130_fd_sc_hd__or3_1
X_16657_ matmul0.matmul_stage_inst.mult1\[5\] VGND VGND VPWR VPWR _08692_ sky130_fd_sc_hd__inv_2
X_13869_ _06125_ _06135_ VGND VGND VPWR VPWR _06136_ sky130_fd_sc_hd__xor2_1
XFILLER_0_14_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15608_ _07674_ _07679_ VGND VGND VPWR VPWR _07680_ sky130_fd_sc_hd__xnor2_1
X_19376_ _11209_ _11210_ _11211_ _11212_ VGND VGND VPWR VPWR _11213_ sky130_fd_sc_hd__o22a_1
XFILLER_0_85_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16588_ _08641_ VGND VGND VPWR VPWR _00235_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_173_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18327_ _10175_ net2543 VGND VGND VPWR VPWR _10178_ sky130_fd_sc_hd__xnor2_1
X_15539_ _07513_ _07521_ _07611_ VGND VGND VPWR VPWR _07612_ sky130_fd_sc_hd__o21a_1
Xfanout8781 net8790 VGND VGND VPWR VPWR net8781 sky130_fd_sc_hd__buf_2
Xfanout8792 net8839 VGND VGND VPWR VPWR net8792 sky130_fd_sc_hd__buf_1
XFILLER_0_151_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18258_ net7032 net7124 net7064 VGND VGND VPWR VPWR _10109_ sky130_fd_sc_hd__and3b_1
XFILLER_0_8_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17209_ _09154_ _09155_ net2587 VGND VGND VPWR VPWR _09159_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18189_ net6953 net6922 VGND VGND VPWR VPWR _10040_ sky130_fd_sc_hd__and2b_2
X_20220_ net8100 _12040_ VGND VGND VPWR VPWR _12041_ sky130_fd_sc_hd__xor2_1
XFILLER_0_142_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20151_ _11971_ _11976_ _11977_ VGND VGND VPWR VPWR _11978_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2909 net2910 VGND VGND VPWR VPWR net2909 sky130_fd_sc_hd__clkbuf_1
X_20082_ _11878_ _11909_ VGND VGND VPWR VPWR _11911_ sky130_fd_sc_hd__nor2_1
XFILLER_0_176_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23910_ pid_q.curr_int\[6\] pid_q.prev_int\[6\] VGND VGND VPWR VPWR _03774_ sky130_fd_sc_hd__xor2_1
X_24890_ _04684_ net4556 net1997 VGND VGND VPWR VPWR _04685_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23841_ _03701_ net2412 _03702_ _03704_ net3741 VGND VGND VPWR VPWR _03706_ sky130_fd_sc_hd__a2111oi_2
XFILLER_0_19_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length7616 net7617 VGND VGND VPWR VPWR net7616 sky130_fd_sc_hd__buf_1
X_23772_ net1164 _03637_ VGND VGND VPWR VPWR _03638_ sky130_fd_sc_hd__xor2_1
X_20984_ _00980_ _00981_ VGND VGND VPWR VPWR _01000_ sky130_fd_sc_hd__nand2_1
XFILLER_0_192_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25511_ clknet_leaf_42_clk _00391_ net8777 VGND VGND VPWR VPWR svm0.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length6915 net6916 VGND VGND VPWR VPWR net6915 sky130_fd_sc_hd__buf_1
X_22723_ _02655_ _02656_ net8084 _02658_ VGND VGND VPWR VPWR _02659_ sky130_fd_sc_hd__or4_1
Xmax_length6926 net6927 VGND VGND VPWR VPWR net6926 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_94_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6937 net6938 VGND VGND VPWR VPWR net6937 sky130_fd_sc_hd__clkbuf_1
Xmax_length6959 net6960 VGND VGND VPWR VPWR net6959 sky130_fd_sc_hd__clkbuf_1
X_25442_ clknet_leaf_113_clk _00325_ net8338 VGND VGND VPWR VPWR cordic0.vec\[1\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_22654_ net5751 net3085 VGND VGND VPWR VPWR _02612_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21605_ _01554_ _01616_ VGND VGND VPWR VPWR _01617_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22585_ net7317 net7306 _02554_ VGND VGND VPWR VPWR _02564_ sky130_fd_sc_hd__or3_1
X_25373_ clknet_leaf_63_clk _00256_ net8708 VGND VGND VPWR VPWR matmul0.alpha_pass\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_164_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24324_ net7506 _04182_ _04183_ VGND VGND VPWR VPWR _04184_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21536_ _01420_ net757 VGND VGND VPWR VPWR _01548_ sky130_fd_sc_hd__nor2_1
Xwire6214 net6212 VGND VGND VPWR VPWR net6214 sky130_fd_sc_hd__buf_1
Xwire6225 net6226 VGND VGND VPWR VPWR net6225 sky130_fd_sc_hd__buf_1
XFILLER_0_62_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6236 net6238 VGND VGND VPWR VPWR net6236 sky130_fd_sc_hd__clkbuf_1
Xwire5502 net5503 VGND VGND VPWR VPWR net5502 sky130_fd_sc_hd__clkbuf_2
X_24255_ net7523 _04042_ net269 net7467 net536 VGND VGND VPWR VPWR _04116_ sky130_fd_sc_hd__a221o_1
X_21467_ net1727 _01479_ VGND VGND VPWR VPWR _01480_ sky130_fd_sc_hd__xor2_1
XFILLER_0_50_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5513 net5514 VGND VGND VPWR VPWR net5513 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_177_Right_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5524 net5525 VGND VGND VPWR VPWR net5524 sky130_fd_sc_hd__buf_1
X_23206_ net5157 net4723 VGND VGND VPWR VPWR _03076_ sky130_fd_sc_hd__nand2_1
Xwire5535 net5536 VGND VGND VPWR VPWR net5535 sky130_fd_sc_hd__buf_1
X_20418_ _12214_ VGND VGND VPWR VPWR _00493_ sky130_fd_sc_hd__clkbuf_1
Xwire4801 net4802 VGND VGND VPWR VPWR net4801 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5546 net5547 VGND VGND VPWR VPWR net5546 sky130_fd_sc_hd__buf_1
Xwire4812 net4810 VGND VGND VPWR VPWR net4812 sky130_fd_sc_hd__buf_1
X_24186_ net739 _04046_ net694 VGND VGND VPWR VPWR _04047_ sky130_fd_sc_hd__a21bo_1
X_21398_ net5455 _00820_ _00821_ _01304_ VGND VGND VPWR VPWR _01412_ sky130_fd_sc_hd__o31a_1
Xwire5557 net5559 VGND VGND VPWR VPWR net5557 sky130_fd_sc_hd__buf_1
Xwire4823 net4824 VGND VGND VPWR VPWR net4823 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4834 net4835 VGND VGND VPWR VPWR net4834 sky130_fd_sc_hd__buf_1
Xwire5579 net5575 VGND VGND VPWR VPWR net5579 sky130_fd_sc_hd__buf_1
X_23137_ _03006_ net1031 _02987_ VGND VGND VPWR VPWR _03007_ sky130_fd_sc_hd__nor3_1
Xwire4845 net4846 VGND VGND VPWR VPWR net4845 sky130_fd_sc_hd__buf_1
X_20349_ _12140_ _12149_ _12148_ VGND VGND VPWR VPWR _12151_ sky130_fd_sc_hd__a21o_1
Xwire4856 net4857 VGND VGND VPWR VPWR net4856 sky130_fd_sc_hd__clkbuf_1
Xwire4867 net4862 VGND VGND VPWR VPWR net4867 sky130_fd_sc_hd__buf_1
XFILLER_0_102_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4889 net4890 VGND VGND VPWR VPWR net4889 sky130_fd_sc_hd__buf_1
XFILLER_0_101_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23068_ _02876_ _02878_ _02877_ VGND VGND VPWR VPWR _02938_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_179_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22019_ net5693 net5498 VGND VGND VPWR VPWR _02026_ sky130_fd_sc_hd__nand2_1
X_14910_ _06969_ VGND VGND VPWR VPWR _06984_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_175_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15890_ _07949_ _07957_ VGND VGND VPWR VPWR _07959_ sky130_fd_sc_hd__nand2_1
X_14841_ _06937_ VGND VGND VPWR VPWR _00192_ sky130_fd_sc_hd__clkbuf_1
X_17560_ svm0.tC\[9\] VGND VGND VPWR VPWR _09442_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14772_ matmul0.sin\[10\] _06898_ VGND VGND VPWR VPWR _06899_ sky130_fd_sc_hd__xor2_1
X_16511_ _08510_ _08519_ net977 VGND VGND VPWR VPWR _08571_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13723_ net621 _05991_ VGND VGND VPWR VPWR _05992_ sky130_fd_sc_hd__xnor2_1
X_25709_ clknet_leaf_4_clk _00582_ net8562 VGND VGND VPWR VPWR pid_d.mult0.b\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_17491_ net4027 _09380_ VGND VGND VPWR VPWR _09381_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19230_ net6201 _11060_ _11065_ _11066_ VGND VGND VPWR VPWR _11067_ sky130_fd_sc_hd__o211a_1
X_16442_ net1086 _08502_ net1078 VGND VGND VPWR VPWR _08503_ sky130_fd_sc_hd__o21a_1
X_13654_ _05793_ _05922_ _05923_ VGND VGND VPWR VPWR _05924_ sky130_fd_sc_hd__a21o_1
XFILLER_0_155_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12605_ _04881_ VGND VGND VPWR VPWR _04882_ sky130_fd_sc_hd__clkbuf_1
X_19161_ net6147 net6101 net3878 VGND VGND VPWR VPWR _10998_ sky130_fd_sc_hd__and3_1
XFILLER_0_183_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16373_ _08418_ net1247 _08434_ VGND VGND VPWR VPWR _08435_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_184_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13585_ _05852_ _05855_ VGND VGND VPWR VPWR _05856_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18112_ _09860_ net2550 _09881_ VGND VGND VPWR VPWR _09963_ sky130_fd_sc_hd__or3_1
Xwire8150 net43 VGND VGND VPWR VPWR net8150 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_186_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8161 net8162 VGND VGND VPWR VPWR net8161 sky130_fd_sc_hd__clkbuf_1
X_15324_ net1868 _07397_ VGND VGND VPWR VPWR _07398_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_183_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19092_ net6246 _10927_ _10928_ VGND VGND VPWR VPWR _10929_ sky130_fd_sc_hd__a21oi_1
Xwire8172 net8173 VGND VGND VPWR VPWR net8172 sky130_fd_sc_hd__clkbuf_1
Xwire8183 net8184 VGND VGND VPWR VPWR net8183 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_170_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8194 net8195 VGND VGND VPWR VPWR net8194 sky130_fd_sc_hd__clkbuf_1
X_18043_ _09860_ net2550 VGND VGND VPWR VPWR _09894_ sky130_fd_sc_hd__xor2_2
Xwire7460 net7461 VGND VGND VPWR VPWR net7460 sky130_fd_sc_hd__buf_1
X_15255_ _07327_ net990 _07328_ net2779 net2705 VGND VGND VPWR VPWR _07329_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_81_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7482 net7479 VGND VGND VPWR VPWR net7482 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_83_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6686 svm0.counter\[14\] VGND VGND VPWR VPWR net6686 sky130_fd_sc_hd__clkbuf_2
Xfanout5941 pid_d.mult0.b\[1\] VGND VGND VPWR VPWR net5941 sky130_fd_sc_hd__clkbuf_1
Xfanout6697 svm0.counter\[12\] VGND VGND VPWR VPWR net6697 sky130_fd_sc_hd__buf_1
Xwire7493 net7494 VGND VGND VPWR VPWR net7493 sky130_fd_sc_hd__clkbuf_1
X_14206_ _06416_ _06450_ _06464_ _06411_ VGND VGND VPWR VPWR _06465_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_144_Right_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire6770 net6769 VGND VGND VPWR VPWR net6770 sky130_fd_sc_hd__buf_1
X_15186_ _07255_ _07257_ _07259_ VGND VGND VPWR VPWR _07260_ sky130_fd_sc_hd__o21a_1
Xwire6781 net6780 VGND VGND VPWR VPWR net6781 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_22_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14137_ _06366_ _06398_ VGND VGND VPWR VPWR _06399_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19994_ _11783_ VGND VGND VPWR VPWR _11825_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14068_ _06329_ _06330_ VGND VGND VPWR VPWR _06331_ sky130_fd_sc_hd__xnor2_1
X_18945_ net9101 net2121 net1450 _10783_ VGND VGND VPWR VPWR _00451_ sky130_fd_sc_hd__a31o_1
XFILLER_0_183_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13019_ net7933 _05288_ _05291_ net1596 VGND VGND VPWR VPWR _05292_ sky130_fd_sc_hd__a211o_1
X_18876_ _10716_ _10717_ VGND VGND VPWR VPWR _10718_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17827_ net2561 VGND VGND VPWR VPWR _09678_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17758_ net6996 net7021 VGND VGND VPWR VPWR _09609_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16709_ net7375 matmul0.matmul_stage_inst.mult1\[13\] VGND VGND VPWR VPWR _08737_
+ sky130_fd_sc_hd__xor2_1
X_17689_ net6701 _09567_ _09568_ VGND VGND VPWR VPWR _09569_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19428_ _10851_ _11264_ VGND VGND VPWR VPWR _11265_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_162_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19359_ _11152_ _11188_ _11195_ VGND VGND VPWR VPWR _11196_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_174_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22370_ net1715 _01964_ VGND VGND VPWR VPWR _02373_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21321_ net4384 _01249_ net561 net4320 _01335_ VGND VGND VPWR VPWR _01336_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24040_ net4652 net4815 _03902_ VGND VGND VPWR VPWR _03903_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_111_Right_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21252_ _01265_ _01266_ VGND VGND VPWR VPWR _01267_ sky130_fd_sc_hd__xor2_1
Xwire4108 net4109 VGND VGND VPWR VPWR net4108 sky130_fd_sc_hd__buf_1
XFILLER_0_40_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20203_ net244 _11967_ VGND VGND VPWR VPWR _12028_ sky130_fd_sc_hd__nand2_1
X_21183_ net5634 net5882 _01172_ _01198_ VGND VGND VPWR VPWR _01199_ sky130_fd_sc_hd__a31o_1
Xwire3407 net3408 VGND VGND VPWR VPWR net3407 sky130_fd_sc_hd__buf_1
XFILLER_0_25_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3418 net3419 VGND VGND VPWR VPWR net3418 sky130_fd_sc_hd__buf_1
Xwire3429 net3430 VGND VGND VPWR VPWR net3429 sky130_fd_sc_hd__buf_1
X_20134_ _11846_ _11960_ _11961_ VGND VGND VPWR VPWR _11962_ sky130_fd_sc_hd__o21a_1
Xwire2706 _07309_ VGND VGND VPWR VPWR net2706 sky130_fd_sc_hd__clkbuf_1
Xwire2717 net2718 VGND VGND VPWR VPWR net2717 sky130_fd_sc_hd__buf_1
XFILLER_0_99_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2728 _07241_ VGND VGND VPWR VPWR net2728 sky130_fd_sc_hd__clkbuf_1
Xwire2739 _07226_ VGND VGND VPWR VPWR net2739 sky130_fd_sc_hd__clkbuf_1
X_24942_ net8866 net8882 VGND VGND VPWR VPWR _04722_ sky130_fd_sc_hd__and2b_1
X_20065_ _11892_ net2493 VGND VGND VPWR VPWR _11894_ sky130_fd_sc_hd__or2_1
X_24873_ _04673_ VGND VGND VPWR VPWR _00734_ sky130_fd_sc_hd__clkbuf_1
X_23824_ _03589_ _03591_ VGND VGND VPWR VPWR _03689_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length7435 matmul0.matmul_stage_inst.b\[1\] VGND VGND VPWR VPWR net7435 sky130_fd_sc_hd__clkbuf_1
X_23755_ _03489_ _03491_ _03490_ VGND VGND VPWR VPWR _03621_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_67_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20967_ _00979_ _00982_ VGND VGND VPWR VPWR _00983_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_49_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22706_ _02645_ net5436 net3094 VGND VGND VPWR VPWR _02646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23686_ _03547_ _03551_ VGND VGND VPWR VPWR _03553_ sky130_fd_sc_hd__nand2_1
XFILLER_0_166_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6778 net6779 VGND VGND VPWR VPWR net6778 sky130_fd_sc_hd__clkbuf_1
X_20898_ _00906_ _00910_ _00891_ VGND VGND VPWR VPWR _00914_ sky130_fd_sc_hd__a21o_1
X_25425_ clknet_leaf_91_clk _00308_ net8428 VGND VGND VPWR VPWR matmul0.cos\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_181_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22637_ net3081 net3092 VGND VGND VPWR VPWR _02603_ sky130_fd_sc_hd__nor2_1
XFILLER_0_165_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13370_ net7947 net1935 VGND VGND VPWR VPWR _05643_ sky130_fd_sc_hd__nand2_1
X_25356_ clknet_leaf_85_clk _00239_ net8513 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult2\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_22568_ net7369 net7352 net7343 VGND VGND VPWR VPWR _02550_ sky130_fd_sc_hd__o21ai_1
Xwire6000 net6001 VGND VGND VPWR VPWR net6000 sky130_fd_sc_hd__buf_1
XFILLER_0_152_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24307_ net692 _04102_ _04101_ VGND VGND VPWR VPWR _04167_ sky130_fd_sc_hd__a21o_1
Xwire6022 net6018 VGND VGND VPWR VPWR net6022 sky130_fd_sc_hd__buf_1
X_21519_ _01342_ _01527_ _01530_ _01531_ VGND VGND VPWR VPWR _01532_ sky130_fd_sc_hd__a211o_1
Xwire6033 net6031 VGND VGND VPWR VPWR net6033 sky130_fd_sc_hd__dlymetal6s2s_1
X_25287_ clknet_leaf_88_clk _00170_ net8444 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.d\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout4503 net4509 VGND VGND VPWR VPWR net4503 sky130_fd_sc_hd__buf_1
X_22499_ _02438_ _02499_ VGND VGND VPWR VPWR _02500_ sky130_fd_sc_hd__nor2_1
Xfanout4514 net4524 VGND VGND VPWR VPWR net4514 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_134_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5310 net5313 VGND VGND VPWR VPWR net5310 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6055 net6056 VGND VGND VPWR VPWR net6055 sky130_fd_sc_hd__buf_1
Xfanout4525 pid_q.mult0.a\[13\] VGND VGND VPWR VPWR net4525 sky130_fd_sc_hd__buf_1
Xwire5321 net5322 VGND VGND VPWR VPWR net5321 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6066 net6067 VGND VGND VPWR VPWR net6066 sky130_fd_sc_hd__buf_1
X_15040_ _07064_ _07113_ VGND VGND VPWR VPWR _07114_ sky130_fd_sc_hd__xnor2_1
X_24238_ net1015 net1658 VGND VGND VPWR VPWR _04099_ sky130_fd_sc_hd__nand2_1
Xwire5332 pid_d.out\[13\] VGND VGND VPWR VPWR net5332 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5343 net5344 VGND VGND VPWR VPWR net5343 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6099 net6096 VGND VGND VPWR VPWR net6099 sky130_fd_sc_hd__buf_1
Xwire4620 net4621 VGND VGND VPWR VPWR net4620 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5365 pid_d.out\[2\] VGND VGND VPWR VPWR net5365 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4631 net4632 VGND VGND VPWR VPWR net4631 sky130_fd_sc_hd__buf_1
Xwire5376 net5377 VGND VGND VPWR VPWR net5376 sky130_fd_sc_hd__buf_1
Xwire4642 net4639 VGND VGND VPWR VPWR net4642 sky130_fd_sc_hd__clkbuf_1
X_24169_ _04029_ _03948_ _04030_ VGND VGND VPWR VPWR _04031_ sky130_fd_sc_hd__a21o_1
Xwire5387 pid_d.mult0.a\[15\] VGND VGND VPWR VPWR net5387 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4653 net4655 VGND VGND VPWR VPWR net4653 sky130_fd_sc_hd__clkbuf_1
Xwire4664 net4665 VGND VGND VPWR VPWR net4664 sky130_fd_sc_hd__buf_1
Xwire4675 net4676 VGND VGND VPWR VPWR net4675 sky130_fd_sc_hd__buf_1
Xwire3930 net3931 VGND VGND VPWR VPWR net3930 sky130_fd_sc_hd__buf_1
Xwire4686 net4680 VGND VGND VPWR VPWR net4686 sky130_fd_sc_hd__clkbuf_1
X_16991_ net2612 net2606 VGND VGND VPWR VPWR _08953_ sky130_fd_sc_hd__or2_1
Xwire3941 _09934_ VGND VGND VPWR VPWR net3941 sky130_fd_sc_hd__buf_1
Xwire4697 net4698 VGND VGND VPWR VPWR net4697 sky130_fd_sc_hd__buf_1
Xwire3952 _09808_ VGND VGND VPWR VPWR net3952 sky130_fd_sc_hd__clkbuf_2
Xwire3974 net3975 VGND VGND VPWR VPWR net3974 sky130_fd_sc_hd__clkbuf_1
X_18730_ net6877 _10533_ _10534_ VGND VGND VPWR VPWR _10575_ sky130_fd_sc_hd__mux2_1
X_15942_ matmul0.matmul_stage_inst.mult1\[5\] net389 _07560_ VGND VGND VPWR VPWR _08011_
+ sky130_fd_sc_hd__mux2_1
Xwire3985 _09661_ VGND VGND VPWR VPWR net3985 sky130_fd_sc_hd__clkbuf_1
Xwire3996 _09617_ VGND VGND VPWR VPWR net3996 sky130_fd_sc_hd__buf_1
X_18661_ net422 _10505_ _10507_ net714 net3923 VGND VGND VPWR VPWR _10508_ sky130_fd_sc_hd__a221o_1
X_15873_ _07846_ net3390 _07941_ VGND VGND VPWR VPWR _07942_ sky130_fd_sc_hd__o21a_1
XFILLER_0_92_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17612_ _09488_ _09489_ _09492_ VGND VGND VPWR VPWR _09493_ sky130_fd_sc_hd__and3b_1
X_14824_ matmul0.a\[1\] matmul0.matmul_stage_inst.e\[1\] net3610 VGND VGND VPWR VPWR
+ _06929_ sky130_fd_sc_hd__mux2_1
X_18592_ net2128 _10439_ VGND VGND VPWR VPWR _10440_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17543_ svm0.tC\[12\] VGND VGND VPWR VPWR _09425_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length8681 net8682 VGND VGND VPWR VPWR net8681 sky130_fd_sc_hd__buf_1
X_14755_ _06826_ net7153 _06839_ VGND VGND VPWR VPWR _06886_ sky130_fd_sc_hd__nand3_1
X_13706_ net7660 net2332 net2326 VGND VGND VPWR VPWR _05975_ sky130_fd_sc_hd__and3_1
XFILLER_0_196_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17474_ net4014 _09360_ VGND VGND VPWR VPWR _09366_ sky130_fd_sc_hd__nand2_1
X_14686_ net9031 net2868 net2262 net2863 VGND VGND VPWR VPWR _00140_ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19213_ net6335 net6287 VGND VGND VPWR VPWR _11050_ sky130_fd_sc_hd__or2b_1
X_16425_ _08485_ _08486_ net303 VGND VGND VPWR VPWR _08487_ sky130_fd_sc_hd__mux2_1
X_13637_ net7657 net1150 VGND VGND VPWR VPWR _05907_ sky130_fd_sc_hd__nand2_1
XFILLER_0_183_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19144_ net2522 net2521 VGND VGND VPWR VPWR _10981_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16356_ net2691 net2210 _08313_ VGND VGND VPWR VPWR _08419_ sky130_fd_sc_hd__and3_1
X_13568_ _05708_ _05837_ _05838_ VGND VGND VPWR VPWR _05839_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15307_ net3501 _07066_ VGND VGND VPWR VPWR _07381_ sky130_fd_sc_hd__nor2_1
Xfanout6450 state\[1\] VGND VGND VPWR VPWR net6450 sky130_fd_sc_hd__clkbuf_1
X_19075_ net6260 net6311 VGND VGND VPWR VPWR _10912_ sky130_fd_sc_hd__or2_1
X_16287_ _08339_ _08350_ VGND VGND VPWR VPWR _08351_ sky130_fd_sc_hd__xnor2_2
X_13499_ _05770_ _05771_ VGND VGND VPWR VPWR _05772_ sky130_fd_sc_hd__nor2_1
XFILLER_0_180_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18026_ net6990 net7035 VGND VGND VPWR VPWR _09877_ sky130_fd_sc_hd__nand2_1
Xwire7290 net7291 VGND VGND VPWR VPWR net7290 sky130_fd_sc_hd__clkbuf_1
X_15238_ net1880 _07311_ VGND VGND VPWR VPWR _07312_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_140_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15169_ _07193_ _07242_ VGND VGND VPWR VPWR _07243_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_157_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19977_ _11806_ _11807_ VGND VGND VPWR VPWR _11808_ sky130_fd_sc_hd__and2_1
XFILLER_0_158_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18928_ net245 _10767_ VGND VGND VPWR VPWR _10768_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18859_ _10686_ _10689_ _10700_ net2125 VGND VGND VPWR VPWR _10701_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_173_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21870_ net1048 net1172 VGND VGND VPWR VPWR _01879_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length6008 net6009 VGND VGND VPWR VPWR net6008 sky130_fd_sc_hd__buf_1
X_20821_ _00834_ net1736 VGND VGND VPWR VPWR _00837_ sky130_fd_sc_hd__xor2_1
XFILLER_0_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23540_ _03397_ _03407_ VGND VGND VPWR VPWR _03408_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20752_ _12521_ _12522_ VGND VGND VPWR VPWR _12523_ sky130_fd_sc_hd__nand2_1
Xwire8908 net8904 VGND VGND VPWR VPWR net8908 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8919 net8920 VGND VGND VPWR VPWR net8919 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23471_ _03338_ _03339_ VGND VGND VPWR VPWR _03340_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_135_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20683_ _12454_ _12457_ VGND VGND VPWR VPWR _12459_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25210_ clknet_leaf_64_clk _00099_ net8670 VGND VGND VPWR VPWR matmul0.op_in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_22422_ _02420_ _02423_ VGND VGND VPWR VPWR _02424_ sky130_fd_sc_hd__xnor2_2
Xwire609 net610 VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length218 net219 VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__buf_1
XFILLER_0_17_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25141_ clknet_leaf_50_clk _00030_ net8757 VGND VGND VPWR VPWR svm0.tC\[13\] sky130_fd_sc_hd__dfrtp_1
X_22353_ _02352_ _02355_ VGND VGND VPWR VPWR _02356_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_61_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21304_ _00868_ _01316_ _01318_ VGND VGND VPWR VPWR _01319_ sky130_fd_sc_hd__o21a_1
X_22284_ _02284_ _02287_ VGND VGND VPWR VPWR _02288_ sky130_fd_sc_hd__xnor2_1
X_25072_ _04817_ _04818_ VGND VGND VPWR VPWR _04819_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24023_ net5011 _03819_ VGND VGND VPWR VPWR _03886_ sky130_fd_sc_hd__xor2_1
XFILLER_0_41_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21235_ _00935_ _01238_ VGND VGND VPWR VPWR _01250_ sky130_fd_sc_hd__and2_1
Xhold240 pid_q.curr_error\[10\] VGND VGND VPWR VPWR net9193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 svm0.tB\[2\] VGND VGND VPWR VPWR net9204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 pid_d.prev_int\[7\] VGND VGND VPWR VPWR net9215 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3215 _10792_ VGND VGND VPWR VPWR net3215 sky130_fd_sc_hd__buf_1
Xhold273 matmul0.b_in\[4\] VGND VGND VPWR VPWR net9226 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3226 net3227 VGND VGND VPWR VPWR net3226 sky130_fd_sc_hd__clkbuf_1
X_21166_ net5882 _01181_ VGND VGND VPWR VPWR _01182_ sky130_fd_sc_hd__nand2_1
Xwire3237 _09851_ VGND VGND VPWR VPWR net3237 sky130_fd_sc_hd__buf_1
Xhold284 matmul0.b\[13\] VGND VGND VPWR VPWR net9237 sky130_fd_sc_hd__dlygate4sd3_1
Xwire2503 _11491_ VGND VGND VPWR VPWR net2503 sky130_fd_sc_hd__clkbuf_1
Xwire3248 net3249 VGND VGND VPWR VPWR net3248 sky130_fd_sc_hd__buf_1
Xwire2514 net2515 VGND VGND VPWR VPWR net2514 sky130_fd_sc_hd__clkbuf_1
Xwire3259 _09638_ VGND VGND VPWR VPWR net3259 sky130_fd_sc_hd__buf_1
Xwire2525 _10899_ VGND VGND VPWR VPWR net2525 sky130_fd_sc_hd__dlymetal6s2s_1
X_20117_ net6006 _11648_ VGND VGND VPWR VPWR _11945_ sky130_fd_sc_hd__nand2_1
Xwire2536 _10770_ VGND VGND VPWR VPWR net2536 sky130_fd_sc_hd__clkbuf_1
Xwire1802 net1803 VGND VGND VPWR VPWR net1802 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2547 _10042_ VGND VGND VPWR VPWR net2547 sky130_fd_sc_hd__buf_1
X_21097_ _01063_ _01058_ VGND VGND VPWR VPWR _01113_ sky130_fd_sc_hd__xnor2_1
Xwire2558 _09691_ VGND VGND VPWR VPWR net2558 sky130_fd_sc_hd__buf_1
Xwire1813 net1814 VGND VGND VPWR VPWR net1813 sky130_fd_sc_hd__buf_1
Xwire1824 net1826 VGND VGND VPWR VPWR net1824 sky130_fd_sc_hd__buf_1
Xwire2569 net2570 VGND VGND VPWR VPWR net2569 sky130_fd_sc_hd__buf_1
X_24925_ pid_q.ki\[4\] _04710_ net1362 VGND VGND VPWR VPWR _04711_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1835 net1836 VGND VGND VPWR VPWR net1835 sky130_fd_sc_hd__buf_1
X_20048_ _11848_ _11870_ _11871_ VGND VGND VPWR VPWR _11877_ sky130_fd_sc_hd__o21ba_1
Xwire1846 _07901_ VGND VGND VPWR VPWR net1846 sky130_fd_sc_hd__buf_1
Xwire1857 net1858 VGND VGND VPWR VPWR net1857 sky130_fd_sc_hd__buf_1
Xwire1868 _07392_ VGND VGND VPWR VPWR net1868 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1879 _07290_ VGND VGND VPWR VPWR net1879 sky130_fd_sc_hd__buf_1
X_24856_ _04661_ VGND VGND VPWR VPWR _00729_ sky130_fd_sc_hd__clkbuf_1
X_12870_ net736 _05142_ VGND VGND VPWR VPWR _05143_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23807_ _03670_ _03580_ _03671_ VGND VGND VPWR VPWR _03672_ sky130_fd_sc_hd__o21a_1
X_24787_ _04608_ _04607_ _04612_ VGND VGND VPWR VPWR _04613_ sky130_fd_sc_hd__o21a_1
X_21999_ net471 _02006_ VGND VGND VPWR VPWR _02007_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14540_ net3639 VGND VGND VPWR VPWR _06719_ sky130_fd_sc_hd__clkbuf_1
X_23738_ _03600_ _03603_ VGND VGND VPWR VPWR _03604_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14471_ net7361 net5305 VGND VGND VPWR VPWR _06658_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23669_ _03530_ _03535_ VGND VGND VPWR VPWR _03536_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length5852 net5853 VGND VGND VPWR VPWR net5852 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16210_ _08187_ _08188_ _08189_ VGND VGND VPWR VPWR _08275_ sky130_fd_sc_hd__a21o_1
X_13422_ _05693_ _05694_ VGND VGND VPWR VPWR _05695_ sky130_fd_sc_hd__and2b_1
X_25408_ clknet_leaf_80_clk _00291_ net8489 VGND VGND VPWR VPWR matmul0.a\[11\] sky130_fd_sc_hd__dfrtp_1
X_17190_ _09139_ _09140_ net6839 VGND VGND VPWR VPWR _09141_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16141_ _08186_ _08206_ VGND VGND VPWR VPWR _08207_ sky130_fd_sc_hd__or2_1
X_13353_ _05612_ _05625_ VGND VGND VPWR VPWR _05626_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25339_ clknet_leaf_85_clk _00222_ net8506 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16072_ _08034_ net1261 _08032_ VGND VGND VPWR VPWR _08139_ sky130_fd_sc_hd__a21bo_1
Xfanout5067 net5074 VGND VGND VPWR VPWR net5067 sky130_fd_sc_hd__clkbuf_1
X_13284_ net3688 net2303 net1321 VGND VGND VPWR VPWR _05557_ sky130_fd_sc_hd__and3_1
XFILLER_0_87_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5140 net5139 VGND VGND VPWR VPWR net5140 sky130_fd_sc_hd__buf_1
Xwire5151 net5152 VGND VGND VPWR VPWR net5151 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19900_ _11667_ net708 _11715_ _11731_ VGND VGND VPWR VPWR _11732_ sky130_fd_sc_hd__o31a_1
X_15023_ net3511 net3506 net4163 net4159 VGND VGND VPWR VPWR _07097_ sky130_fd_sc_hd__o22a_1
Xwire5162 net5163 VGND VGND VPWR VPWR net5162 sky130_fd_sc_hd__buf_1
XFILLER_0_121_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5173 pid_q.curr_int\[13\] VGND VGND VPWR VPWR net5173 sky130_fd_sc_hd__buf_1
Xwire5184 pid_q.curr_int\[0\] VGND VGND VPWR VPWR net5184 sky130_fd_sc_hd__buf_1
XFILLER_0_20_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5195 net5196 VGND VGND VPWR VPWR net5195 sky130_fd_sc_hd__buf_1
Xwire4450 net4451 VGND VGND VPWR VPWR net4450 sky130_fd_sc_hd__clkbuf_1
Xwire4461 pid_q.out\[3\] VGND VGND VPWR VPWR net4461 sky130_fd_sc_hd__clkbuf_1
X_19831_ _11543_ _11662_ _11664_ VGND VGND VPWR VPWR _11665_ sky130_fd_sc_hd__o21ai_1
Xwire4472 net4473 VGND VGND VPWR VPWR net4472 sky130_fd_sc_hd__clkbuf_1
Xwire4483 net4486 VGND VGND VPWR VPWR net4483 sky130_fd_sc_hd__buf_1
Xwire3760 net3761 VGND VGND VPWR VPWR net3760 sky130_fd_sc_hd__clkbuf_1
Xwire3771 net3772 VGND VGND VPWR VPWR net3771 sky130_fd_sc_hd__clkbuf_1
X_19762_ _11594_ _11596_ VGND VGND VPWR VPWR _11597_ sky130_fd_sc_hd__nor2_1
Xwire3782 net3783 VGND VGND VPWR VPWR net3782 sky130_fd_sc_hd__clkbuf_1
X_16974_ net5989 _08919_ VGND VGND VPWR VPWR _08937_ sky130_fd_sc_hd__nor2_1
Xwire3793 net3794 VGND VGND VPWR VPWR net3793 sky130_fd_sc_hd__clkbuf_1
X_18713_ _10554_ _10557_ VGND VGND VPWR VPWR _10559_ sky130_fd_sc_hd__nor2_1
X_15925_ net1527 net1262 VGND VGND VPWR VPWR _07994_ sky130_fd_sc_hd__xnor2_1
X_19693_ net1058 _11528_ VGND VGND VPWR VPWR _11529_ sky130_fd_sc_hd__nor2_1
Xinput8 angle_in[1] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_1
XFILLER_0_190_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15856_ net827 _07888_ _07862_ VGND VGND VPWR VPWR _07925_ sky130_fd_sc_hd__o21ba_1
X_18644_ net3223 _10487_ _10489_ net6817 _10490_ VGND VGND VPWR VPWR _10491_ sky130_fd_sc_hd__o221a_1
X_14807_ net9008 net3004 _06920_ VGND VGND VPWR VPWR _00175_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18575_ net6972 _10421_ _10422_ VGND VGND VPWR VPWR _10423_ sky130_fd_sc_hd__o21ai_1
X_15787_ net1264 _07856_ VGND VGND VPWR VPWR _07857_ sky130_fd_sc_hd__nor2_1
X_12999_ _05156_ _05157_ VGND VGND VPWR VPWR _05272_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17526_ net6742 _09405_ _09409_ VGND VGND VPWR VPWR _09410_ sky130_fd_sc_hd__o21a_1
XFILLER_0_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14738_ net9104 net2861 net2865 _06872_ VGND VGND VPWR VPWR _00154_ sky130_fd_sc_hd__a22o_1
XFILLER_0_188_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17457_ svm0.counter\[3\] net2577 VGND VGND VPWR VPWR _09352_ sky130_fd_sc_hd__nor2_1
XFILLER_0_184_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14669_ net7455 net7163 VGND VGND VPWR VPWR _06821_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16408_ net2654 net2218 net1840 _08469_ VGND VGND VPWR VPWR _08470_ sky130_fd_sc_hd__o31a_1
XFILLER_0_7_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17388_ svm0.delta\[5\] _09292_ VGND VGND VPWR VPWR _09296_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19127_ net3187 _10963_ VGND VGND VPWR VPWR _10964_ sky130_fd_sc_hd__xor2_1
X_16339_ net1248 _08401_ VGND VGND VPWR VPWR _08402_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19058_ net6360 _10811_ _10894_ net6293 _10830_ VGND VGND VPWR VPWR _10895_ sky130_fd_sc_hd__o221a_1
Xfanout6291 net6304 VGND VGND VPWR VPWR net6291 sky130_fd_sc_hd__buf_1
XFILLER_0_125_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18009_ net7052 _09859_ VGND VGND VPWR VPWR _09860_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_2_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21020_ _01032_ _01035_ VGND VGND VPWR VPWR _01036_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1109 net1110 VGND VGND VPWR VPWR net1109 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_184_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22971_ _02853_ VGND VGND VPWR VPWR _00652_ sky130_fd_sc_hd__clkbuf_1
X_24710_ _04536_ _04544_ _04545_ VGND VGND VPWR VPWR _04546_ sky130_fd_sc_hd__a21o_1
X_21922_ net5540 net5669 VGND VGND VPWR VPWR _01930_ sky130_fd_sc_hd__nand2_1
X_25690_ clknet_leaf_6_clk _00563_ net8562 VGND VGND VPWR VPWR pid_d.curr_error\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_24641_ _04492_ _04495_ VGND VGND VPWR VPWR _04496_ sky130_fd_sc_hd__xnor2_1
X_21853_ _01770_ _01773_ _01861_ VGND VGND VPWR VPWR _01862_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_167_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20804_ net5936 net5425 VGND VGND VPWR VPWR _00820_ sky130_fd_sc_hd__nand2_2
X_24572_ _04424_ _04427_ VGND VGND VPWR VPWR _04428_ sky130_fd_sc_hd__xnor2_2
X_21784_ net1048 _01793_ VGND VGND VPWR VPWR _01794_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_38_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length5126 net5117 VGND VGND VPWR VPWR net5126 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23523_ pid_q.curr_int\[1\] pid_q.prev_int\[1\] _03390_ VGND VGND VPWR VPWR _03391_
+ sky130_fd_sc_hd__o21a_1
X_20735_ net5544 net5810 VGND VGND VPWR VPWR _12506_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8738 net8739 VGND VGND VPWR VPWR net8738 sky130_fd_sc_hd__buf_1
X_23454_ net4575 net5054 VGND VGND VPWR VPWR _03323_ sky130_fd_sc_hd__nand2_1
Xwire406 net407 VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__clkbuf_1
Xmax_length4447 pid_q.out\[6\] VGND VGND VPWR VPWR net4447 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20666_ net6755 net3305 _09143_ _12264_ _12442_ VGND VGND VPWR VPWR _12443_ sky130_fd_sc_hd__o221a_1
Xwire417 net418 VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__clkbuf_1
Xwire428 net429 VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__clkbuf_1
X_22405_ _04872_ _02406_ VGND VGND VPWR VPWR _02407_ sky130_fd_sc_hd__nor2_1
Xwire439 _07740_ VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__clkbuf_1
X_23385_ _03193_ _03190_ _03194_ VGND VGND VPWR VPWR _03255_ sky130_fd_sc_hd__a21o_1
X_20597_ net6196 net1396 VGND VGND VPWR VPWR _12379_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_144_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length3768 net3769 VGND VGND VPWR VPWR net3768 sky130_fd_sc_hd__buf_1
XFILLER_0_190_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3779 _01873_ VGND VGND VPWR VPWR net3779 sky130_fd_sc_hd__buf_1
X_25124_ net4391 _04849_ net2391 net5975 VGND VGND VPWR VPWR _00805_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22336_ _02320_ _02318_ _02338_ VGND VGND VPWR VPWR _02339_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_162_Left_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25055_ net239 net1630 _04803_ net9173 _04804_ VGND VGND VPWR VPWR _00785_ sky130_fd_sc_hd__a221o_1
X_22267_ _02269_ _02185_ _02270_ VGND VGND VPWR VPWR _02271_ sky130_fd_sc_hd__o21a_1
XFILLER_0_130_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire3001 net3002 VGND VGND VPWR VPWR net3001 sky130_fd_sc_hd__clkbuf_1
X_24006_ net932 _03867_ _03868_ VGND VGND VPWR VPWR _03869_ sky130_fd_sc_hd__o21ai_2
Xwire3012 net3013 VGND VGND VPWR VPWR net3012 sky130_fd_sc_hd__clkbuf_1
X_21218_ net861 _01233_ VGND VGND VPWR VPWR _01234_ sky130_fd_sc_hd__xnor2_1
Xwire3023 net3024 VGND VGND VPWR VPWR net3023 sky130_fd_sc_hd__clkbuf_1
X_22198_ net1036 _02202_ net1168 VGND VGND VPWR VPWR _02203_ sky130_fd_sc_hd__a21bo_1
Xwire3034 net3035 VGND VGND VPWR VPWR net3034 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2300 net2301 VGND VGND VPWR VPWR net2300 sky130_fd_sc_hd__clkbuf_1
Xwire3045 net3046 VGND VGND VPWR VPWR net3045 sky130_fd_sc_hd__buf_1
Xwire3056 net3057 VGND VGND VPWR VPWR net3056 sky130_fd_sc_hd__clkbuf_1
Xwire2311 net2312 VGND VGND VPWR VPWR net2311 sky130_fd_sc_hd__buf_1
Xwire2322 net2323 VGND VGND VPWR VPWR net2322 sky130_fd_sc_hd__buf_1
XFILLER_0_40_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3067 _02722_ VGND VGND VPWR VPWR net3067 sky130_fd_sc_hd__clkbuf_1
Xwire2333 net2334 VGND VGND VPWR VPWR net2333 sky130_fd_sc_hd__clkbuf_1
X_21149_ _01157_ _01164_ VGND VGND VPWR VPWR _01165_ sky130_fd_sc_hd__xnor2_1
Xwire3078 _02604_ VGND VGND VPWR VPWR net3078 sky130_fd_sc_hd__buf_1
Xwire2344 net2345 VGND VGND VPWR VPWR net2344 sky130_fd_sc_hd__buf_1
Xwire3089 _02553_ VGND VGND VPWR VPWR net3089 sky130_fd_sc_hd__buf_1
Xwire2355 _04912_ VGND VGND VPWR VPWR net2355 sky130_fd_sc_hd__clkbuf_1
Xwire1621 net1626 VGND VGND VPWR VPWR net1621 sky130_fd_sc_hd__buf_1
Xwire2366 net2367 VGND VGND VPWR VPWR net2366 sky130_fd_sc_hd__clkbuf_1
X_13971_ net1961 net1583 VGND VGND VPWR VPWR _06236_ sky130_fd_sc_hd__nor2_1
Xwire2377 net2378 VGND VGND VPWR VPWR net2377 sky130_fd_sc_hd__clkbuf_1
Xwire1632 _04752_ VGND VGND VPWR VPWR net1632 sky130_fd_sc_hd__buf_1
Xwire1643 _04529_ VGND VGND VPWR VPWR net1643 sky130_fd_sc_hd__buf_1
Xwire2388 net2389 VGND VGND VPWR VPWR net2388 sky130_fd_sc_hd__buf_1
Xwire2399 net2400 VGND VGND VPWR VPWR net2399 sky130_fd_sc_hd__clkbuf_2
Xwire1654 _04141_ VGND VGND VPWR VPWR net1654 sky130_fd_sc_hd__buf_1
X_15710_ net2647 net3465 VGND VGND VPWR VPWR _07781_ sky130_fd_sc_hd__nor2_1
X_24908_ net122 net125 net124 net8886 VGND VGND VPWR VPWR _04698_ sky130_fd_sc_hd__or4_1
X_12922_ net1957 _05111_ VGND VGND VPWR VPWR _05195_ sky130_fd_sc_hd__nor2_1
Xwire1676 _03004_ VGND VGND VPWR VPWR net1676 sky130_fd_sc_hd__dlymetal6s2s_1
X_16690_ matmul0.alpha_pass\[10\] net528 net6550 VGND VGND VPWR VPWR _08721_ sky130_fd_sc_hd__mux2_1
X_25888_ clknet_leaf_17_clk _00761_ net8628 VGND VGND VPWR VPWR pid_q.kp\[0\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_171_Left_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1687 _02695_ VGND VGND VPWR VPWR net1687 sky130_fd_sc_hd__buf_1
Xwire1698 _02568_ VGND VGND VPWR VPWR net1698 sky130_fd_sc_hd__buf_1
XFILLER_0_77_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15641_ matmul0.matmul_stage_inst.e\[15\] _07151_ _07152_ net7378 VGND VGND VPWR
+ VPWR _07713_ sky130_fd_sc_hd__a22o_1
X_24839_ net4933 net2008 net2001 net586 VGND VGND VPWR VPWR _00721_ sky130_fd_sc_hd__a22o_1
X_12853_ _05047_ _05124_ _05125_ VGND VGND VPWR VPWR _05126_ sky130_fd_sc_hd__a21oi_2
X_18360_ net6842 net6789 VGND VGND VPWR VPWR _10211_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15572_ _07631_ _07633_ VGND VGND VPWR VPWR _07644_ sky130_fd_sc_hd__or2b_1
X_12784_ net1958 VGND VGND VPWR VPWR _05057_ sky130_fd_sc_hd__buf_1
XFILLER_0_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17311_ net4024 _09224_ VGND VGND VPWR VPWR _09225_ sky130_fd_sc_hd__nand2_1
Xmax_length6350 net6344 VGND VGND VPWR VPWR net6350 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_56_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14523_ net7282 net5253 VGND VGND VPWR VPWR _06703_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18291_ net963 _09834_ _10141_ VGND VGND VPWR VPWR _10142_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_138_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17242_ _09188_ VGND VGND VPWR VPWR _09189_ sky130_fd_sc_hd__buf_1
Xmax_length5671 net5672 VGND VGND VPWR VPWR net5671 sky130_fd_sc_hd__dlymetal6s2s_1
X_14454_ _06644_ matmul0.b_in\[15\] net995 VGND VGND VPWR VPWR _06645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length4970 net4971 VGND VGND VPWR VPWR net4970 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13405_ _05668_ net581 _05674_ VGND VGND VPWR VPWR _05678_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17173_ _09122_ _09124_ VGND VGND VPWR VPWR _09125_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4981 net4982 VGND VGND VPWR VPWR net4981 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_180_Left_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14385_ net7198 net1296 net2893 net5315 _06591_ VGND VGND VPWR VPWR _06592_ sky130_fd_sc_hd__a221o_1
Xwire940 _02587_ VGND VGND VPWR VPWR net940 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire951 _12122_ VGND VGND VPWR VPWR net951 sky130_fd_sc_hd__buf_1
XFILLER_0_84_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire962 _09949_ VGND VGND VPWR VPWR net962 sky130_fd_sc_hd__buf_1
X_16124_ _08188_ _08189_ VGND VGND VPWR VPWR _08190_ sky130_fd_sc_hd__xnor2_1
X_13336_ net2964 VGND VGND VPWR VPWR _05609_ sky130_fd_sc_hd__buf_1
XFILLER_0_107_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire973 net974 VGND VGND VPWR VPWR net973 sky130_fd_sc_hd__clkbuf_1
Xwire984 net985 VGND VGND VPWR VPWR net984 sky130_fd_sc_hd__buf_1
Xclkbuf_4_5__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_4_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16055_ net2747 net2656 VGND VGND VPWR VPWR _08122_ sky130_fd_sc_hd__nor2_1
X_13267_ _05412_ _05415_ VGND VGND VPWR VPWR _05540_ sky130_fd_sc_hd__xor2_1
XFILLER_0_122_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15006_ net3573 net3569 VGND VGND VPWR VPWR _07080_ sky130_fd_sc_hd__or2_1
X_13198_ net733 net682 VGND VGND VPWR VPWR _05471_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_47_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4280 net4281 VGND VGND VPWR VPWR net4280 sky130_fd_sc_hd__clkbuf_1
X_19814_ net6068 net6041 VGND VGND VPWR VPWR _11648_ sky130_fd_sc_hd__nand2_1
Xwire4291 net4292 VGND VGND VPWR VPWR net4291 sky130_fd_sc_hd__buf_1
X_19745_ _11576_ _11579_ net6176 VGND VGND VPWR VPWR _11580_ sky130_fd_sc_hd__mux2_1
X_16957_ net2177 net1825 net7138 VGND VGND VPWR VPWR _08920_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_194_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15908_ _07967_ _07976_ VGND VGND VPWR VPWR _07977_ sky130_fd_sc_hd__xnor2_1
X_19676_ net3162 _11177_ _11511_ VGND VGND VPWR VPWR _11512_ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16888_ net6368 net6390 VGND VGND VPWR VPWR _08852_ sky130_fd_sc_hd__or2b_1
XFILLER_0_154_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18627_ _10472_ _10473_ VGND VGND VPWR VPWR _10474_ sky130_fd_sc_hd__nand2_1
X_15839_ _07890_ _07908_ VGND VGND VPWR VPWR _07909_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18558_ net765 _10404_ _10405_ VGND VGND VPWR VPWR _10406_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17509_ svm0.delta\[11\] _09395_ VGND VGND VPWR VPWR _09396_ sky130_fd_sc_hd__xnor2_1
X_18489_ net765 VGND VGND VPWR VPWR _10339_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20520_ net6324 net1470 VGND VGND VPWR VPWR _12307_ sky130_fd_sc_hd__nand2_1
Xmax_length3009 _00008_ VGND VGND VPWR VPWR net3009 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_170_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20451_ _12236_ _12235_ _12240_ _12243_ VGND VGND VPWR VPWR _12244_ sky130_fd_sc_hd__o31a_1
XFILLER_0_132_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23170_ net5116 net4719 _03039_ VGND VGND VPWR VPWR _03040_ sky130_fd_sc_hd__a21o_1
XFILLER_0_113_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20382_ cordic0.slte0.opA\[7\] VGND VGND VPWR VPWR _12181_ sky130_fd_sc_hd__inv_2
Xmax_length1618 _04901_ VGND VGND VPWR VPWR net1618 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22121_ _02025_ _02027_ _02026_ VGND VGND VPWR VPWR _02127_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22052_ net2067 _02058_ VGND VGND VPWR VPWR _02059_ sky130_fd_sc_hd__xnor2_2
X_21003_ _00889_ _00892_ VGND VGND VPWR VPWR _01019_ sky130_fd_sc_hd__xor2_1
X_25811_ clknet_leaf_36_clk _00684_ net8797 VGND VGND VPWR VPWR pid_q.prev_error\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_25742_ clknet_leaf_8_clk _00615_ net8554 VGND VGND VPWR VPWR pid_d.kp\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22954_ _02835_ _02837_ _02841_ _02513_ VGND VGND VPWR VPWR _02842_ sky130_fd_sc_hd__a31o_1
X_21905_ net4352 _01912_ _01913_ VGND VGND VPWR VPWR _01914_ sky130_fd_sc_hd__and3_1
X_25673_ clknet_leaf_4_clk _00546_ net8563 VGND VGND VPWR VPWR pid_d.prev_error\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_22885_ net5977 _02779_ VGND VGND VPWR VPWR _02780_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_195_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24624_ net4823 net4498 _04426_ _04478_ net4490 VGND VGND VPWR VPWR _04479_ sky130_fd_sc_hd__o32a_1
X_21836_ _01755_ _01760_ _01844_ VGND VGND VPWR VPWR _01845_ sky130_fd_sc_hd__o21a_1
XFILLER_0_194_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout8429 net8434 VGND VGND VPWR VPWR net8429 sky130_fd_sc_hd__clkbuf_2
X_24555_ _04355_ _04364_ _04339_ VGND VGND VPWR VPWR _04411_ sky130_fd_sc_hd__o21a_1
X_21767_ _01748_ _01776_ VGND VGND VPWR VPWR _01777_ sky130_fd_sc_hd__xnor2_1
Xwire8502 net8503 VGND VGND VPWR VPWR net8502 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout7717 net7729 VGND VGND VPWR VPWR net7717 sky130_fd_sc_hd__clkbuf_1
Xwire8513 net8514 VGND VGND VPWR VPWR net8513 sky130_fd_sc_hd__clkbuf_1
Xwire8524 net8529 VGND VGND VPWR VPWR net8524 sky130_fd_sc_hd__clkbuf_1
X_23506_ _03371_ _03374_ VGND VGND VPWR VPWR _03375_ sky130_fd_sc_hd__xor2_1
XFILLER_0_19_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8535 net8536 VGND VGND VPWR VPWR net8535 sky130_fd_sc_hd__clkbuf_1
X_20718_ net966 _12489_ VGND VGND VPWR VPWR _12490_ sky130_fd_sc_hd__nand2_1
Xwire8546 net8547 VGND VGND VPWR VPWR net8546 sky130_fd_sc_hd__clkbuf_1
X_24486_ net4523 net4825 VGND VGND VPWR VPWR _04343_ sky130_fd_sc_hd__nand2_2
X_21698_ net5396 VGND VGND VPWR VPWR _01709_ sky130_fd_sc_hd__inv_2
Xwire203 _02842_ VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_1
Xwire8557 net8558 VGND VGND VPWR VPWR net8557 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7823 net7824 VGND VGND VPWR VPWR net7823 sky130_fd_sc_hd__buf_1
Xwire8568 net8564 VGND VGND VPWR VPWR net8568 sky130_fd_sc_hd__buf_1
Xwire214 net215 VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_1
Xwire225 net226 VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__clkbuf_1
Xwire7834 net7827 VGND VGND VPWR VPWR net7834 sky130_fd_sc_hd__buf_1
Xwire8579 net8580 VGND VGND VPWR VPWR net8579 sky130_fd_sc_hd__buf_1
XFILLER_0_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length3521 _07066_ VGND VGND VPWR VPWR net3521 sky130_fd_sc_hd__buf_1
XFILLER_0_92_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23437_ _03306_ VGND VGND VPWR VPWR _03307_ sky130_fd_sc_hd__inv_2
Xwire7845 net7846 VGND VGND VPWR VPWR net7845 sky130_fd_sc_hd__clkbuf_1
Xwire236 net237 VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__buf_1
XFILLER_0_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20649_ net6757 net3327 net2168 _12315_ VGND VGND VPWR VPWR _12427_ sky130_fd_sc_hd__a22o_1
Xwire247 net248 VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__clkbuf_1
Xwire7867 net7868 VGND VGND VPWR VPWR net7867 sky130_fd_sc_hd__clkbuf_1
Xwire258 _04656_ VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__clkbuf_1
Xmax_length2820 _07092_ VGND VGND VPWR VPWR net2820 sky130_fd_sc_hd__buf_1
Xwire269 net270 VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__buf_1
X_14170_ _06421_ _06430_ VGND VGND VPWR VPWR _06431_ sky130_fd_sc_hd__xor2_1
Xwire7889 net7899 VGND VGND VPWR VPWR net7889 sky130_fd_sc_hd__buf_1
X_23368_ net697 net755 _03236_ _03237_ VGND VGND VPWR VPWR _03238_ sky130_fd_sc_hd__a211o_1
XFILLER_0_104_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13121_ _05390_ _05393_ VGND VGND VPWR VPWR _05394_ sky130_fd_sc_hd__xor2_1
X_25107_ net4297 net9248 net4308 VGND VGND VPWR VPWR _04849_ sky130_fd_sc_hd__a21oi_2
Xmax_length2875 _06805_ VGND VGND VPWR VPWR net2875 sky130_fd_sc_hd__buf_1
X_22319_ _02318_ _02322_ VGND VGND VPWR VPWR _02323_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2886 net2887 VGND VGND VPWR VPWR net2886 sky130_fd_sc_hd__clkbuf_2
X_23299_ _03149_ _03167_ _03168_ VGND VGND VPWR VPWR _03169_ sky130_fd_sc_hd__o21ai_1
Xmax_length2897 net2899 VGND VGND VPWR VPWR net2897 sky130_fd_sc_hd__clkbuf_1
X_25038_ net3739 net1157 _04789_ VGND VGND VPWR VPWR _04790_ sky130_fd_sc_hd__a21o_1
X_13052_ _05030_ _05321_ _05324_ VGND VGND VPWR VPWR _05325_ sky130_fd_sc_hd__o21ai_1
X_17860_ net7091 net7027 VGND VGND VPWR VPWR _09711_ sky130_fd_sc_hd__nand2_1
Xwire2130 _10363_ VGND VGND VPWR VPWR net2130 sky130_fd_sc_hd__buf_1
Xwire2141 _09719_ VGND VGND VPWR VPWR net2141 sky130_fd_sc_hd__buf_1
Xwire2152 _09503_ VGND VGND VPWR VPWR net2152 sky130_fd_sc_hd__clkbuf_1
X_16811_ cordic0.cos\[8\] matmul0.cos\[8\] net3367 VGND VGND VPWR VPWR _08796_ sky130_fd_sc_hd__mux2_1
Xwire2163 _09189_ VGND VGND VPWR VPWR net2163 sky130_fd_sc_hd__dlymetal6s2s_1
X_17791_ net7133 net7120 VGND VGND VPWR VPWR _09642_ sky130_fd_sc_hd__nand2b_1
Xclkbuf_4_13__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_4_13__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xwire2174 net2175 VGND VGND VPWR VPWR net2174 sky130_fd_sc_hd__buf_1
Xwire2185 net2186 VGND VGND VPWR VPWR net2185 sky130_fd_sc_hd__clkbuf_1
Xwire1440 _10306_ VGND VGND VPWR VPWR net1440 sky130_fd_sc_hd__buf_1
X_19530_ _11303_ _11364_ _11365_ _11366_ VGND VGND VPWR VPWR _11367_ sky130_fd_sc_hd__o22a_1
Xwire2196 net2197 VGND VGND VPWR VPWR net2196 sky130_fd_sc_hd__buf_1
Xwire1462 net1463 VGND VGND VPWR VPWR net1462 sky130_fd_sc_hd__clkbuf_1
X_13954_ net7664 net1125 VGND VGND VPWR VPWR _06219_ sky130_fd_sc_hd__nand2_1
X_16742_ net7567 matmul0.b\[7\] net3381 VGND VGND VPWR VPWR _08760_ sky130_fd_sc_hd__mux2_1
Xwire1473 net1474 VGND VGND VPWR VPWR net1473 sky130_fd_sc_hd__buf_1
Xwire1484 net1485 VGND VGND VPWR VPWR net1484 sky130_fd_sc_hd__clkbuf_2
X_12905_ net7779 _04905_ _04907_ VGND VGND VPWR VPWR _05178_ sky130_fd_sc_hd__and3_1
Xwire1495 net1496 VGND VGND VPWR VPWR net1495 sky130_fd_sc_hd__buf_1
X_19461_ _11294_ _11297_ VGND VGND VPWR VPWR _11298_ sky130_fd_sc_hd__xnor2_1
X_16673_ _08704_ _08700_ _08705_ VGND VGND VPWR VPWR _08706_ sky130_fd_sc_hd__o21a_1
X_13885_ _06142_ _06151_ VGND VGND VPWR VPWR _06152_ sky130_fd_sc_hd__xnor2_1
X_18412_ net9059 net2289 _09598_ _10262_ VGND VGND VPWR VPWR _00439_ sky130_fd_sc_hd__a31o_1
XFILLER_0_97_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12836_ _05034_ _05036_ VGND VGND VPWR VPWR _05109_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15624_ _07606_ _07693_ _07695_ VGND VGND VPWR VPWR _07696_ sky130_fd_sc_hd__a21o_1
X_19392_ _11222_ _11224_ _11226_ _11228_ VGND VGND VPWR VPWR _11229_ sky130_fd_sc_hd__a211o_1
XFILLER_0_33_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15555_ net1273 _07496_ _07500_ VGND VGND VPWR VPWR _07628_ sky130_fd_sc_hd__o21ba_1
X_18343_ _10132_ _10135_ VGND VGND VPWR VPWR _10194_ sky130_fd_sc_hd__or2b_1
X_12767_ net7758 net2345 net2342 VGND VGND VPWR VPWR _05040_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6180 net6177 VGND VGND VPWR VPWR net6180 sky130_fd_sc_hd__clkbuf_1
X_14506_ _06686_ _06687_ VGND VGND VPWR VPWR _06688_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18274_ _10121_ net3228 VGND VGND VPWR VPWR _10125_ sky130_fd_sc_hd__xnor2_1
X_15486_ net3478 VGND VGND VPWR VPWR _07560_ sky130_fd_sc_hd__buf_1
XFILLER_0_154_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12698_ _04955_ _04970_ VGND VGND VPWR VPWR _04971_ sky130_fd_sc_hd__xnor2_1
X_14437_ matmul0.beta_pass\[11\] net1294 net2890 net4413 _06631_ VGND VGND VPWR VPWR
+ _06632_ sky130_fd_sc_hd__a221o_1
X_17225_ net6806 _09163_ VGND VGND VPWR VPWR _09173_ sky130_fd_sc_hd__nand2_1
Xinput11 angle_in[4] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_1
XFILLER_0_86_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput22 currA_in[14] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput33 currB_in[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput44 currB_in[5] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17156_ net3301 net1234 _09107_ _09109_ VGND VGND VPWR VPWR _00335_ sky130_fd_sc_hd__a31o_1
Xinput55 currT_in[15] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_1
Xwire770 _09378_ VGND VGND VPWR VPWR net770 sky130_fd_sc_hd__buf_1
X_14368_ net8300 net3637 VGND VGND VPWR VPWR _06579_ sky130_fd_sc_hd__and2_1
Xwire781 _05978_ VGND VGND VPWR VPWR net781 sky130_fd_sc_hd__buf_1
Xinput66 periodTop[10] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput77 periodTop[6] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire792 _04309_ VGND VGND VPWR VPWR net792 sky130_fd_sc_hd__buf_2
X_16107_ net3561 net3394 VGND VGND VPWR VPWR _08173_ sky130_fd_sc_hd__nand2_1
Xinput88 pid_d_addr[1] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_1
X_13319_ net7722 net2321 net2317 VGND VGND VPWR VPWR _05592_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput99 pid_d_data[11] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_1
X_17087_ net7039 _09014_ _09041_ VGND VGND VPWR VPWR _09045_ sky130_fd_sc_hd__or3b_1
XFILLER_0_40_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14299_ net4236 net1991 _06520_ VGND VGND VPWR VPWR _06521_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16038_ _08098_ _08104_ VGND VGND VPWR VPWR _08105_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17989_ _09830_ _09833_ _09838_ net963 VGND VGND VPWR VPWR _09840_ sky130_fd_sc_hd__a31oi_1
X_19728_ _11431_ _11501_ VGND VGND VPWR VPWR _11563_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19659_ net6012 net2504 VGND VGND VPWR VPWR _11495_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_181_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22670_ _02621_ VGND VGND VPWR VPWR _00583_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21621_ _01632_ VGND VGND VPWR VPWR _01633_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_158_Right_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24340_ _04144_ _04150_ _04198_ VGND VGND VPWR VPWR _04199_ sky130_fd_sc_hd__a21oi_1
X_21552_ net5729 net5549 VGND VGND VPWR VPWR _01564_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20503_ net3169 net2088 net6350 VGND VGND VPWR VPWR _12290_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24271_ net4917 net4502 VGND VGND VPWR VPWR _04131_ sky130_fd_sc_hd__nand2_2
Xwire6407 net6408 VGND VGND VPWR VPWR net6407 sky130_fd_sc_hd__buf_1
X_21483_ _01366_ _01368_ _01364_ VGND VGND VPWR VPWR _01496_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_133_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6418 cordic0.slte0.opB\[4\] VGND VGND VPWR VPWR net6418 sky130_fd_sc_hd__buf_1
XFILLER_0_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6429 cordic0.sin\[3\] VGND VGND VPWR VPWR net6429 sky130_fd_sc_hd__clkbuf_1
X_23222_ _02993_ _03091_ VGND VGND VPWR VPWR _03092_ sky130_fd_sc_hd__xnor2_2
X_20434_ _12226_ _12228_ VGND VGND VPWR VPWR _12229_ sky130_fd_sc_hd__xor2_1
Xwire5717 net5712 VGND VGND VPWR VPWR net5717 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5728 net5729 VGND VGND VPWR VPWR net5728 sky130_fd_sc_hd__clkbuf_1
X_23153_ _03021_ _03022_ VGND VGND VPWR VPWR _03023_ sky130_fd_sc_hd__xnor2_1
X_20365_ _12159_ net1054 _12156_ VGND VGND VPWR VPWR _12165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22104_ _02108_ _02019_ _02109_ VGND VGND VPWR VPWR _02110_ sky130_fd_sc_hd__o21a_1
X_23084_ _02871_ _02873_ VGND VGND VPWR VPWR _02954_ sky130_fd_sc_hd__nand2_1
X_20296_ _12089_ _12100_ VGND VGND VPWR VPWR _12102_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22035_ _02040_ _02041_ VGND VGND VPWR VPWR _02042_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23986_ _03848_ _03849_ VGND VGND VPWR VPWR _03850_ sky130_fd_sc_hd__nor2_1
X_25725_ clknet_leaf_13_clk _00598_ net8609 VGND VGND VPWR VPWR pid_d.mult0.a\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_22937_ _02826_ VGND VGND VPWR VPWR _00645_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13670_ net7700 net2308 net1953 VGND VGND VPWR VPWR _05939_ sky130_fd_sc_hd__and3_2
X_25656_ clknet_leaf_2_clk _00529_ net8573 VGND VGND VPWR VPWR pid_d.curr_int\[10\]
+ sky130_fd_sc_hd__dfrtp_4
X_22868_ _02762_ _02763_ VGND VGND VPWR VPWR _02765_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24607_ _04423_ _04461_ VGND VGND VPWR VPWR _04462_ sky130_fd_sc_hd__nand2_1
X_12621_ _04893_ VGND VGND VPWR VPWR _04894_ sky130_fd_sc_hd__clkbuf_2
X_21819_ _01748_ _01775_ _01762_ VGND VGND VPWR VPWR _01828_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_167_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25587_ clknet_leaf_99_clk _00460_ net8382 VGND VGND VPWR VPWR cordic0.cos\[7\] sky130_fd_sc_hd__dfrtp_1
X_22799_ _02707_ VGND VGND VPWR VPWR _00626_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_125_Right_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8310 net8311 VGND VGND VPWR VPWR net8310 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15340_ _07310_ _07312_ VGND VGND VPWR VPWR _07414_ sky130_fd_sc_hd__xnor2_1
Xwire8321 net8322 VGND VGND VPWR VPWR net8321 sky130_fd_sc_hd__clkbuf_1
X_24538_ _04315_ _04373_ _04393_ net792 VGND VGND VPWR VPWR _04394_ sky130_fd_sc_hd__a22o_1
Xfanout7525 net7528 VGND VGND VPWR VPWR net7525 sky130_fd_sc_hd__clkbuf_1
Xwire8332 net8328 VGND VGND VPWR VPWR net8332 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_80_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length4041 _09032_ VGND VGND VPWR VPWR net4041 sky130_fd_sc_hd__buf_1
Xwire8354 net8356 VGND VGND VPWR VPWR net8354 sky130_fd_sc_hd__buf_1
Xwire7620 net7621 VGND VGND VPWR VPWR net7620 sky130_fd_sc_hd__clkbuf_1
Xmax_length4052 _08943_ VGND VGND VPWR VPWR net4052 sky130_fd_sc_hd__clkbuf_1
Xwire8365 net8366 VGND VGND VPWR VPWR net8365 sky130_fd_sc_hd__buf_1
Xwire7631 net7632 VGND VGND VPWR VPWR net7631 sky130_fd_sc_hd__buf_1
XFILLER_0_108_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15271_ net2838 net3466 VGND VGND VPWR VPWR _07345_ sky130_fd_sc_hd__nor2_1
X_24469_ net4001 _04326_ VGND VGND VPWR VPWR _04327_ sky130_fd_sc_hd__nor2_1
Xwire8376 net8377 VGND VGND VPWR VPWR net8376 sky130_fd_sc_hd__buf_1
XFILLER_0_53_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7642 net7641 VGND VGND VPWR VPWR net7642 sky130_fd_sc_hd__buf_1
Xwire8387 net8385 VGND VGND VPWR VPWR net8387 sky130_fd_sc_hd__buf_1
XFILLER_0_108_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17010_ net4060 VGND VGND VPWR VPWR _08971_ sky130_fd_sc_hd__clkbuf_2
Xmax_length3340 _08967_ VGND VGND VPWR VPWR net3340 sky130_fd_sc_hd__buf_1
X_14222_ _06434_ _06436_ _06437_ _06460_ _06459_ VGND VGND VPWR VPWR _06480_ sky130_fd_sc_hd__a41o_1
Xwire7664 net7660 VGND VGND VPWR VPWR net7664 sky130_fd_sc_hd__buf_1
XFILLER_0_11_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7675 net7676 VGND VGND VPWR VPWR net7675 sky130_fd_sc_hd__buf_1
Xwire7686 net7687 VGND VGND VPWR VPWR net7686 sky130_fd_sc_hd__clkbuf_1
Xwire6941 net6944 VGND VGND VPWR VPWR net6941 sky130_fd_sc_hd__buf_1
Xfanout6879 net6883 VGND VGND VPWR VPWR net6879 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7697 net7698 VGND VGND VPWR VPWR net7697 sky130_fd_sc_hd__buf_1
Xwire6963 net6964 VGND VGND VPWR VPWR net6963 sky130_fd_sc_hd__buf_1
Xmax_length3395 _07688_ VGND VGND VPWR VPWR net3395 sky130_fd_sc_hd__buf_1
X_14153_ net7666 _06405_ _06412_ _06413_ VGND VGND VPWR VPWR _06414_ sky130_fd_sc_hd__a31o_1
Xwire6974 net6978 VGND VGND VPWR VPWR net6974 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_100_clk clknet_4_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_100_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_46_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6996 net6993 VGND VGND VPWR VPWR net6996 sky130_fd_sc_hd__clkbuf_4
X_13104_ _05373_ _05376_ VGND VGND VPWR VPWR _05377_ sky130_fd_sc_hd__xnor2_1
X_14084_ _06298_ _06303_ _06295_ VGND VGND VPWR VPWR _06347_ sky130_fd_sc_hd__a21bo_1
X_18961_ net6189 net6142 VGND VGND VPWR VPWR _10798_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13035_ _05247_ net735 _05307_ VGND VGND VPWR VPWR _05308_ sky130_fd_sc_hd__o21ai_1
X_17912_ net2562 _09652_ net3260 VGND VGND VPWR VPWR _09763_ sky130_fd_sc_hd__a21o_1
X_18892_ _10705_ net1194 VGND VGND VPWR VPWR _10733_ sky130_fd_sc_hd__or2_1
X_17843_ net7103 net7123 VGND VGND VPWR VPWR _09694_ sky130_fd_sc_hd__and2b_1
XFILLER_0_156_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17774_ _09622_ _09623_ net3265 net3994 net7092 VGND VGND VPWR VPWR _09625_ sky130_fd_sc_hd__a32o_1
X_14986_ net3544 _07059_ VGND VGND VPWR VPWR _07060_ sky130_fd_sc_hd__xnor2_2
Xwire1270 net1271 VGND VGND VPWR VPWR net1270 sky130_fd_sc_hd__clkbuf_2
X_19513_ _11347_ net3155 VGND VGND VPWR VPWR _11350_ sky130_fd_sc_hd__xnor2_1
Xwire1281 net1282 VGND VGND VPWR VPWR net1281 sky130_fd_sc_hd__clkbuf_1
Xwire1292 _06655_ VGND VGND VPWR VPWR net1292 sky130_fd_sc_hd__clkbuf_2
X_16725_ matmul0.alpha_pass\[15\] _08750_ net6557 VGND VGND VPWR VPWR _08751_ sky130_fd_sc_hd__mux2_1
X_13937_ _06198_ _06202_ VGND VGND VPWR VPWR _06203_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_53_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19444_ _11278_ _11279_ net2507 VGND VGND VPWR VPWR _11281_ sky130_fd_sc_hd__a21oi_2
X_13868_ _06128_ _06134_ VGND VGND VPWR VPWR _06135_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16656_ _08691_ VGND VGND VPWR VPWR _00253_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12819_ _05090_ _05091_ VGND VGND VPWR VPWR _05092_ sky130_fd_sc_hd__xnor2_1
X_15607_ net1851 net1537 VGND VGND VPWR VPWR _07679_ sky130_fd_sc_hd__xnor2_1
X_19375_ net3166 net2523 VGND VGND VPWR VPWR _11212_ sky130_fd_sc_hd__or2_1
X_13799_ net782 _06065_ _06066_ VGND VGND VPWR VPWR _06067_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_146_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16587_ matmul0.matmul_stage_inst.mult2\[4\] net396 net2617 VGND VGND VPWR VPWR _08641_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18326_ net6945 _09680_ _10176_ net3986 _09796_ VGND VGND VPWR VPWR _10177_ sky130_fd_sc_hd__a221o_1
XFILLER_0_84_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8760 net8766 VGND VGND VPWR VPWR net8760 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15538_ _07513_ _07521_ _07510_ VGND VGND VPWR VPWR _07611_ sky130_fd_sc_hd__a21o_1
XFILLER_0_173_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15469_ _07502_ _07542_ VGND VGND VPWR VPWR _07543_ sky130_fd_sc_hd__xnor2_2
X_18257_ net7012 net7115 VGND VGND VPWR VPWR _10108_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_114_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17208_ net3285 VGND VGND VPWR VPWR _09158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18188_ net6847 net6875 VGND VGND VPWR VPWR _10039_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_8_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17139_ _09092_ VGND VGND VPWR VPWR _09093_ sky130_fd_sc_hd__clkbuf_1
X_20150_ net6079 _11491_ _11971_ _11976_ VGND VGND VPWR VPWR _11977_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_122_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20081_ _11878_ _11909_ VGND VGND VPWR VPWR _11910_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23840_ net4490 VGND VGND VPWR VPWR _03705_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23771_ _03629_ _03636_ VGND VGND VPWR VPWR _03637_ sky130_fd_sc_hd__xnor2_2
X_20983_ _00980_ _00981_ VGND VGND VPWR VPWR _00999_ sky130_fd_sc_hd__nor2_1
X_25510_ clknet_leaf_36_clk _00390_ net8758 VGND VGND VPWR VPWR svm0.delta\[15\] sky130_fd_sc_hd__dfrtp_1
X_22722_ net8101 net92 net8099 net94 VGND VGND VPWR VPWR _02658_ sky130_fd_sc_hd__or4_1
XFILLER_0_67_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25441_ clknet_leaf_113_clk _00324_ net8340 VGND VGND VPWR VPWR cordic0.vec\[1\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_22653_ net9171 net3086 _02611_ net522 net8894 VGND VGND VPWR VPWR _00576_ sky130_fd_sc_hd__o221a_1
XFILLER_0_76_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21604_ _01603_ _01615_ VGND VGND VPWR VPWR _01616_ sky130_fd_sc_hd__xor2_1
XFILLER_0_146_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25372_ clknet_leaf_81_clk _00255_ net8709 VGND VGND VPWR VPWR matmul0.alpha_pass\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_22584_ _02563_ VGND VGND VPWR VPWR _00555_ sky130_fd_sc_hd__clkbuf_1
Xfanout6109 net6123 VGND VGND VPWR VPWR net6109 sky130_fd_sc_hd__buf_1
XFILLER_0_91_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24323_ _04180_ _04181_ VGND VGND VPWR VPWR _04183_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21535_ net702 _01546_ VGND VGND VPWR VPWR _01547_ sky130_fd_sc_hd__xor2_1
XFILLER_0_16_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6226 net6227 VGND VGND VPWR VPWR net6226 sky130_fd_sc_hd__dlymetal6s2s_1
X_24254_ net7505 _04113_ _04114_ VGND VGND VPWR VPWR _04115_ sky130_fd_sc_hd__and3_1
X_21466_ _01477_ _01478_ VGND VGND VPWR VPWR _01479_ sky130_fd_sc_hd__and2b_1
Xwire5503 net5504 VGND VGND VPWR VPWR net5503 sky130_fd_sc_hd__clkbuf_1
Xwire6248 net6249 VGND VGND VPWR VPWR net6248 sky130_fd_sc_hd__buf_1
Xwire5514 net5515 VGND VGND VPWR VPWR net5514 sky130_fd_sc_hd__buf_1
Xwire6259 net6258 VGND VGND VPWR VPWR net6259 sky130_fd_sc_hd__buf_1
X_23205_ net5158 net4742 _03073_ _03074_ net3752 VGND VGND VPWR VPWR _03075_ sky130_fd_sc_hd__a32o_1
Xwire5525 net5526 VGND VGND VPWR VPWR net5525 sky130_fd_sc_hd__buf_1
Xwire5536 net5537 VGND VGND VPWR VPWR net5536 sky130_fd_sc_hd__clkbuf_1
X_20417_ _12212_ _12213_ _08865_ VGND VGND VPWR VPWR _12214_ sky130_fd_sc_hd__mux2_1
Xwire4802 net4803 VGND VGND VPWR VPWR net4802 sky130_fd_sc_hd__buf_1
X_24185_ net930 VGND VGND VPWR VPWR _04046_ sky130_fd_sc_hd__inv_2
Xwire5547 net5541 VGND VGND VPWR VPWR net5547 sky130_fd_sc_hd__clkbuf_1
X_21397_ _01396_ _01410_ VGND VGND VPWR VPWR _01411_ sky130_fd_sc_hd__xnor2_1
Xwire4813 net4810 VGND VGND VPWR VPWR net4813 sky130_fd_sc_hd__buf_1
Xwire4824 net4825 VGND VGND VPWR VPWR net4824 sky130_fd_sc_hd__buf_1
Xwire5569 net5574 VGND VGND VPWR VPWR net5569 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23136_ _02990_ _03002_ _03005_ VGND VGND VPWR VPWR _03006_ sky130_fd_sc_hd__a21o_1
Xwire4846 net4847 VGND VGND VPWR VPWR net4846 sky130_fd_sc_hd__buf_1
X_20348_ _12140_ _12148_ _12149_ VGND VGND VPWR VPWR _12150_ sky130_fd_sc_hd__and3_1
Xwire4857 net4858 VGND VGND VPWR VPWR net4857 sky130_fd_sc_hd__buf_1
Xwire4868 net4869 VGND VGND VPWR VPWR net4868 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23067_ _02933_ _02936_ VGND VGND VPWR VPWR _02937_ sky130_fd_sc_hd__xnor2_1
X_20279_ net3314 net6476 net2604 _12085_ net2608 VGND VGND VPWR VPWR _12086_ sky130_fd_sc_hd__o311a_1
X_22018_ net5540 net5649 VGND VGND VPWR VPWR _02025_ sky130_fd_sc_hd__nand2b_1
X_14840_ net9227 matmul0.matmul_stage_inst.e\[9\] net3612 VGND VGND VPWR VPWR _06937_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14771_ net4224 net1908 VGND VGND VPWR VPWR _06898_ sky130_fd_sc_hd__and2_1
XFILLER_0_187_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23969_ _03831_ _03832_ net4704 VGND VGND VPWR VPWR _03833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13722_ _05984_ _05990_ VGND VGND VPWR VPWR _05991_ sky130_fd_sc_hd__xnor2_1
X_16510_ net881 _08569_ VGND VGND VPWR VPWR _08570_ sky130_fd_sc_hd__xnor2_1
X_25708_ clknet_leaf_6_clk _00581_ net8564 VGND VGND VPWR VPWR pid_d.mult0.b\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_17490_ net2574 _09379_ net6660 VGND VGND VPWR VPWR _09380_ sky130_fd_sc_hd__o21a_1
Xmax_length8896 net8897 VGND VGND VPWR VPWR net8896 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13653_ net7832 net1328 _05794_ VGND VGND VPWR VPWR _05923_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16441_ net976 _08465_ VGND VGND VPWR VPWR _08502_ sky130_fd_sc_hd__xnor2_1
X_25639_ clknet_leaf_102_clk _00512_ net8364 VGND VGND VPWR VPWR cordic0.vec\[0\]\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_151_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12604_ net8872 net7490 VGND VGND VPWR VPWR _04881_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19160_ net6138 net6101 net3878 VGND VGND VPWR VPWR _10997_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16372_ _08418_ net1247 _08415_ VGND VGND VPWR VPWR _08434_ sky130_fd_sc_hd__a21o_1
X_13584_ net367 _05853_ _05854_ VGND VGND VPWR VPWR _05855_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_186_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8140 net45 VGND VGND VPWR VPWR net8140 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18111_ _09860_ net2550 _09881_ VGND VGND VPWR VPWR _09962_ sky130_fd_sc_hd__o21ai_1
X_15323_ net2229 net1866 VGND VGND VPWR VPWR _07397_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8151 net8152 VGND VGND VPWR VPWR net8151 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_170_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8162 net41 VGND VGND VPWR VPWR net8162 sky130_fd_sc_hd__clkbuf_1
X_19091_ net3209 _10917_ net6300 VGND VGND VPWR VPWR _10928_ sky130_fd_sc_hd__a21oi_1
Xwire8173 net39 VGND VGND VPWR VPWR net8173 sky130_fd_sc_hd__clkbuf_1
Xfanout6632 net6648 VGND VGND VPWR VPWR net6632 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8184 net8185 VGND VGND VPWR VPWR net8184 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7450 net7451 VGND VGND VPWR VPWR net7450 sky130_fd_sc_hd__clkbuf_1
Xwire8195 net8196 VGND VGND VPWR VPWR net8195 sky130_fd_sc_hd__clkbuf_1
X_18042_ _09891_ _09892_ VGND VGND VPWR VPWR _09893_ sky130_fd_sc_hd__xnor2_4
X_15254_ _07312_ VGND VGND VPWR VPWR _07328_ sky130_fd_sc_hd__inv_2
Xwire7461 net7458 VGND VGND VPWR VPWR net7461 sky130_fd_sc_hd__clkbuf_1
Xwire7472 net7473 VGND VGND VPWR VPWR net7472 sky130_fd_sc_hd__buf_1
Xfanout5931 net5938 VGND VGND VPWR VPWR net5931 sky130_fd_sc_hd__buf_1
XFILLER_0_151_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14205_ _06415_ _06450_ VGND VGND VPWR VPWR _06464_ sky130_fd_sc_hd__or2b_1
Xwire7494 net7495 VGND VGND VPWR VPWR net7494 sky130_fd_sc_hd__clkbuf_1
Xfanout5953 net5959 VGND VGND VPWR VPWR net5953 sky130_fd_sc_hd__buf_1
Xwire6760 net6761 VGND VGND VPWR VPWR net6760 sky130_fd_sc_hd__buf_1
X_15185_ net1278 _07258_ VGND VGND VPWR VPWR _07259_ sky130_fd_sc_hd__xnor2_2
Xwire6771 net6769 VGND VGND VPWR VPWR net6771 sky130_fd_sc_hd__buf_1
XFILLER_0_2_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6793 net6792 VGND VGND VPWR VPWR net6793 sky130_fd_sc_hd__buf_1
X_14136_ _06368_ _06397_ VGND VGND VPWR VPWR _06398_ sky130_fd_sc_hd__xnor2_1
X_19993_ _11822_ _11823_ VGND VGND VPWR VPWR _11824_ sky130_fd_sc_hd__or2_1
X_14067_ net7701 net1567 VGND VGND VPWR VPWR _06330_ sky130_fd_sc_hd__nand2_1
X_18944_ _10781_ _10782_ net2133 VGND VGND VPWR VPWR _10783_ sky130_fd_sc_hd__o21a_1
X_13018_ net4259 net7878 _05290_ VGND VGND VPWR VPWR _05291_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18875_ net6770 _10436_ VGND VGND VPWR VPWR _10717_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17826_ net3246 _09676_ VGND VGND VPWR VPWR _09677_ sky130_fd_sc_hd__xor2_1
X_17757_ net6996 net7028 VGND VGND VPWR VPWR _09608_ sky130_fd_sc_hd__or2b_1
X_14969_ net4154 net4149 VGND VGND VPWR VPWR _07043_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16708_ _08734_ net383 _08735_ VGND VGND VPWR VPWR _08736_ sky130_fd_sc_hd__a21o_1
X_17688_ net6701 _09567_ svm0.tA\[12\] VGND VGND VPWR VPWR _09568_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_76_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19427_ _11262_ _11263_ VGND VGND VPWR VPWR _11264_ sky130_fd_sc_hd__nor2_2
XFILLER_0_71_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16639_ _08675_ _08676_ VGND VGND VPWR VPWR _08677_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19358_ _11146_ _11150_ _11194_ net6362 VGND VGND VPWR VPWR _11195_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18309_ net7071 _10158_ _10159_ VGND VGND VPWR VPWR _10160_ sky130_fd_sc_hd__o21ai_1
Xfanout8590 net8815 VGND VGND VPWR VPWR net8590 sky130_fd_sc_hd__buf_1
XFILLER_0_73_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19289_ net6313 net3898 _11125_ net6261 net6293 VGND VGND VPWR VPWR _11126_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21320_ _01333_ _01334_ net4356 VGND VGND VPWR VPWR _01335_ sky130_fd_sc_hd__o21a_1
X_21251_ net5415 net5945 VGND VGND VPWR VPWR _01266_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4109 net4110 VGND VGND VPWR VPWR net4109 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20202_ _12020_ net866 VGND VGND VPWR VPWR _12027_ sky130_fd_sc_hd__xnor2_1
X_21182_ _01176_ _01179_ VGND VGND VPWR VPWR _01198_ sky130_fd_sc_hd__nand2_1
Xwire3408 _07571_ VGND VGND VPWR VPWR net3408 sky130_fd_sc_hd__clkbuf_1
Xwire3419 _07516_ VGND VGND VPWR VPWR net3419 sky130_fd_sc_hd__buf_1
XFILLER_0_99_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20133_ _11873_ _11913_ _11846_ VGND VGND VPWR VPWR _11961_ sky130_fd_sc_hd__or3b_1
XFILLER_0_1_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2707 net2708 VGND VGND VPWR VPWR net2707 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_187_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24941_ _04721_ VGND VGND VPWR VPWR _00754_ sky130_fd_sc_hd__clkbuf_1
X_20064_ net3144 _11436_ net6005 VGND VGND VPWR VPWR _11893_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24872_ _04672_ net4687 net1996 VGND VGND VPWR VPWR _04673_ sky130_fd_sc_hd__mux2_1
X_23823_ net4527 net5057 _03686_ _03687_ VGND VGND VPWR VPWR _03688_ sky130_fd_sc_hd__a31o_1
XFILLER_0_174_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6702 svm0.counter\[12\] VGND VGND VPWR VPWR net6702 sky130_fd_sc_hd__clkbuf_1
X_23754_ _03616_ _03619_ VGND VGND VPWR VPWR _03620_ sky130_fd_sc_hd__xnor2_2
Xmax_length7447 net7443 VGND VGND VPWR VPWR net7447 sky130_fd_sc_hd__clkbuf_1
X_20966_ _00980_ _00981_ VGND VGND VPWR VPWR _00982_ sky130_fd_sc_hd__xor2_1
XFILLER_0_177_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22705_ pid_d.ki\[12\] net3705 _04886_ pid_d.kp\[12\] VGND VGND VPWR VPWR _02645_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23685_ _03547_ _03551_ VGND VGND VPWR VPWR _03552_ sky130_fd_sc_hd__nor2_1
X_20897_ _00891_ _00893_ _00912_ VGND VGND VPWR VPWR _00913_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25424_ clknet_leaf_91_clk _00307_ net8427 VGND VGND VPWR VPWR matmul0.cos\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_22636_ net5941 net3082 _02602_ _01335_ net8893 VGND VGND VPWR VPWR _00568_ sky130_fd_sc_hd__o221a_1
XFILLER_0_119_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25355_ clknet_leaf_42_clk _00238_ net8771 VGND VGND VPWR VPWR svm0.delta\[0\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_152_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22567_ net9037 net2043 _02548_ _02549_ VGND VGND VPWR VPWR _00552_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24306_ _04121_ _04165_ VGND VGND VPWR VPWR _04166_ sky130_fd_sc_hd__xnor2_1
Xwire6001 net6002 VGND VGND VPWR VPWR net6001 sky130_fd_sc_hd__buf_1
XFILLER_0_91_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6012 net6013 VGND VGND VPWR VPWR net6012 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_63_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21518_ _01528_ _01526_ _01418_ VGND VGND VPWR VPWR _01531_ sky130_fd_sc_hd__mux2_1
X_25286_ clknet_leaf_89_clk _00169_ net8443 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.d\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_22498_ _02443_ _02439_ VGND VGND VPWR VPWR _02499_ sky130_fd_sc_hd__nand2_1
Xwire6034 net6031 VGND VGND VPWR VPWR net6034 sky130_fd_sc_hd__buf_1
Xwire5300 net5301 VGND VGND VPWR VPWR net5300 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5311 net5312 VGND VGND VPWR VPWR net5311 sky130_fd_sc_hd__buf_1
X_24237_ net1015 net1658 VGND VGND VPWR VPWR _04098_ sky130_fd_sc_hd__nor2_1
Xwire5322 net5323 VGND VGND VPWR VPWR net5322 sky130_fd_sc_hd__clkbuf_1
X_21449_ _01349_ VGND VGND VPWR VPWR _01462_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_39_Left_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire6067 net6064 VGND VGND VPWR VPWR net6067 sky130_fd_sc_hd__clkbuf_2
Xwire5333 net5334 VGND VGND VPWR VPWR net5333 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5344 net5345 VGND VGND VPWR VPWR net5344 sky130_fd_sc_hd__clkbuf_1
Xwire4610 net4613 VGND VGND VPWR VPWR net4610 sky130_fd_sc_hd__buf_1
Xwire5355 net5356 VGND VGND VPWR VPWR net5355 sky130_fd_sc_hd__clkbuf_1
Xwire4621 net4622 VGND VGND VPWR VPWR net4621 sky130_fd_sc_hd__clkbuf_1
X_24168_ _04029_ _03948_ pid_q.prev_error\[7\] VGND VGND VPWR VPWR _04030_ sky130_fd_sc_hd__o21ba_1
Xwire5366 pid_d.out\[1\] VGND VGND VPWR VPWR net5366 sky130_fd_sc_hd__clkbuf_2
Xwire4632 net4633 VGND VGND VPWR VPWR net4632 sky130_fd_sc_hd__clkbuf_1
Xwire5377 net5378 VGND VGND VPWR VPWR net5377 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4643 net4644 VGND VGND VPWR VPWR net4643 sky130_fd_sc_hd__clkbuf_1
Xwire5399 net5400 VGND VGND VPWR VPWR net5399 sky130_fd_sc_hd__buf_1
X_23119_ _02973_ _02978_ VGND VGND VPWR VPWR _02989_ sky130_fd_sc_hd__xnor2_1
Xwire4665 net4666 VGND VGND VPWR VPWR net4665 sky130_fd_sc_hd__buf_1
Xwire3920 net3921 VGND VGND VPWR VPWR net3920 sky130_fd_sc_hd__clkbuf_2
Xwire4676 net4673 VGND VGND VPWR VPWR net4676 sky130_fd_sc_hd__buf_1
Xwire3931 _10122_ VGND VGND VPWR VPWR net3931 sky130_fd_sc_hd__buf_1
X_24099_ _03941_ _03960_ VGND VGND VPWR VPWR _03961_ sky130_fd_sc_hd__nand2_1
X_16990_ net1809 VGND VGND VPWR VPWR _08952_ sky130_fd_sc_hd__buf_1
Xwire3942 _09910_ VGND VGND VPWR VPWR net3942 sky130_fd_sc_hd__buf_1
XFILLER_0_101_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4698 net4699 VGND VGND VPWR VPWR net4698 sky130_fd_sc_hd__buf_1
Xwire3953 net3954 VGND VGND VPWR VPWR net3953 sky130_fd_sc_hd__clkbuf_1
Xwire3964 net3965 VGND VGND VPWR VPWR net3964 sky130_fd_sc_hd__buf_1
X_15941_ net425 _08009_ VGND VGND VPWR VPWR _08010_ sky130_fd_sc_hd__xnor2_1
Xwire3975 _09682_ VGND VGND VPWR VPWR net3975 sky130_fd_sc_hd__clkbuf_1
Xwire3986 net3987 VGND VGND VPWR VPWR net3986 sky130_fd_sc_hd__buf_1
Xwire3997 _09606_ VGND VGND VPWR VPWR net3997 sky130_fd_sc_hd__buf_2
X_18660_ net422 _10503_ _10505_ VGND VGND VPWR VPWR _10507_ sky130_fd_sc_hd__a21o_1
X_15872_ net2842 net3432 net3390 net2683 net3523 VGND VGND VPWR VPWR _07941_ sky130_fd_sc_hd__a32o_1
X_17611_ net6695 _09490_ svm0.tB\[8\] net4025 _09491_ VGND VGND VPWR VPWR _09492_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_99_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14823_ net4285 VGND VGND VPWR VPWR _06928_ sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_48_Left_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18591_ net2539 _10438_ VGND VGND VPWR VPWR _10439_ sky130_fd_sc_hd__xnor2_2
X_17542_ net6691 _09421_ _09422_ _09423_ VGND VGND VPWR VPWR _09424_ sky130_fd_sc_hd__a211o_1
XFILLER_0_153_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length8671 net8672 VGND VGND VPWR VPWR net8671 sky130_fd_sc_hd__buf_1
Xmax_length8682 net8683 VGND VGND VPWR VPWR net8682 sky130_fd_sc_hd__buf_1
X_14754_ net8974 net2870 net1906 VGND VGND VPWR VPWR _00157_ sky130_fd_sc_hd__a21bo_1
X_13705_ net7697 net3685 net2967 VGND VGND VPWR VPWR _05974_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17473_ net4020 net2569 _09363_ _09365_ VGND VGND VPWR VPWR _00396_ sky130_fd_sc_hd__a31o_1
X_14685_ matmul0.sin\[4\] _06833_ VGND VGND VPWR VPWR _06834_ sky130_fd_sc_hd__xnor2_1
X_19212_ net6258 net6313 VGND VGND VPWR VPWR _11049_ sky130_fd_sc_hd__and2_1
X_13636_ _05900_ _05905_ VGND VGND VPWR VPWR _05906_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16424_ net490 _08484_ _08428_ _08381_ VGND VGND VPWR VPWR _08486_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_6_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19143_ net6232 net3908 _10979_ net3206 _10804_ VGND VGND VPWR VPWR _10980_ sky130_fd_sc_hd__a221o_1
X_13567_ net7865 net1577 _05710_ VGND VGND VPWR VPWR _05838_ sky130_fd_sc_hd__and3_1
X_16355_ _08416_ _08417_ VGND VGND VPWR VPWR _08418_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15306_ _06968_ net3598 _07379_ VGND VGND VPWR VPWR _07380_ sky130_fd_sc_hd__o21a_1
XFILLER_0_124_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19074_ _10827_ VGND VGND VPWR VPWR _10911_ sky130_fd_sc_hd__buf_1
X_16286_ _08348_ _08349_ VGND VGND VPWR VPWR _08350_ sky130_fd_sc_hd__nor2_1
X_13498_ net578 net785 VGND VGND VPWR VPWR _05771_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_57_Left_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18025_ net6918 VGND VGND VPWR VPWR _09876_ sky130_fd_sc_hd__inv_2
Xwire7280 net7281 VGND VGND VPWR VPWR net7280 sky130_fd_sc_hd__buf_1
XFILLER_0_1_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15237_ net1881 net1879 VGND VGND VPWR VPWR _07311_ sky130_fd_sc_hd__xnor2_1
Xwire7291 net7292 VGND VGND VPWR VPWR net7291 sky130_fd_sc_hd__buf_1
XFILLER_0_140_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout5783 net5786 VGND VGND VPWR VPWR net5783 sky130_fd_sc_hd__buf_1
X_15168_ net2730 net2729 VGND VGND VPWR VPWR _07242_ sky130_fd_sc_hd__nand2_1
X_14119_ _06379_ _06380_ VGND VGND VPWR VPWR _06381_ sky130_fd_sc_hd__xnor2_1
X_15099_ net4163 net4159 net4169 net4164 VGND VGND VPWR VPWR _07173_ sky130_fd_sc_hd__o22a_1
X_19976_ net5999 net2092 VGND VGND VPWR VPWR _11807_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18927_ net275 _10747_ net6376 VGND VGND VPWR VPWR _10767_ sky130_fd_sc_hd__o21a_1
XFILLER_0_157_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18858_ _10686_ _10688_ VGND VGND VPWR VPWR _10700_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_66_Left_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17809_ net6982 VGND VGND VPWR VPWR _09660_ sky130_fd_sc_hd__inv_2
X_18789_ net3967 _10580_ _10579_ VGND VGND VPWR VPWR _10633_ sky130_fd_sc_hd__mux2_1
X_20820_ _12555_ _12557_ _00835_ VGND VGND VPWR VPWR _00836_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20751_ net5546 net5873 VGND VGND VPWR VPWR _12522_ sky130_fd_sc_hd__nand2_1
Xwire8909 net8915 VGND VGND VPWR VPWR net8909 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23470_ net4619 net4996 VGND VGND VPWR VPWR _03339_ sky130_fd_sc_hd__nand2_1
XFILLER_0_174_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20682_ _12454_ _12457_ VGND VGND VPWR VPWR _12458_ sky130_fd_sc_hd__and2_1
Xmax_length4629 net4623 VGND VGND VPWR VPWR net4629 sky130_fd_sc_hd__buf_1
XFILLER_0_162_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22421_ _02421_ _02422_ VGND VGND VPWR VPWR _02423_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_75_Left_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3939 _10045_ VGND VGND VPWR VPWR net3939 sky130_fd_sc_hd__clkbuf_1
X_25140_ clknet_leaf_50_clk _00029_ net8757 VGND VGND VPWR VPWR svm0.tC\[12\] sky130_fd_sc_hd__dfrtp_1
X_22352_ _02353_ _02354_ VGND VGND VPWR VPWR _02355_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21303_ _00862_ _00868_ _00864_ net3796 VGND VGND VPWR VPWR _01318_ sky130_fd_sc_hd__a211o_1
XFILLER_0_171_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25071_ net4418 net5176 VGND VGND VPWR VPWR _04818_ sky130_fd_sc_hd__xor2_1
X_22283_ _02285_ _02286_ VGND VGND VPWR VPWR _02287_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24022_ _03876_ _03884_ VGND VGND VPWR VPWR _03885_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_14_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold230 matmul0.a\[13\] VGND VGND VPWR VPWR net9183 sky130_fd_sc_hd__dlygate4sd3_1
X_21234_ _01247_ _01248_ VGND VGND VPWR VPWR _01249_ sky130_fd_sc_hd__xnor2_1
Xhold241 svm0.tC\[15\] VGND VGND VPWR VPWR net9194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 pid_d.prev_int\[9\] VGND VGND VPWR VPWR net9205 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3205 net3206 VGND VGND VPWR VPWR net3205 sky130_fd_sc_hd__buf_1
Xwire3216 net3217 VGND VGND VPWR VPWR net3216 sky130_fd_sc_hd__clkbuf_2
Xhold263 cordic0.slte0.opA\[17\] VGND VGND VPWR VPWR net9216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 matmul0.a\[9\] VGND VGND VPWR VPWR net9227 sky130_fd_sc_hd__dlygate4sd3_1
X_21165_ _01168_ _01169_ VGND VGND VPWR VPWR _01181_ sky130_fd_sc_hd__or2_1
Xwire3227 _10165_ VGND VGND VPWR VPWR net3227 sky130_fd_sc_hd__clkbuf_1
Xhold285 matmul0.beta_pass\[5\] VGND VGND VPWR VPWR net9238 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3238 _09802_ VGND VGND VPWR VPWR net3238 sky130_fd_sc_hd__buf_1
Xwire2504 net2505 VGND VGND VPWR VPWR net2504 sky130_fd_sc_hd__clkbuf_2
Xwire3249 net3250 VGND VGND VPWR VPWR net3249 sky130_fd_sc_hd__clkbuf_1
Xwire2515 _11127_ VGND VGND VPWR VPWR net2515 sky130_fd_sc_hd__buf_1
Xwire2526 _10894_ VGND VGND VPWR VPWR net2526 sky130_fd_sc_hd__clkbuf_1
X_20116_ net6079 _11943_ VGND VGND VPWR VPWR _11944_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21096_ _01104_ _01110_ _01111_ VGND VGND VPWR VPWR _01112_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_84_Left_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1803 _09010_ VGND VGND VPWR VPWR net1803 sky130_fd_sc_hd__clkbuf_1
Xwire2548 _09931_ VGND VGND VPWR VPWR net2548 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_102_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1814 net1815 VGND VGND VPWR VPWR net1814 sky130_fd_sc_hd__clkbuf_1
Xwire2559 net2560 VGND VGND VPWR VPWR net2559 sky130_fd_sc_hd__clkbuf_2
Xwire1825 net1826 VGND VGND VPWR VPWR net1825 sky130_fd_sc_hd__buf_1
X_24924_ net8868 net140 VGND VGND VPWR VPWR _04710_ sky130_fd_sc_hd__and2b_1
Xwire1836 net1837 VGND VGND VPWR VPWR net1836 sky130_fd_sc_hd__clkbuf_1
X_20047_ net9038 net1202 _11876_ net1771 VGND VGND VPWR VPWR _00460_ sky130_fd_sc_hd__a22o_1
XFILLER_0_176_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1847 net1848 VGND VGND VPWR VPWR net1847 sky130_fd_sc_hd__clkbuf_1
Xwire1858 _07600_ VGND VGND VPWR VPWR net1858 sky130_fd_sc_hd__clkbuf_1
Xwire1869 net1870 VGND VGND VPWR VPWR net1869 sky130_fd_sc_hd__dlymetal6s2s_1
X_24855_ _04660_ net4779 net2003 VGND VGND VPWR VPWR _04661_ sky130_fd_sc_hd__mux2_1
Xmax_length7211 net7212 VGND VGND VPWR VPWR net7211 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23806_ pid_q.curr_int\[4\] VGND VGND VPWR VPWR _03671_ sky130_fd_sc_hd__inv_2
X_24786_ _04608_ _04607_ _04609_ VGND VGND VPWR VPWR _04612_ sky130_fd_sc_hd__a21bo_1
X_21998_ _02003_ _02005_ VGND VGND VPWR VPWR _02006_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23737_ _03601_ _03602_ VGND VGND VPWR VPWR _03603_ sky130_fd_sc_hd__xnor2_1
Xmax_length6543 net6539 VGND VGND VPWR VPWR net6543 sky130_fd_sc_hd__buf_1
X_20949_ _00920_ _00964_ net3840 VGND VGND VPWR VPWR _00965_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_80_clk clknet_4_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_80_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14470_ net7361 net5305 VGND VGND VPWR VPWR _06657_ sky130_fd_sc_hd__or2_1
X_23668_ _03532_ _03534_ VGND VGND VPWR VPWR _03535_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_93_Left_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13421_ net7921 net1929 _05692_ VGND VGND VPWR VPWR _05694_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22619_ net7218 _02586_ VGND VGND VPWR VPWR _02590_ sky130_fd_sc_hd__or2_1
X_25407_ clknet_leaf_72_clk _00290_ net8465 VGND VGND VPWR VPWR matmul0.a\[10\] sky130_fd_sc_hd__dfrtp_1
X_23599_ _03465_ net1020 VGND VGND VPWR VPWR _03467_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16140_ _08200_ _08205_ VGND VGND VPWR VPWR _08206_ sky130_fd_sc_hd__xnor2_1
X_13352_ _05623_ _05624_ VGND VGND VPWR VPWR _05625_ sky130_fd_sc_hd__and2b_1
X_25338_ clknet_leaf_84_clk _00221_ net8506 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16071_ net776 _08137_ VGND VGND VPWR VPWR _08138_ sky130_fd_sc_hd__xnor2_2
X_13283_ net1575 VGND VGND VPWR VPWR _05556_ sky130_fd_sc_hd__clkbuf_1
X_25269_ clknet_leaf_88_clk _00152_ net8421 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.b\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire5130 net5131 VGND VGND VPWR VPWR net5130 sky130_fd_sc_hd__clkbuf_1
Xfanout4334 net4340 VGND VGND VPWR VPWR net4334 sky130_fd_sc_hd__clkbuf_1
X_15022_ _06998_ VGND VGND VPWR VPWR _07096_ sky130_fd_sc_hd__buf_1
Xwire5152 net5153 VGND VGND VPWR VPWR net5152 sky130_fd_sc_hd__clkbuf_1
Xwire5163 net5164 VGND VGND VPWR VPWR net5163 sky130_fd_sc_hd__buf_1
XFILLER_0_47_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5174 net5175 VGND VGND VPWR VPWR net5174 sky130_fd_sc_hd__clkbuf_2
Xwire4440 net4441 VGND VGND VPWR VPWR net4440 sky130_fd_sc_hd__clkbuf_1
Xwire5185 net5186 VGND VGND VPWR VPWR net5185 sky130_fd_sc_hd__buf_1
X_19830_ _11608_ _11606_ VGND VGND VPWR VPWR _11664_ sky130_fd_sc_hd__or2b_1
Xwire5196 net5197 VGND VGND VPWR VPWR net5196 sky130_fd_sc_hd__clkbuf_1
Xwire4473 net4474 VGND VGND VPWR VPWR net4473 sky130_fd_sc_hd__clkbuf_1
Xwire4484 net4485 VGND VGND VPWR VPWR net4484 sky130_fd_sc_hd__buf_1
Xwire4495 net4496 VGND VGND VPWR VPWR net4495 sky130_fd_sc_hd__buf_1
Xwire3750 net3751 VGND VGND VPWR VPWR net3750 sky130_fd_sc_hd__clkbuf_1
Xwire3761 net3762 VGND VGND VPWR VPWR net3761 sky130_fd_sc_hd__buf_1
X_19761_ _11517_ _11524_ _11595_ VGND VGND VPWR VPWR _11596_ sky130_fd_sc_hd__o21ai_1
X_16973_ _08925_ _08935_ VGND VGND VPWR VPWR _08936_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3772 net3773 VGND VGND VPWR VPWR net3772 sky130_fd_sc_hd__clkbuf_1
Xwire3783 net3784 VGND VGND VPWR VPWR net3783 sky130_fd_sc_hd__clkbuf_1
Xwire3794 net3795 VGND VGND VPWR VPWR net3794 sky130_fd_sc_hd__clkbuf_1
X_18712_ _10554_ _10557_ VGND VGND VPWR VPWR _10558_ sky130_fd_sc_hd__and2_1
X_15924_ _07989_ _07991_ _07992_ VGND VGND VPWR VPWR _07993_ sky130_fd_sc_hd__o21ba_1
X_19692_ _11458_ net2101 _11527_ VGND VGND VPWR VPWR _11528_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 angle_in[2] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
X_18643_ net6770 net6792 net2539 _10436_ VGND VGND VPWR VPWR _10490_ sky130_fd_sc_hd__or4_1
XFILLER_0_188_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15855_ _07831_ _07919_ _07920_ VGND VGND VPWR VPWR _07924_ sky130_fd_sc_hd__o21a_1
X_14806_ net3626 net7175 net3622 VGND VGND VPWR VPWR _06920_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18574_ _10171_ _10364_ net3308 net6934 VGND VGND VPWR VPWR _10422_ sky130_fd_sc_hd__a211o_1
X_15786_ _07850_ _07855_ VGND VGND VPWR VPWR _07856_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12998_ _05178_ _05179_ VGND VGND VPWR VPWR _05271_ sky130_fd_sc_hd__or2_1
X_17525_ net6742 _09405_ net6694 VGND VGND VPWR VPWR _09409_ sky130_fd_sc_hd__a21o_1
X_14737_ net7158 _06871_ VGND VGND VPWR VPWR _06872_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_71_clk clknet_4_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_129_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17456_ net3274 _09350_ net6662 VGND VGND VPWR VPWR _09351_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14668_ net3630 VGND VGND VPWR VPWR _06820_ sky130_fd_sc_hd__buf_1
X_16407_ net2654 net2209 VGND VGND VPWR VPWR _08469_ sky130_fd_sc_hd__nand2_1
X_13619_ _05791_ _05796_ VGND VGND VPWR VPWR _05889_ sky130_fd_sc_hd__or2_1
X_17387_ svm0.delta\[6\] VGND VGND VPWR VPWR _09295_ sky130_fd_sc_hd__inv_2
XFILLER_0_184_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14599_ _06768_ _06772_ VGND VGND VPWR VPWR _06773_ sky130_fd_sc_hd__xnor2_1
X_19126_ net3910 _10791_ VGND VGND VPWR VPWR _10963_ sky130_fd_sc_hd__nor2_1
X_16338_ _08399_ _08400_ VGND VGND VPWR VPWR _08401_ sky130_fd_sc_hd__nand2_1
X_19057_ net6314 _10829_ net3211 VGND VGND VPWR VPWR _10894_ sky130_fd_sc_hd__o21ai_1
X_16269_ _08323_ _08332_ VGND VGND VPWR VPWR _08333_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_168_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18008_ _09641_ _09858_ VGND VGND VPWR VPWR _09859_ sky130_fd_sc_hd__xnor2_2
Xfanout5580 net5586 VGND VGND VPWR VPWR net5580 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19959_ _11755_ _11758_ net3153 net6107 VGND VGND VPWR VPWR _11790_ sky130_fd_sc_hd__a211o_1
X_22970_ matmul0.beta_pass\[4\] net1838 net6567 VGND VGND VPWR VPWR _02853_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21921_ net5693 net5514 VGND VGND VPWR VPWR _01929_ sky130_fd_sc_hd__nand2_1
XFILLER_0_179_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24640_ net2016 _04493_ _04494_ VGND VGND VPWR VPWR _04495_ sky130_fd_sc_hd__a21o_1
X_21852_ _01770_ _01773_ _01767_ VGND VGND VPWR VPWR _01861_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_132_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20803_ net5913 net5455 VGND VGND VPWR VPWR _00819_ sky130_fd_sc_hd__nand2_1
X_24571_ _04425_ _04426_ VGND VGND VPWR VPWR _04427_ sky130_fd_sc_hd__xnor2_1
X_21783_ net1172 _01792_ VGND VGND VPWR VPWR _01793_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_62_clk clknet_4_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_62_clk sky130_fd_sc_hd__clkbuf_16
X_23522_ pid_q.curr_int\[0\] pid_q.prev_int\[0\] pid_q.prev_int\[1\] pid_q.curr_int\[1\]
+ VGND VGND VPWR VPWR _03390_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20734_ net5524 net5838 VGND VGND VPWR VPWR _12505_ sky130_fd_sc_hd__nand2_1
Xwire8706 net8707 VGND VGND VPWR VPWR net8706 sky130_fd_sc_hd__buf_1
Xwire8728 net8729 VGND VGND VPWR VPWR net8728 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_9_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8739 net8740 VGND VGND VPWR VPWR net8739 sky130_fd_sc_hd__clkbuf_1
X_23453_ net4597 net5024 VGND VGND VPWR VPWR _03322_ sky130_fd_sc_hd__nand2_2
X_20665_ net6483 _12441_ VGND VGND VPWR VPWR _12442_ sky130_fd_sc_hd__nand2_1
XFILLER_0_163_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire418 net419 VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__clkbuf_1
X_22404_ _02402_ _02405_ VGND VGND VPWR VPWR _02406_ sky130_fd_sc_hd__xor2_1
XFILLER_0_45_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire429 net430 VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__clkbuf_1
Xmax_length3736 _04117_ VGND VGND VPWR VPWR net3736 sky130_fd_sc_hd__buf_1
XFILLER_0_34_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23384_ _03245_ _03253_ VGND VGND VPWR VPWR _03254_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_162_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length3758 _02866_ VGND VGND VPWR VPWR net3758 sky130_fd_sc_hd__buf_1
X_20596_ net6756 _09035_ _12377_ net2609 VGND VGND VPWR VPWR _12378_ sky130_fd_sc_hd__a22oi_1
X_25123_ net9224 net3033 _04852_ pid_d.curr_int\[11\] VGND VGND VPWR VPWR _00804_
+ sky130_fd_sc_hd__a22o_1
X_22335_ _02320_ _02318_ _02321_ VGND VGND VPWR VPWR _02338_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_21_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25054_ pid_q.out\[8\] net1995 _04802_ VGND VGND VPWR VPWR _04804_ sky130_fd_sc_hd__nor3_1
X_22266_ pid_d.curr_int\[11\] VGND VGND VPWR VPWR _02270_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24005_ net795 _03835_ VGND VGND VPWR VPWR _03868_ sky130_fd_sc_hd__nand2_1
Xwire3002 _00000_ VGND VGND VPWR VPWR net3002 sky130_fd_sc_hd__clkbuf_1
X_21217_ _00938_ _00968_ VGND VGND VPWR VPWR _01233_ sky130_fd_sc_hd__xnor2_1
Xwire3013 net3014 VGND VGND VPWR VPWR net3013 sky130_fd_sc_hd__clkbuf_1
Xwire3024 net3025 VGND VGND VPWR VPWR net3024 sky130_fd_sc_hd__clkbuf_1
X_22197_ net1708 _02201_ VGND VGND VPWR VPWR _02202_ sky130_fd_sc_hd__xnor2_1
Xwire3035 net3036 VGND VGND VPWR VPWR net3035 sky130_fd_sc_hd__clkbuf_1
Xwire2301 net2302 VGND VGND VPWR VPWR net2301 sky130_fd_sc_hd__buf_1
Xwire3046 net3047 VGND VGND VPWR VPWR net3046 sky130_fd_sc_hd__buf_1
Xwire3057 net3058 VGND VGND VPWR VPWR net3057 sky130_fd_sc_hd__clkbuf_1
Xwire2312 net2313 VGND VGND VPWR VPWR net2312 sky130_fd_sc_hd__buf_1
X_21148_ _01161_ _01163_ VGND VGND VPWR VPWR _01164_ sky130_fd_sc_hd__xnor2_1
Xwire3068 _02684_ VGND VGND VPWR VPWR net3068 sky130_fd_sc_hd__buf_1
Xwire2323 net2324 VGND VGND VPWR VPWR net2323 sky130_fd_sc_hd__buf_1
Xwire2334 _04957_ VGND VGND VPWR VPWR net2334 sky130_fd_sc_hd__buf_1
Xwire1600 net1601 VGND VGND VPWR VPWR net1600 sky130_fd_sc_hd__clkbuf_1
Xwire2345 _04923_ VGND VGND VPWR VPWR net2345 sky130_fd_sc_hd__buf_1
Xwire2356 net2357 VGND VGND VPWR VPWR net2356 sky130_fd_sc_hd__buf_1
Xwire1611 net1612 VGND VGND VPWR VPWR net1611 sky130_fd_sc_hd__clkbuf_2
X_13970_ _06117_ net7604 VGND VGND VPWR VPWR _06235_ sky130_fd_sc_hd__and2_1
Xwire2367 _04899_ VGND VGND VPWR VPWR net2367 sky130_fd_sc_hd__buf_1
Xwire1622 net1623 VGND VGND VPWR VPWR net1622 sky130_fd_sc_hd__buf_1
X_21079_ _01088_ _01090_ VGND VGND VPWR VPWR _01095_ sky130_fd_sc_hd__nand2_1
Xwire2378 _04891_ VGND VGND VPWR VPWR net2378 sky130_fd_sc_hd__buf_1
Xwire1633 _04752_ VGND VGND VPWR VPWR net1633 sky130_fd_sc_hd__buf_1
Xwire2389 net2390 VGND VGND VPWR VPWR net2389 sky130_fd_sc_hd__buf_1
Xwire1655 _04139_ VGND VGND VPWR VPWR net1655 sky130_fd_sc_hd__buf_1
X_24907_ net8869 net121 net123 net126 VGND VGND VPWR VPWR _04697_ sky130_fd_sc_hd__or4_1
Xwire1666 _03505_ VGND VGND VPWR VPWR net1666 sky130_fd_sc_hd__buf_1
X_12921_ net7931 net1958 net1957 _05111_ VGND VGND VPWR VPWR _05194_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_38_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25887_ clknet_leaf_40_clk _00760_ net8769 VGND VGND VPWR VPWR pid_q.ki\[15\] sky130_fd_sc_hd__dfrtp_1
Xwire1677 _02983_ VGND VGND VPWR VPWR net1677 sky130_fd_sc_hd__buf_1
Xwire1688 net1689 VGND VGND VPWR VPWR net1688 sky130_fd_sc_hd__clkbuf_2
Xwire1699 net1700 VGND VGND VPWR VPWR net1699 sky130_fd_sc_hd__buf_1
X_15640_ _07590_ _07625_ _07711_ VGND VGND VPWR VPWR _07712_ sky130_fd_sc_hd__o21ai_2
X_24838_ net7482 net690 _04035_ VGND VGND VPWR VPWR _04652_ sky130_fd_sc_hd__a21o_1
X_12852_ _05068_ _05069_ _05067_ VGND VGND VPWR VPWR _05125_ sky130_fd_sc_hd__a21boi_1
X_12783_ _05055_ VGND VGND VPWR VPWR _05056_ sky130_fd_sc_hd__clkbuf_1
X_15571_ _07633_ _07631_ VGND VGND VPWR VPWR _07643_ sky130_fd_sc_hd__and2b_1
X_24769_ _04596_ _04593_ net5235 VGND VGND VPWR VPWR _04597_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_53_clk clknet_4_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_150_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17310_ net6709 net7719 VGND VGND VPWR VPWR _09224_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14522_ _06692_ _06695_ _06701_ net7302 net2389 VGND VGND VPWR VPWR _06702_ sky130_fd_sc_hd__o221a_1
X_18290_ net3245 net1215 _10140_ VGND VGND VPWR VPWR _10141_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_127_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17241_ net3387 _09186_ _09187_ VGND VGND VPWR VPWR _09188_ sky130_fd_sc_hd__mux2_1
X_14453_ net5192 net1550 net3648 net4394 _06643_ VGND VGND VPWR VPWR _06644_ sky130_fd_sc_hd__a221o_1
XFILLER_0_83_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length5694 net5689 VGND VGND VPWR VPWR net5694 sky130_fd_sc_hd__buf_1
XFILLER_0_37_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13404_ _05668_ net581 net583 VGND VGND VPWR VPWR _05677_ sky130_fd_sc_hd__o21bai_1
Xwire930 net931 VGND VGND VPWR VPWR net930 sky130_fd_sc_hd__buf_1
X_14384_ net8280 net3637 VGND VGND VPWR VPWR _06591_ sky130_fd_sc_hd__and2_1
X_17172_ net1076 _09123_ VGND VGND VPWR VPWR _09124_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4993 net4994 VGND VGND VPWR VPWR net4993 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire941 net942 VGND VGND VPWR VPWR net941 sky130_fd_sc_hd__buf_1
XFILLER_0_135_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire952 _11977_ VGND VGND VPWR VPWR net952 sky130_fd_sc_hd__buf_1
X_13335_ net2304 VGND VGND VPWR VPWR _05608_ sky130_fd_sc_hd__buf_1
XFILLER_0_49_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16123_ net2656 net2764 VGND VGND VPWR VPWR _08189_ sky130_fd_sc_hd__nor2_1
Xwire963 _09824_ VGND VGND VPWR VPWR net963 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire974 _08696_ VGND VGND VPWR VPWR net974 sky130_fd_sc_hd__clkbuf_1
Xwire985 net986 VGND VGND VPWR VPWR net985 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire996 _06070_ VGND VGND VPWR VPWR net996 sky130_fd_sc_hd__buf_1
X_13266_ _05417_ _05418_ VGND VGND VPWR VPWR _05539_ sky130_fd_sc_hd__and2_1
X_16054_ net2652 net2764 VGND VGND VPWR VPWR _08121_ sky130_fd_sc_hd__nor2_2
XFILLER_0_11_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15005_ net2831 _07078_ net3553 net3545 VGND VGND VPWR VPWR _07079_ sky130_fd_sc_hd__a211o_1
X_13197_ _05466_ _05469_ VGND VGND VPWR VPWR _05470_ sky130_fd_sc_hd__xor2_1
Xwire4270 net4271 VGND VGND VPWR VPWR net4270 sky130_fd_sc_hd__clkbuf_1
X_19813_ _11645_ _10975_ _11453_ _11646_ VGND VGND VPWR VPWR _11647_ sky130_fd_sc_hd__a211o_1
Xwire4281 net4286 VGND VGND VPWR VPWR net4281 sky130_fd_sc_hd__buf_1
Xwire4292 _04876_ VGND VGND VPWR VPWR net4292 sky130_fd_sc_hd__buf_1
XFILLER_0_138_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3580 net3581 VGND VGND VPWR VPWR net3580 sky130_fd_sc_hd__buf_1
XFILLER_0_194_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19744_ _11577_ _11578_ VGND VGND VPWR VPWR _11579_ sky130_fd_sc_hd__nand2_1
X_16956_ _08838_ net1808 VGND VGND VPWR VPWR _08919_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire3591 net3593 VGND VGND VPWR VPWR net3591 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2890 _06603_ VGND VGND VPWR VPWR net2890 sky130_fd_sc_hd__buf_1
X_15907_ _07970_ net1522 VGND VGND VPWR VPWR _07976_ sky130_fd_sc_hd__xor2_1
X_19675_ net3162 _11177_ _11466_ VGND VGND VPWR VPWR _11511_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_139_Right_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16887_ net5989 net2612 _08850_ VGND VGND VPWR VPWR _08851_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18626_ net6999 net3296 net6920 VGND VGND VPWR VPWR _10473_ sky130_fd_sc_hd__or3_1
XFILLER_0_189_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15838_ _07906_ _07907_ VGND VGND VPWR VPWR _07908_ sky130_fd_sc_hd__nor2_1
X_18557_ _10334_ _10339_ _10397_ VGND VGND VPWR VPWR _10405_ sky130_fd_sc_hd__and3_1
X_15769_ net2700 net2671 net3526 VGND VGND VPWR VPWR _07839_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_44_clk clknet_4_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_188_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17508_ _09311_ _09388_ _09394_ VGND VGND VPWR VPWR _09395_ sky130_fd_sc_hd__a21o_1
X_18488_ _10249_ _10254_ _10337_ VGND VGND VPWR VPWR _10338_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17439_ net6744 _09335_ VGND VGND VPWR VPWR _09336_ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20450_ net950 _12232_ _12241_ _08857_ _12242_ VGND VGND VPWR VPWR _12243_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19109_ net6226 VGND VGND VPWR VPWR _10946_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20381_ net949 _12178_ _12179_ VGND VGND VPWR VPWR _12180_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_179_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22120_ _02122_ _02125_ VGND VGND VPWR VPWR _02126_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22051_ _01966_ _02055_ VGND VGND VPWR VPWR _02058_ sky130_fd_sc_hd__nor2_1
X_21002_ _00996_ _01016_ _01017_ VGND VGND VPWR VPWR _01018_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25810_ clknet_leaf_36_clk _00683_ net8797 VGND VGND VPWR VPWR pid_q.prev_error\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25741_ clknet_leaf_13_clk _00614_ net8608 VGND VGND VPWR VPWR pid_d.ki\[15\] sky130_fd_sc_hd__dfrtp_1
X_22953_ _02388_ _02838_ _02840_ VGND VGND VPWR VPWR _02841_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_106_Right_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21904_ _01910_ _01911_ VGND VGND VPWR VPWR _01913_ sky130_fd_sc_hd__or2_1
X_25672_ clknet_leaf_4_clk _00545_ net8567 VGND VGND VPWR VPWR pid_d.prev_error\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22884_ _01917_ _02770_ _02778_ VGND VGND VPWR VPWR _02779_ sky130_fd_sc_hd__a21o_1
XFILLER_0_179_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24623_ net4503 net4807 VGND VGND VPWR VPWR _04478_ sky130_fd_sc_hd__nand2_1
X_21835_ _01755_ _01760_ _01753_ VGND VGND VPWR VPWR _01844_ sky130_fd_sc_hd__a21bo_1
Xclkbuf_leaf_35_clk clknet_4_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_16
X_24554_ _04408_ _04409_ VGND VGND VPWR VPWR _04410_ sky130_fd_sc_hd__and2b_1
X_21766_ _01762_ _01775_ VGND VGND VPWR VPWR _01776_ sky130_fd_sc_hd__xnor2_1
Xwire8503 net8504 VGND VGND VPWR VPWR net8503 sky130_fd_sc_hd__clkbuf_2
Xwire8514 net8515 VGND VGND VPWR VPWR net8514 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23505_ net3750 net3050 VGND VGND VPWR VPWR _03374_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20717_ net2583 _12269_ _12479_ VGND VGND VPWR VPWR _12489_ sky130_fd_sc_hd__a21o_1
Xwire8525 net8526 VGND VGND VPWR VPWR net8525 sky130_fd_sc_hd__clkbuf_1
X_24485_ _04298_ _04304_ _04341_ net4873 VGND VGND VPWR VPWR _04342_ sky130_fd_sc_hd__a2bb2o_2
Xwire8536 net8530 VGND VGND VPWR VPWR net8536 sky130_fd_sc_hd__clkbuf_1
Xwire7802 net7803 VGND VGND VPWR VPWR net7802 sky130_fd_sc_hd__buf_1
X_21697_ net1174 _01707_ VGND VGND VPWR VPWR _01708_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_53_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8547 net8548 VGND VGND VPWR VPWR net8547 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire204 _02516_ VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_1
Xwire7813 net7819 VGND VGND VPWR VPWR net7813 sky130_fd_sc_hd__buf_1
Xwire8558 net8559 VGND VGND VPWR VPWR net8558 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7824 net7825 VGND VGND VPWR VPWR net7824 sky130_fd_sc_hd__buf_1
XFILLER_0_19_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3511 net3512 VGND VGND VPWR VPWR net3511 sky130_fd_sc_hd__buf_1
X_23436_ net749 net796 VGND VGND VPWR VPWR _03306_ sky130_fd_sc_hd__xnor2_1
Xmax_length4267 _04928_ VGND VGND VPWR VPWR net4267 sky130_fd_sc_hd__clkbuf_1
Xwire215 net216 VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_1
Xwire226 _06011_ VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__clkbuf_1
X_20648_ net6757 net2597 _09082_ net3124 VGND VGND VPWR VPWR _12426_ sky130_fd_sc_hd__a22o_1
Xwire7846 net7848 VGND VGND VPWR VPWR net7846 sky130_fd_sc_hd__clkbuf_1
Xwire237 _04320_ VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__clkbuf_1
Xwire7857 net7858 VGND VGND VPWR VPWR net7857 sky130_fd_sc_hd__clkbuf_1
Xwire248 net249 VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7868 net7856 VGND VGND VPWR VPWR net7868 sky130_fd_sc_hd__buf_1
Xwire259 net260 VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__buf_1
Xmax_length3555 _07042_ VGND VGND VPWR VPWR net3555 sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_length2810 net2812 VGND VGND VPWR VPWR net2810 sky130_fd_sc_hd__clkbuf_1
Xwire7879 net7878 VGND VGND VPWR VPWR net7879 sky130_fd_sc_hd__clkbuf_1
X_23367_ _03231_ _03235_ VGND VGND VPWR VPWR _03237_ sky130_fd_sc_hd__nor2_1
Xmax_length3577 net3578 VGND VGND VPWR VPWR net3577 sky130_fd_sc_hd__buf_1
XFILLER_0_132_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20579_ net6255 _12357_ _12358_ VGND VGND VPWR VPWR _12362_ sky130_fd_sc_hd__o21ai_1
X_13120_ _05391_ _05392_ VGND VGND VPWR VPWR _05393_ sky130_fd_sc_hd__or2_1
X_22318_ _02320_ _02321_ VGND VGND VPWR VPWR _02322_ sky130_fd_sc_hd__xor2_1
X_25106_ net4393 net1633 net1627 _04847_ _04848_ VGND VGND VPWR VPWR _00792_ sky130_fd_sc_hd__a221o_1
XFILLER_0_103_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23298_ _03154_ _03151_ VGND VGND VPWR VPWR _03168_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2898 net2899 VGND VGND VPWR VPWR net2898 sky130_fd_sc_hd__buf_1
X_25037_ net3739 net1157 pid_q.out\[5\] VGND VGND VPWR VPWR _04789_ sky130_fd_sc_hd__o21ba_1
X_13051_ _05030_ _05322_ _05323_ VGND VGND VPWR VPWR _05324_ sky130_fd_sc_hd__a21o_1
X_22249_ pid_d.curr_error\[10\] VGND VGND VPWR VPWR _02254_ sky130_fd_sc_hd__inv_2
Xwire2120 _10874_ VGND VGND VPWR VPWR net2120 sky130_fd_sc_hd__clkbuf_1
X_16810_ _08795_ VGND VGND VPWR VPWR _00303_ sky130_fd_sc_hd__clkbuf_1
Xwire2131 _10277_ VGND VGND VPWR VPWR net2131 sky130_fd_sc_hd__clkbuf_2
Xwire2142 _09706_ VGND VGND VPWR VPWR net2142 sky130_fd_sc_hd__clkbuf_1
Xwire2153 _09476_ VGND VGND VPWR VPWR net2153 sky130_fd_sc_hd__buf_1
X_17790_ net7107 net7081 VGND VGND VPWR VPWR _09641_ sky130_fd_sc_hd__nor2b_2
Xwire2164 net2165 VGND VGND VPWR VPWR net2164 sky130_fd_sc_hd__buf_1
Xwire2175 _08899_ VGND VGND VPWR VPWR net2175 sky130_fd_sc_hd__clkbuf_1
Xwire1430 _10537_ VGND VGND VPWR VPWR net1430 sky130_fd_sc_hd__buf_1
Xwire1441 net1442 VGND VGND VPWR VPWR net1441 sky130_fd_sc_hd__buf_1
Xwire2186 net2187 VGND VGND VPWR VPWR net2186 sky130_fd_sc_hd__buf_1
X_16741_ net4291 VGND VGND VPWR VPWR _08759_ sky130_fd_sc_hd__clkbuf_1
X_13953_ _05873_ VGND VGND VPWR VPWR _06218_ sky130_fd_sc_hd__buf_1
Xwire1452 net1453 VGND VGND VPWR VPWR net1452 sky130_fd_sc_hd__buf_1
X_25939_ clknet_leaf_24_clk _00004_ net8588 VGND VGND VPWR VPWR pid_d.state\[3\] sky130_fd_sc_hd__dfrtp_1
Xwire2197 net2198 VGND VGND VPWR VPWR net2197 sky130_fd_sc_hd__buf_1
Xwire1463 net1464 VGND VGND VPWR VPWR net1463 sky130_fd_sc_hd__clkbuf_1
Xwire1474 net1475 VGND VGND VPWR VPWR net1474 sky130_fd_sc_hd__clkbuf_1
Xwire1485 net1486 VGND VGND VPWR VPWR net1485 sky130_fd_sc_hd__buf_1
X_12904_ net7803 _04902_ VGND VGND VPWR VPWR _05177_ sky130_fd_sc_hd__nand2_1
X_19460_ net2522 _11295_ _11296_ VGND VGND VPWR VPWR _11297_ sky130_fd_sc_hd__o21a_1
Xwire1496 net1497 VGND VGND VPWR VPWR net1496 sky130_fd_sc_hd__buf_1
X_16672_ _08704_ _08700_ matmul0.matmul_stage_inst.mult2\[7\] VGND VGND VPWR VPWR
+ _08705_ sky130_fd_sc_hd__a21bo_1
X_13884_ net283 _06146_ _06149_ _06150_ VGND VGND VPWR VPWR _06151_ sky130_fd_sc_hd__o211a_1
X_18411_ net606 _10261_ VGND VGND VPWR VPWR _10262_ sky130_fd_sc_hd__nor2_1
XFILLER_0_186_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15623_ _07377_ _07694_ _07605_ VGND VGND VPWR VPWR _07695_ sky130_fd_sc_hd__and3_1
X_12835_ net7849 _04901_ _05034_ _05036_ VGND VGND VPWR VPWR _05108_ sky130_fd_sc_hd__a22oi_4
X_19391_ net6358 _11225_ _11227_ VGND VGND VPWR VPWR _11228_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_26_clk clknet_4_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18342_ _10135_ _10132_ VGND VGND VPWR VPWR _10193_ sky130_fd_sc_hd__and2b_1
X_15554_ _07590_ _07626_ VGND VGND VPWR VPWR _07627_ sky130_fd_sc_hd__xnor2_2
X_12766_ net7784 _04920_ VGND VGND VPWR VPWR _05039_ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length6181 net6177 VGND VGND VPWR VPWR net6181 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_84_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14505_ net7302 net5262 VGND VGND VPWR VPWR _06687_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6192 net6193 VGND VGND VPWR VPWR net6192 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18273_ net3928 net3926 VGND VGND VPWR VPWR _10124_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12697_ net1343 _04969_ VGND VGND VPWR VPWR _04970_ sky130_fd_sc_hd__xnor2_1
X_15485_ _07556_ _07558_ VGND VGND VPWR VPWR _07559_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length5480 net5481 VGND VGND VPWR VPWR net5480 sky130_fd_sc_hd__buf_1
XFILLER_0_25_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17224_ _09165_ VGND VGND VPWR VPWR _09172_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14436_ net8190 net3632 VGND VGND VPWR VPWR _06631_ sky130_fd_sc_hd__and2_1
Xinput12 angle_in[5] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_1
Xinput23 currA_in[15] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput34 currB_in[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
Xinput45 currB_in[6] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
X_17155_ net3301 _09108_ VGND VGND VPWR VPWR _09109_ sky130_fd_sc_hd__nor2_1
X_14367_ _06578_ VGND VGND VPWR VPWR _00077_ sky130_fd_sc_hd__clkbuf_1
Xwire760 _01219_ VGND VGND VPWR VPWR net760 sky130_fd_sc_hd__buf_1
Xinput56 currT_in[1] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_1
Xwire771 _09266_ VGND VGND VPWR VPWR net771 sky130_fd_sc_hd__buf_1
XFILLER_0_3_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire782 _05959_ VGND VGND VPWR VPWR net782 sky130_fd_sc_hd__buf_1
Xinput67 periodTop[11] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_1
Xwire793 net794 VGND VGND VPWR VPWR net793 sky130_fd_sc_hd__buf_1
Xinput78 periodTop[7] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_1
X_16106_ net2707 _07932_ VGND VGND VPWR VPWR _08172_ sky130_fd_sc_hd__nor2_1
Xinput89 pid_d_addr[2] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_1
X_13318_ net7769 net1598 VGND VGND VPWR VPWR _05591_ sky130_fd_sc_hd__nand2_1
X_14298_ net6455 net6445 VGND VGND VPWR VPWR _06520_ sky130_fd_sc_hd__xor2_1
X_17086_ _08978_ _08979_ _09015_ _09042_ _09043_ VGND VGND VPWR VPWR _09044_ sky130_fd_sc_hd__a32o_1
XFILLER_0_58_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16037_ net1516 _08103_ VGND VGND VPWR VPWR _08104_ sky130_fd_sc_hd__xor2_1
XFILLER_0_149_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13249_ _05521_ VGND VGND VPWR VPWR _05522_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_122_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17988_ net963 _09830_ _09833_ _09838_ VGND VGND VPWR VPWR _09839_ sky130_fd_sc_hd__and4_1
X_19727_ net6030 _11449_ VGND VGND VPWR VPWR _11562_ sky130_fd_sc_hd__nand2_1
X_16939_ net4054 _08902_ cordic0.slte0.opA\[17\] VGND VGND VPWR VPWR _08903_ sky130_fd_sc_hd__a21o_1
XFILLER_0_165_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19658_ net2504 _11492_ _11493_ net3135 VGND VGND VPWR VPWR _11494_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18609_ net605 _10456_ VGND VGND VPWR VPWR _10457_ sky130_fd_sc_hd__xnor2_1
X_19589_ net653 _11424_ _11425_ VGND VGND VPWR VPWR _11426_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_17_clk clknet_4_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_16
X_21620_ _01628_ net701 VGND VGND VPWR VPWR _01632_ sky130_fd_sc_hd__and2_1
XFILLER_0_192_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21551_ net5704 net5565 VGND VGND VPWR VPWR _01563_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7109 net7106 VGND VGND VPWR VPWR net7109 sky130_fd_sc_hd__buf_1
XFILLER_0_30_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20502_ net6363 net1823 _12282_ net2086 VGND VGND VPWR VPWR _12289_ sky130_fd_sc_hd__or4_1
X_24270_ _04061_ _04063_ _04129_ VGND VGND VPWR VPWR _04130_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_56_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21482_ _01487_ _01494_ VGND VGND VPWR VPWR _01495_ sky130_fd_sc_hd__xnor2_2
Xwire6408 net6409 VGND VGND VPWR VPWR net6408 sky130_fd_sc_hd__clkbuf_1
Xwire6419 cordic0.slte0.opB\[3\] VGND VGND VPWR VPWR net6419 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23221_ net2431 _03000_ VGND VGND VPWR VPWR _03091_ sky130_fd_sc_hd__xor2_1
X_20433_ cordic0.slte0.opA\[11\] net863 _12227_ VGND VGND VPWR VPWR _12228_ sky130_fd_sc_hd__o21a_1
XFILLER_0_71_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5707 net5708 VGND VGND VPWR VPWR net5707 sky130_fd_sc_hd__buf_1
XFILLER_0_31_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5729 net5724 VGND VGND VPWR VPWR net5729 sky130_fd_sc_hd__buf_1
X_23152_ net5039 net4738 VGND VGND VPWR VPWR _03022_ sky130_fd_sc_hd__nand2_1
X_20364_ net949 _12159_ _12156_ VGND VGND VPWR VPWR _12164_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22103_ net5976 VGND VGND VPWR VPWR _02109_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23083_ _02949_ _02952_ VGND VGND VPWR VPWR _02953_ sky130_fd_sc_hd__xnor2_2
X_20295_ _12089_ _12100_ VGND VGND VPWR VPWR _12101_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22034_ net5779 net5389 VGND VGND VPWR VPWR _02041_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23985_ _03753_ net511 _03779_ VGND VGND VPWR VPWR _03849_ sky130_fd_sc_hd__and3_1
X_25724_ clknet_leaf_11_clk _00597_ net8603 VGND VGND VPWR VPWR pid_d.mult0.a\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_11_Left_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22936_ net8908 _02825_ VGND VGND VPWR VPWR _02826_ sky130_fd_sc_hd__and2_1
XFILLER_0_196_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25655_ clknet_leaf_2_clk _00528_ net8573 VGND VGND VPWR VPWR pid_d.curr_int\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22867_ _02762_ _02763_ VGND VGND VPWR VPWR _02764_ sky130_fd_sc_hd__nand2_1
XFILLER_0_196_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24606_ _04409_ _04438_ VGND VGND VPWR VPWR _04461_ sky130_fd_sc_hd__nor2_1
X_12620_ net6664 net6673 net6678 VGND VGND VPWR VPWR _04893_ sky130_fd_sc_hd__nor3b_1
X_21818_ _01825_ _01826_ VGND VGND VPWR VPWR _01827_ sky130_fd_sc_hd__nand2_1
X_22798_ pid_d.kp\[11\] net3068 net2035 VGND VGND VPWR VPWR _02707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25586_ clknet_leaf_90_clk _00459_ net8425 VGND VGND VPWR VPWR cordic0.cos\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8300 net8301 VGND VGND VPWR VPWR net8300 sky130_fd_sc_hd__clkbuf_1
Xwire8311 net18 VGND VGND VPWR VPWR net8311 sky130_fd_sc_hd__clkbuf_1
Xwire8322 net8323 VGND VGND VPWR VPWR net8322 sky130_fd_sc_hd__clkbuf_1
X_24537_ _04314_ _04372_ VGND VGND VPWR VPWR _04393_ sky130_fd_sc_hd__nand2_1
X_21749_ _01757_ _01758_ VGND VGND VPWR VPWR _01759_ sky130_fd_sc_hd__xor2_1
Xwire8333 net8328 VGND VGND VPWR VPWR net8333 sky130_fd_sc_hd__clkbuf_1
Xwire8344 net8345 VGND VGND VPWR VPWR net8344 sky130_fd_sc_hd__buf_1
Xfanout6803 cordic0.vec\[1\]\[16\] VGND VGND VPWR VPWR net6803 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7610 net7605 VGND VGND VPWR VPWR net7610 sky130_fd_sc_hd__buf_1
Xmax_length4042 _09032_ VGND VGND VPWR VPWR net4042 sky130_fd_sc_hd__buf_1
Xwire7621 net7622 VGND VGND VPWR VPWR net7621 sky130_fd_sc_hd__buf_1
X_15270_ _07008_ net1286 net1287 VGND VGND VPWR VPWR _07344_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_0_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8366 net8367 VGND VGND VPWR VPWR net8366 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout6825 net6835 VGND VGND VPWR VPWR net6825 sky130_fd_sc_hd__clkbuf_2
Xwire7632 net7628 VGND VGND VPWR VPWR net7632 sky130_fd_sc_hd__buf_1
X_24468_ _04323_ _04325_ VGND VGND VPWR VPWR _04326_ sky130_fd_sc_hd__xnor2_1
Xwire8377 net8378 VGND VGND VPWR VPWR net8377 sky130_fd_sc_hd__clkbuf_1
Xwire7643 net7644 VGND VGND VPWR VPWR net7643 sky130_fd_sc_hd__buf_1
Xmax_length3330 net3331 VGND VGND VPWR VPWR net3330 sky130_fd_sc_hd__buf_1
Xwire7654 net7655 VGND VGND VPWR VPWR net7654 sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_length3341 net3342 VGND VGND VPWR VPWR net3341 sky130_fd_sc_hd__clkbuf_1
X_14221_ net9157 _05779_ net156 net2373 VGND VGND VPWR VPWR _00030_ sky130_fd_sc_hd__a22o_1
Xfanout6858 net6861 VGND VGND VPWR VPWR net6858 sky130_fd_sc_hd__buf_1
Xwire6920 net6921 VGND VGND VPWR VPWR net6920 sky130_fd_sc_hd__buf_1
Xwire8399 net8400 VGND VGND VPWR VPWR net8399 sky130_fd_sc_hd__buf_1
XFILLER_0_190_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23419_ _03217_ _03218_ _03288_ VGND VGND VPWR VPWR _03289_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_20_Left_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire7676 net7677 VGND VGND VPWR VPWR net7676 sky130_fd_sc_hd__clkbuf_1
X_24399_ net7522 _04191_ net292 net7465 net374 VGND VGND VPWR VPWR _04258_ sky130_fd_sc_hd__a221o_1
Xwire6931 cordic0.vec\[1\]\[10\] VGND VGND VPWR VPWR net6931 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7687 net7690 VGND VGND VPWR VPWR net7687 sky130_fd_sc_hd__buf_1
XFILLER_0_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6942 net6943 VGND VGND VPWR VPWR net6942 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7698 net7699 VGND VGND VPWR VPWR net7698 sky130_fd_sc_hd__buf_1
XFILLER_0_123_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire6953 net6957 VGND VGND VPWR VPWR net6953 sky130_fd_sc_hd__clkbuf_1
Xmax_length2640 _07843_ VGND VGND VPWR VPWR net2640 sky130_fd_sc_hd__buf_1
X_14152_ _06378_ _06380_ VGND VGND VPWR VPWR _06413_ sky130_fd_sc_hd__nor2_1
Xwire6964 net6965 VGND VGND VPWR VPWR net6964 sky130_fd_sc_hd__buf_1
Xwire6975 net6976 VGND VGND VPWR VPWR net6975 sky130_fd_sc_hd__buf_1
XFILLER_0_10_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6986 net6987 VGND VGND VPWR VPWR net6986 sky130_fd_sc_hd__clkbuf_1
Xwire6997 net6993 VGND VGND VPWR VPWR net6997 sky130_fd_sc_hd__buf_1
X_13103_ _05374_ _05375_ VGND VGND VPWR VPWR _05376_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length1961 _04976_ VGND VGND VPWR VPWR net1961 sky130_fd_sc_hd__buf_1
X_14083_ _06340_ _06345_ VGND VGND VPWR VPWR _06346_ sky130_fd_sc_hd__xnor2_1
X_18960_ net6209 _10796_ VGND VGND VPWR VPWR _10797_ sky130_fd_sc_hd__xnor2_4
X_13034_ net1140 net1004 VGND VGND VPWR VPWR _05307_ sky130_fd_sc_hd__or2_1
X_17911_ net3260 _09653_ _09667_ VGND VGND VPWR VPWR _09762_ sky130_fd_sc_hd__and3_1
X_18891_ net9076 net2287 net1450 _10732_ VGND VGND VPWR VPWR _00448_ sky130_fd_sc_hd__a31o_1
X_17842_ net7104 _09643_ _09620_ VGND VGND VPWR VPWR _09693_ sky130_fd_sc_hd__o21a_1
X_17773_ net7133 net7120 VGND VGND VPWR VPWR _09624_ sky130_fd_sc_hd__nor2b_1
X_14985_ net3539 net3541 VGND VGND VPWR VPWR _07059_ sky130_fd_sc_hd__xnor2_1
Xwire1260 _08058_ VGND VGND VPWR VPWR net1260 sky130_fd_sc_hd__dlymetal6s2s_1
X_19512_ net4045 _11348_ VGND VGND VPWR VPWR _11349_ sky130_fd_sc_hd__xnor2_1
Xwire1271 _07610_ VGND VGND VPWR VPWR net1271 sky130_fd_sc_hd__clkbuf_1
X_16724_ _08746_ _08749_ VGND VGND VPWR VPWR _08750_ sky130_fd_sc_hd__xnor2_1
X_13936_ net906 _06201_ VGND VGND VPWR VPWR _06202_ sky130_fd_sc_hd__xor2_1
Xwire1282 _07161_ VGND VGND VPWR VPWR net1282 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1293 net1294 VGND VGND VPWR VPWR net1293 sky130_fd_sc_hd__buf_1
XFILLER_0_92_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19443_ net2507 _11278_ _11279_ VGND VGND VPWR VPWR _11280_ sky130_fd_sc_hd__and3_1
X_16655_ net7316 net1240 net6554 VGND VGND VPWR VPWR _08691_ sky130_fd_sc_hd__mux2_1
X_13867_ _06132_ _06133_ VGND VGND VPWR VPWR _06134_ sky130_fd_sc_hd__xor2_1
X_15606_ _07613_ _07615_ _07677_ VGND VGND VPWR VPWR _07678_ sky130_fd_sc_hd__o21a_1
XFILLER_0_174_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12818_ net7779 net2354 net2316 VGND VGND VPWR VPWR _05091_ sky130_fd_sc_hd__and3_1
X_19374_ _11046_ _11207_ VGND VGND VPWR VPWR _11211_ sky130_fd_sc_hd__nor2_1
X_16586_ _08640_ VGND VGND VPWR VPWR _00234_ sky130_fd_sc_hd__clkbuf_1
X_13798_ _05954_ _05957_ VGND VGND VPWR VPWR _06066_ sky130_fd_sc_hd__nand2_1
XFILLER_0_158_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18325_ _09680_ net3955 VGND VGND VPWR VPWR _10176_ sky130_fd_sc_hd__or2b_1
X_15537_ _07597_ _07609_ VGND VGND VPWR VPWR _07610_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12749_ net4260 _05021_ VGND VGND VPWR VPWR _05022_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18256_ _10105_ _10100_ _10101_ VGND VGND VPWR VPWR _10107_ sky130_fd_sc_hd__nand3_1
XFILLER_0_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15468_ _07504_ _07541_ VGND VGND VPWR VPWR _07542_ sky130_fd_sc_hd__xor2_1
XFILLER_0_115_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17207_ net4036 VGND VGND VPWR VPWR _09157_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14419_ _06618_ VGND VGND VPWR VPWR _00089_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18187_ _10037_ net2554 VGND VGND VPWR VPWR _10038_ sky130_fd_sc_hd__xnor2_4
X_15399_ _07403_ _07404_ _07407_ VGND VGND VPWR VPWR _07473_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17138_ net6906 VGND VGND VPWR VPWR _09092_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire590 net591 VGND VGND VPWR VPWR net590 sky130_fd_sc_hd__buf_1
XFILLER_0_12_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17069_ _09027_ VGND VGND VPWR VPWR _00330_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_6_clk clknet_4_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_176_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20080_ _11904_ _11908_ VGND VGND VPWR VPWR _11909_ sky130_fd_sc_hd__xor2_2
XFILLER_0_176_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_191_Right_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23770_ _03634_ _03635_ VGND VGND VPWR VPWR _03636_ sky130_fd_sc_hd__or2b_1
X_20982_ _00997_ _00943_ VGND VGND VPWR VPWR _00998_ sky130_fd_sc_hd__xnor2_2
X_22721_ net8921 net8102 net90 net93 VGND VGND VPWR VPWR _02657_ sky130_fd_sc_hd__or4_1
XFILLER_0_189_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6928 net6929 VGND VGND VPWR VPWR net6928 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25440_ clknet_leaf_91_clk _00323_ net8432 VGND VGND VPWR VPWR matmul0.sin\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_22652_ _02553_ _02578_ net3081 VGND VGND VPWR VPWR _02611_ sky130_fd_sc_hd__a21o_1
XFILLER_0_165_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21603_ _01605_ _01614_ VGND VGND VPWR VPWR _01615_ sky130_fd_sc_hd__xnor2_2
X_22583_ net8891 _02562_ VGND VGND VPWR VPWR _02563_ sky130_fd_sc_hd__and2_1
X_25371_ clknet_leaf_57_clk _00254_ net8711 VGND VGND VPWR VPWR matmul0.alpha_pass\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24322_ _04180_ _04181_ VGND VGND VPWR VPWR _04182_ sky130_fd_sc_hd__nand2_1
X_21534_ net860 net806 _01545_ VGND VGND VPWR VPWR _01546_ sky130_fd_sc_hd__o21a_1
Xfanout5409 net5422 VGND VGND VPWR VPWR net5409 sky130_fd_sc_hd__buf_1
Xwire6205 net6204 VGND VGND VPWR VPWR net6205 sky130_fd_sc_hd__buf_1
XFILLER_0_8_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24253_ _04111_ _04112_ VGND VGND VPWR VPWR _04114_ sky130_fd_sc_hd__or2_1
Xwire6216 net6217 VGND VGND VPWR VPWR net6216 sky130_fd_sc_hd__buf_1
XFILLER_0_172_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21465_ net1726 _01476_ VGND VGND VPWR VPWR _01478_ sky130_fd_sc_hd__nand2_1
Xwire6227 net6223 VGND VGND VPWR VPWR net6227 sky130_fd_sc_hd__buf_1
XFILLER_0_133_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6238 net6233 VGND VGND VPWR VPWR net6238 sky130_fd_sc_hd__buf_1
Xwire5504 net5496 VGND VGND VPWR VPWR net5504 sky130_fd_sc_hd__clkbuf_1
X_23204_ net5111 net5083 VGND VGND VPWR VPWR _03074_ sky130_fd_sc_hd__and2_1
Xwire6249 net6247 VGND VGND VPWR VPWR net6249 sky130_fd_sc_hd__buf_1
Xwire5515 net5516 VGND VGND VPWR VPWR net5515 sky130_fd_sc_hd__buf_1
X_20416_ net1915 _12211_ VGND VGND VPWR VPWR _12213_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24184_ _03941_ _03960_ _04043_ _04044_ VGND VGND VPWR VPWR _04045_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5537 net5538 VGND VGND VPWR VPWR net5537 sky130_fd_sc_hd__buf_1
X_21396_ _01398_ _01409_ VGND VGND VPWR VPWR _01410_ sky130_fd_sc_hd__xnor2_1
Xwire4803 net4804 VGND VGND VPWR VPWR net4803 sky130_fd_sc_hd__buf_1
Xwire5559 net5562 VGND VGND VPWR VPWR net5559 sky130_fd_sc_hd__buf_1
X_23135_ _02990_ _03002_ net1676 VGND VGND VPWR VPWR _03005_ sky130_fd_sc_hd__o21a_1
Xwire4825 net4821 VGND VGND VPWR VPWR net4825 sky130_fd_sc_hd__buf_1
X_20347_ _12126_ _12137_ _12138_ cordic0.slte0.opA\[4\] VGND VGND VPWR VPWR _12149_
+ sky130_fd_sc_hd__a31o_1
Xwire4836 net4837 VGND VGND VPWR VPWR net4836 sky130_fd_sc_hd__buf_1
XFILLER_0_102_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4858 net4849 VGND VGND VPWR VPWR net4858 sky130_fd_sc_hd__clkbuf_1
Xwire4869 net4870 VGND VGND VPWR VPWR net4869 sky130_fd_sc_hd__clkbuf_1
X_23066_ _02934_ _02935_ VGND VGND VPWR VPWR _02936_ sky130_fd_sc_hd__xnor2_1
X_20278_ net6516 _12084_ VGND VGND VPWR VPWR _12085_ sky130_fd_sc_hd__or2_1
X_22017_ _01928_ _01930_ _02023_ VGND VGND VPWR VPWR _02024_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_41_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14770_ net8954 net2867 _06897_ VGND VGND VPWR VPWR _00161_ sky130_fd_sc_hd__a21bo_1
X_23968_ net4811 _03711_ _03830_ VGND VGND VPWR VPWR _03832_ sky130_fd_sc_hd__a21o_1
X_13721_ net780 _05989_ VGND VGND VPWR VPWR _05990_ sky130_fd_sc_hd__xnor2_2
Xmax_length8875 net8876 VGND VGND VPWR VPWR net8875 sky130_fd_sc_hd__clkbuf_1
X_25707_ clknet_leaf_6_clk _00580_ net8561 VGND VGND VPWR VPWR pid_d.mult0.b\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22919_ _02270_ _02802_ net5340 VGND VGND VPWR VPWR _02810_ sky130_fd_sc_hd__o21ba_1
X_23899_ _03762_ _03664_ _03763_ VGND VGND VPWR VPWR _03764_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16440_ _08466_ _08474_ _08500_ VGND VGND VPWR VPWR _08501_ sky130_fd_sc_hd__o21ai_1
X_13652_ net7832 net1328 _05794_ VGND VGND VPWR VPWR _05922_ sky130_fd_sc_hd__a21o_1
X_25638_ clknet_leaf_103_clk _00511_ net8375 VGND VGND VPWR VPWR cordic0.vec\[0\]\[10\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_195_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12603_ _04880_ VGND VGND VPWR VPWR _00009_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout8046 net8065 VGND VGND VPWR VPWR net8046 sky130_fd_sc_hd__clkbuf_1
X_16371_ _08433_ VGND VGND VPWR VPWR _00226_ sky130_fd_sc_hd__clkbuf_1
X_13583_ net504 _05773_ VGND VGND VPWR VPWR _05854_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25569_ clknet_leaf_99_clk _00442_ net8387 VGND VGND VPWR VPWR cordic0.sin\[3\] sky130_fd_sc_hd__dfrtp_1
X_18110_ _09875_ _09881_ _09894_ net2551 VGND VGND VPWR VPWR _09961_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_66_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8130 net8131 VGND VGND VPWR VPWR net8130 sky130_fd_sc_hd__clkbuf_1
Xwire8141 net8142 VGND VGND VPWR VPWR net8141 sky130_fd_sc_hd__clkbuf_1
X_15322_ _07024_ _07031_ _07395_ VGND VGND VPWR VPWR _07396_ sky130_fd_sc_hd__o21a_1
XFILLER_0_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19090_ _10827_ net6318 net3898 VGND VGND VPWR VPWR _10927_ sky130_fd_sc_hd__a21o_1
Xwire8152 net8153 VGND VGND VPWR VPWR net8152 sky130_fd_sc_hd__clkbuf_1
Xwire8163 net8164 VGND VGND VPWR VPWR net8163 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout6622 matmul0.matmul_stage_inst.state\[2\] VGND VGND VPWR VPWR net6622 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_136_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8174 net8175 VGND VGND VPWR VPWR net8174 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8185 net37 VGND VGND VPWR VPWR net8185 sky130_fd_sc_hd__clkbuf_1
X_18041_ net3963 _09843_ VGND VGND VPWR VPWR _09892_ sky130_fd_sc_hd__xnor2_2
Xwire8196 net8197 VGND VGND VPWR VPWR net8196 sky130_fd_sc_hd__clkbuf_1
X_15253_ net1878 net1275 VGND VGND VPWR VPWR _07327_ sky130_fd_sc_hd__nand2_1
Xwire7473 net7474 VGND VGND VPWR VPWR net7473 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout6677 net6679 VGND VGND VPWR VPWR net6677 sky130_fd_sc_hd__clkbuf_2
X_14204_ _06438_ _06459_ _06460_ VGND VGND VPWR VPWR _06463_ sky130_fd_sc_hd__o21ai_1
Xwire7484 net7485 VGND VGND VPWR VPWR net7484 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7495 pid_q.state\[3\] VGND VGND VPWR VPWR net7495 sky130_fd_sc_hd__clkbuf_1
Xwire6750 net6751 VGND VGND VPWR VPWR net6750 sky130_fd_sc_hd__buf_1
XFILLER_0_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15184_ net1277 _07183_ VGND VGND VPWR VPWR _07258_ sky130_fd_sc_hd__xor2_1
Xwire6761 net6764 VGND VGND VPWR VPWR net6761 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6783 net6782 VGND VGND VPWR VPWR net6783 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14135_ _06369_ _06396_ VGND VGND VPWR VPWR _06397_ sky130_fd_sc_hd__xor2_1
Xwire6794 net6792 VGND VGND VPWR VPWR net6794 sky130_fd_sc_hd__buf_1
X_19992_ _11819_ _11821_ VGND VGND VPWR VPWR _11823_ sky130_fd_sc_hd__and2_1
X_14066_ _06327_ _06328_ VGND VGND VPWR VPWR _06329_ sky130_fd_sc_hd__and2_1
X_18943_ net6375 net207 _10772_ VGND VGND VPWR VPWR _10782_ sky130_fd_sc_hd__and3_1
X_13017_ _05289_ VGND VGND VPWR VPWR _05290_ sky130_fd_sc_hd__clkbuf_2
X_18874_ net6860 _10715_ VGND VGND VPWR VPWR _10716_ sky130_fd_sc_hd__xnor2_2
X_17825_ net6926 net6875 VGND VGND VPWR VPWR _09676_ sky130_fd_sc_hd__xor2_2
Xhold1 matmul0.matmul_stage_inst.c\[9\] VGND VGND VPWR VPWR net8954 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_146_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17756_ net6963 net6925 VGND VGND VPWR VPWR _09607_ sky130_fd_sc_hd__xnor2_1
X_14968_ net4136 net4129 VGND VGND VPWR VPWR _07042_ sky130_fd_sc_hd__nor2_1
XFILLER_0_178_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1090 _08202_ VGND VGND VPWR VPWR net1090 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16707_ _08734_ net383 matmul0.matmul_stage_inst.mult2\[12\] VGND VGND VPWR VPWR
+ _08735_ sky130_fd_sc_hd__o21ba_1
X_13919_ net7681 _05873_ VGND VGND VPWR VPWR _06185_ sky130_fd_sc_hd__nand2_1
XFILLER_0_159_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17687_ net3272 svm0.tA\[11\] _09566_ VGND VGND VPWR VPWR _09567_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14899_ net4213 net4211 net4210 net4208 VGND VGND VPWR VPWR _06973_ sky130_fd_sc_hd__o22a_1
XFILLER_0_71_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19426_ net6241 net6346 VGND VGND VPWR VPWR _11263_ sky130_fd_sc_hd__and2b_1
XFILLER_0_147_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16638_ matmul0.matmul_stage_inst.mult2\[3\] matmul0.matmul_stage_inst.mult1\[3\]
+ VGND VGND VPWR VPWR _08676_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19357_ net6202 net2515 net2508 _11193_ VGND VGND VPWR VPWR _11194_ sky130_fd_sc_hd__a31o_1
X_16569_ _08582_ _08585_ VGND VGND VPWR VPWR _08628_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18308_ _09675_ _10108_ _08967_ net7040 VGND VGND VPWR VPWR _10159_ sky130_fd_sc_hd__a211o_1
XFILLER_0_73_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19288_ net3909 net3209 VGND VGND VPWR VPWR _11125_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18239_ _10087_ _10088_ _10089_ net7095 net3340 VGND VGND VPWR VPWR _10090_ sky130_fd_sc_hd__a221o_1
XFILLER_0_154_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21250_ net5426 net5922 VGND VGND VPWR VPWR _01265_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20201_ _12010_ _12025_ VGND VGND VPWR VPWR _12026_ sky130_fd_sc_hd__xnor2_1
X_21181_ _01188_ _01196_ VGND VGND VPWR VPWR _01197_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_187_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3409 net3410 VGND VGND VPWR VPWR net3409 sky130_fd_sc_hd__buf_1
XFILLER_0_187_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20132_ _11959_ _11915_ _11913_ VGND VGND VPWR VPWR _11960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2708 net2709 VGND VGND VPWR VPWR net2708 sky130_fd_sc_hd__buf_1
XFILLER_0_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2719 net2720 VGND VGND VPWR VPWR net2719 sky130_fd_sc_hd__buf_1
X_24940_ pid_q.ki\[9\] _04720_ net1360 VGND VGND VPWR VPWR _04721_ sky130_fd_sc_hd__mux2_1
X_20063_ _11889_ _11891_ VGND VGND VPWR VPWR _11892_ sky130_fd_sc_hd__xor2_1
X_24871_ net4481 net2397 net3009 net4478 VGND VGND VPWR VPWR _04672_ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23822_ _03600_ _03602_ VGND VGND VPWR VPWR _03687_ sky130_fd_sc_hd__nor2_1
XFILLER_0_174_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23753_ _03617_ _03618_ VGND VGND VPWR VPWR _03619_ sky130_fd_sc_hd__xnor2_1
X_20965_ net5506 net5950 VGND VGND VPWR VPWR _00981_ sky130_fd_sc_hd__nand2_1
Xmax_length7459 net7460 VGND VGND VPWR VPWR net7459 sky130_fd_sc_hd__buf_1
X_22704_ _02644_ VGND VGND VPWR VPWR _00594_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23684_ _03548_ _03550_ VGND VGND VPWR VPWR _03551_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20896_ _00895_ _00911_ VGND VGND VPWR VPWR _00912_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25423_ clknet_leaf_90_clk _00306_ net8424 VGND VGND VPWR VPWR matmul0.cos\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_192_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22635_ net3090 _02549_ net3080 VGND VGND VPWR VPWR _02602_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22566_ net7368 net7353 VGND VGND VPWR VPWR _02549_ sky130_fd_sc_hd__xor2_1
X_25354_ clknet_leaf_84_clk _00237_ net8506 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult2\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24305_ _04162_ _04164_ VGND VGND VPWR VPWR _04165_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21517_ _01528_ _01529_ _01342_ VGND VGND VPWR VPWR _01530_ sky130_fd_sc_hd__o21ba_1
Xwire6013 net6011 VGND VGND VPWR VPWR net6013 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_161_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22497_ _02471_ _02497_ VGND VGND VPWR VPWR _02498_ sky130_fd_sc_hd__xnor2_1
X_25285_ clknet_leaf_89_clk _00168_ net8421 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.d\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire5301 net5302 VGND VGND VPWR VPWR net5301 sky130_fd_sc_hd__clkbuf_1
Xwire6046 net6044 VGND VGND VPWR VPWR net6046 sky130_fd_sc_hd__buf_1
XFILLER_0_181_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24236_ net793 _04096_ VGND VGND VPWR VPWR _04097_ sky130_fd_sc_hd__xnor2_1
X_21448_ _01452_ _01460_ VGND VGND VPWR VPWR _01461_ sky130_fd_sc_hd__xnor2_1
Xwire5312 net5313 VGND VGND VPWR VPWR net5312 sky130_fd_sc_hd__buf_1
Xwire5323 net5324 VGND VGND VPWR VPWR net5323 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5334 net5335 VGND VGND VPWR VPWR net5334 sky130_fd_sc_hd__clkbuf_1
Xwire6079 net6077 VGND VGND VPWR VPWR net6079 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4600 net4601 VGND VGND VPWR VPWR net4600 sky130_fd_sc_hd__clkbuf_1
Xwire5345 pid_d.out\[11\] VGND VGND VPWR VPWR net5345 sky130_fd_sc_hd__clkbuf_1
Xwire4611 net4612 VGND VGND VPWR VPWR net4611 sky130_fd_sc_hd__clkbuf_1
X_24167_ pid_q.curr_error\[7\] VGND VGND VPWR VPWR _04029_ sky130_fd_sc_hd__inv_2
Xwire5356 pid_d.out\[8\] VGND VGND VPWR VPWR net5356 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5367 net5368 VGND VGND VPWR VPWR net5367 sky130_fd_sc_hd__clkbuf_1
X_21379_ _01288_ _01289_ _01298_ VGND VGND VPWR VPWR _01393_ sky130_fd_sc_hd__a21o_1
Xwire4633 net4634 VGND VGND VPWR VPWR net4633 sky130_fd_sc_hd__buf_1
Xwire5378 net5379 VGND VGND VPWR VPWR net5378 sky130_fd_sc_hd__buf_1
Xwire4644 net4645 VGND VGND VPWR VPWR net4644 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5389 net5390 VGND VGND VPWR VPWR net5389 sky130_fd_sc_hd__buf_1
Xwire3910 net3911 VGND VGND VPWR VPWR net3910 sky130_fd_sc_hd__buf_1
Xwire4655 net4646 VGND VGND VPWR VPWR net4655 sky130_fd_sc_hd__buf_1
X_23118_ net1031 _02987_ _02984_ VGND VGND VPWR VPWR _02988_ sky130_fd_sc_hd__a21o_1
Xwire4666 net4667 VGND VGND VPWR VPWR net4666 sky130_fd_sc_hd__buf_1
X_24098_ net376 _03942_ VGND VGND VPWR VPWR _03960_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4677 net4678 VGND VGND VPWR VPWR net4677 sky130_fd_sc_hd__buf_1
Xwire3932 _10103_ VGND VGND VPWR VPWR net3932 sky130_fd_sc_hd__buf_1
Xwire4688 net4689 VGND VGND VPWR VPWR net4688 sky130_fd_sc_hd__buf_1
Xwire3943 net3944 VGND VGND VPWR VPWR net3943 sky130_fd_sc_hd__clkbuf_1
Xwire4699 net4700 VGND VGND VPWR VPWR net4699 sky130_fd_sc_hd__clkbuf_1
Xwire3954 net3955 VGND VGND VPWR VPWR net3954 sky130_fd_sc_hd__clkbuf_1
X_23049_ _02913_ _02915_ _02918_ VGND VGND VPWR VPWR _02919_ sky130_fd_sc_hd__a21oi_1
X_15940_ _08007_ _08008_ VGND VGND VPWR VPWR _08009_ sky130_fd_sc_hd__or2_1
Xwire3965 _09735_ VGND VGND VPWR VPWR net3965 sky130_fd_sc_hd__clkbuf_1
Xwire3976 _09679_ VGND VGND VPWR VPWR net3976 sky130_fd_sc_hd__buf_1
Xwire3987 _09660_ VGND VGND VPWR VPWR net3987 sky130_fd_sc_hd__buf_1
Xwire3998 _09604_ VGND VGND VPWR VPWR net3998 sky130_fd_sc_hd__buf_1
X_15871_ _07935_ _07939_ VGND VGND VPWR VPWR _07940_ sky130_fd_sc_hd__xnor2_1
X_17610_ net6701 svm0.tB\[12\] VGND VGND VPWR VPWR _09491_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_192_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14822_ _06927_ VGND VGND VPWR VPWR _00183_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18590_ net6786 _10437_ VGND VGND VPWR VPWR _10438_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17541_ svm0.tC\[14\] net6687 VGND VGND VPWR VPWR _09423_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_103_Left_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14753_ net7448 _06883_ _06884_ net7454 net3621 VGND VGND VPWR VPWR _06885_ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13704_ net4248 net1961 VGND VGND VPWR VPWR _05973_ sky130_fd_sc_hd__nor2_1
X_17472_ net4020 _09364_ VGND VGND VPWR VPWR _09365_ sky130_fd_sc_hd__nor2_1
X_14684_ net7454 _06832_ VGND VGND VPWR VPWR _06833_ sky130_fd_sc_hd__nand2_1
X_19211_ _11046_ _11047_ VGND VGND VPWR VPWR _11048_ sky130_fd_sc_hd__nor2_2
XFILLER_0_6_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16423_ net571 _08427_ _08484_ net490 VGND VGND VPWR VPWR _08485_ sky130_fd_sc_hd__o22a_1
XFILLER_0_168_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13635_ _05902_ _05904_ VGND VGND VPWR VPWR _05905_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19142_ net3908 net3906 VGND VGND VPWR VPWR _10979_ sky130_fd_sc_hd__or2_1
Xfanout7131 net7137 VGND VGND VPWR VPWR net7131 sky130_fd_sc_hd__clkbuf_1
X_16354_ net2651 net3587 net3431 net1848 VGND VGND VPWR VPWR _08417_ sky130_fd_sc_hd__and4_1
X_13566_ net7865 net1577 _05710_ VGND VGND VPWR VPWR _05837_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15305_ net2233 _07378_ net3598 _06978_ VGND VGND VPWR VPWR _07379_ sky130_fd_sc_hd__a31o_1
XFILLER_0_81_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19073_ net2527 _10855_ VGND VGND VPWR VPWR _10910_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16285_ net1253 _08346_ _08340_ VGND VGND VPWR VPWR _08349_ sky130_fd_sc_hd__nor3_1
X_13497_ net785 net578 VGND VGND VPWR VPWR _05770_ sky130_fd_sc_hd__and2b_1
Xfanout6452 state\[0\] VGND VGND VPWR VPWR net6452 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout6463 cordic0.gm0.iter\[4\] VGND VGND VPWR VPWR net6463 sky130_fd_sc_hd__buf_1
Xwire7270 net7271 VGND VGND VPWR VPWR net7270 sky130_fd_sc_hd__buf_1
X_18024_ net2549 _09874_ VGND VGND VPWR VPWR _09875_ sky130_fd_sc_hd__xnor2_2
X_15236_ net2705 net2779 VGND VGND VPWR VPWR _07310_ sky130_fd_sc_hd__nor2_1
Xwire7281 matmul0.alpha_pass\[8\] VGND VGND VPWR VPWR net7281 sky130_fd_sc_hd__buf_1
Xwire7292 net7293 VGND VGND VPWR VPWR net7292 sky130_fd_sc_hd__clkbuf_1
Xfanout5751 pid_d.mult0.b\[10\] VGND VGND VPWR VPWR net5751 sky130_fd_sc_hd__buf_1
XFILLER_0_23_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout5762 net5765 VGND VGND VPWR VPWR net5762 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_50_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15167_ _07194_ VGND VGND VPWR VPWR _07241_ sky130_fd_sc_hd__clkbuf_1
Xfanout5795 net5803 VGND VGND VPWR VPWR net5795 sky130_fd_sc_hd__buf_1
XFILLER_0_23_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14118_ net7627 _05348_ VGND VGND VPWR VPWR _06380_ sky130_fd_sc_hd__nand2_1
Xwire5890 net5894 VGND VGND VPWR VPWR net5890 sky130_fd_sc_hd__buf_1
XFILLER_0_120_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19975_ net5999 net2092 VGND VGND VPWR VPWR _11806_ sky130_fd_sc_hd__nand2_1
X_15098_ net3511 net3506 _07026_ _07028_ VGND VGND VPWR VPWR _07172_ sky130_fd_sc_hd__o22a_1
XFILLER_0_66_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14049_ net7742 net1570 _06253_ VGND VGND VPWR VPWR _06313_ sky130_fd_sc_hd__and3_1
X_18926_ _10764_ _10765_ VGND VGND VPWR VPWR _10766_ sky130_fd_sc_hd__xor2_1
XFILLER_0_157_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18857_ net658 _10664_ VGND VGND VPWR VPWR _10699_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17808_ _09640_ _09653_ net1781 VGND VGND VPWR VPWR _09659_ sky130_fd_sc_hd__o21a_1
X_18788_ net6862 net3967 _10579_ _10631_ VGND VGND VPWR VPWR _10632_ sky130_fd_sc_hd__o31a_1
XFILLER_0_55_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17739_ _06530_ _06646_ _09593_ VGND VGND VPWR VPWR _00435_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_173_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20750_ net5558 net5836 VGND VGND VPWR VPWR _12521_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19409_ _11094_ _11045_ VGND VGND VPWR VPWR _11246_ sky130_fd_sc_hd__nand2_1
X_20681_ _12435_ _12446_ _12455_ _12456_ VGND VGND VPWR VPWR _12457_ sky130_fd_sc_hd__o31a_1
XFILLER_0_169_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22420_ net5412 net5676 VGND VGND VPWR VPWR _02422_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3907 _10801_ VGND VGND VPWR VPWR net3907 sky130_fd_sc_hd__buf_1
XFILLER_0_61_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22351_ net5694 net5411 VGND VGND VPWR VPWR _02354_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21302_ net5487 VGND VGND VPWR VPWR _01317_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25070_ net3734 _04811_ _04816_ VGND VGND VPWR VPWR _04817_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22282_ net5722 net5388 VGND VGND VPWR VPWR _02286_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24021_ _03878_ _03883_ VGND VGND VPWR VPWR _03884_ sky130_fd_sc_hd__xnor2_1
Xhold220 pid_q.out\[8\] VGND VGND VPWR VPWR net9173 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21233_ net5985 pid_d.prev_int\[1\] VGND VGND VPWR VPWR _01248_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold231 pid_q.prev_error\[11\] VGND VGND VPWR VPWR net9184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 pid_d.curr_int\[15\] VGND VGND VPWR VPWR net9195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 pid_d.curr_int\[0\] VGND VGND VPWR VPWR net9206 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3206 _10836_ VGND VGND VPWR VPWR net3206 sky130_fd_sc_hd__buf_1
Xhold264 pid_d.prev_int\[8\] VGND VGND VPWR VPWR net9217 sky130_fd_sc_hd__dlygate4sd3_1
X_21164_ _01176_ _01179_ VGND VGND VPWR VPWR _01180_ sky130_fd_sc_hd__nor2_1
Xwire3217 net3218 VGND VGND VPWR VPWR net3217 sky130_fd_sc_hd__clkbuf_1
Xhold275 pid_q.prev_error\[1\] VGND VGND VPWR VPWR net9228 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3228 _10124_ VGND VGND VPWR VPWR net3228 sky130_fd_sc_hd__buf_1
Xhold286 pid_q.prev_int\[4\] VGND VGND VPWR VPWR net9239 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3239 _09801_ VGND VGND VPWR VPWR net3239 sky130_fd_sc_hd__buf_1
Xwire2505 _11446_ VGND VGND VPWR VPWR net2505 sky130_fd_sc_hd__buf_1
X_20115_ _11292_ _11942_ net6027 VGND VGND VPWR VPWR _11943_ sky130_fd_sc_hd__mux2_1
Xwire2516 net2517 VGND VGND VPWR VPWR net2516 sky130_fd_sc_hd__buf_1
X_21095_ _01103_ _01102_ _01100_ net5793 net5642 VGND VGND VPWR VPWR _01111_ sky130_fd_sc_hd__o2111ai_2
Xwire2527 _10852_ VGND VGND VPWR VPWR net2527 sky130_fd_sc_hd__buf_1
Xwire2538 _10486_ VGND VGND VPWR VPWR net2538 sky130_fd_sc_hd__clkbuf_1
Xwire1804 net1805 VGND VGND VPWR VPWR net1804 sky130_fd_sc_hd__clkbuf_2
Xwire2549 _09869_ VGND VGND VPWR VPWR net2549 sky130_fd_sc_hd__clkbuf_2
Xwire1815 _08915_ VGND VGND VPWR VPWR net1815 sky130_fd_sc_hd__buf_1
X_24923_ _04709_ VGND VGND VPWR VPWR _00748_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20046_ _11840_ _11875_ VGND VGND VPWR VPWR _11876_ sky130_fd_sc_hd__xnor2_1
Xwire1826 net1827 VGND VGND VPWR VPWR net1826 sky130_fd_sc_hd__buf_1
Xwire1837 _08819_ VGND VGND VPWR VPWR net1837 sky130_fd_sc_hd__buf_1
Xwire1859 _07578_ VGND VGND VPWR VPWR net1859 sky130_fd_sc_hd__buf_1
X_24854_ pid_q.ki\[0\] net3022 net3007 pid_q.kp\[0\] VGND VGND VPWR VPWR _04660_ sky130_fd_sc_hd__a22o_1
Xmax_length7201 net7202 VGND VGND VPWR VPWR net7201 sky130_fd_sc_hd__clkbuf_1
X_23805_ pid_q.prev_int\[4\] VGND VGND VPWR VPWR _03670_ sky130_fd_sc_hd__inv_2
X_24785_ pid_q.curr_error\[11\] net1643 _04543_ net455 VGND VGND VPWR VPWR _00708_
+ sky130_fd_sc_hd__a22o_1
Xmax_length7245 net7246 VGND VGND VPWR VPWR net7245 sky130_fd_sc_hd__clkbuf_1
X_21997_ _02004_ VGND VGND VPWR VPWR _02005_ sky130_fd_sc_hd__inv_2
XFILLER_0_178_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23736_ net4543 net5031 VGND VGND VPWR VPWR _03602_ sky130_fd_sc_hd__nand2_1
Xmax_length6522 net6523 VGND VGND VPWR VPWR net6522 sky130_fd_sc_hd__buf_1
X_20948_ _00896_ _00898_ net5905 VGND VGND VPWR VPWR _00964_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23667_ _03400_ _03401_ _03533_ VGND VGND VPWR VPWR _03534_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_48_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20879_ _12530_ _00894_ VGND VGND VPWR VPWR _00895_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13420_ net7921 net1929 _05692_ VGND VGND VPWR VPWR _05693_ sky130_fd_sc_hd__and3_1
X_25406_ clknet_leaf_76_clk _00289_ net8472 VGND VGND VPWR VPWR matmul0.a\[9\] sky130_fd_sc_hd__dfrtp_1
X_22618_ _02589_ VGND VGND VPWR VPWR _00563_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23598_ _03371_ _03374_ VGND VGND VPWR VPWR _03466_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length5887 net5883 VGND VGND VPWR VPWR net5887 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13351_ _05621_ _05622_ _05613_ _05614_ VGND VGND VPWR VPWR _05624_ sky130_fd_sc_hd__a211o_1
X_25337_ clknet_leaf_83_clk _00220_ net8507 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22549_ pid_d.curr_error\[12\] net3017 net2460 VGND VGND VPWR VPWR _02537_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5036 net5047 VGND VGND VPWR VPWR net5036 sky130_fd_sc_hd__buf_1
X_16070_ _08131_ _08136_ VGND VGND VPWR VPWR _08137_ sky130_fd_sc_hd__xor2_1
X_13282_ _05527_ VGND VGND VPWR VPWR _05555_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25268_ clknet_leaf_77_clk _00151_ net8437 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.b\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire5120 net5121 VGND VGND VPWR VPWR net5120 sky130_fd_sc_hd__buf_1
Xfanout4324 pid_d.state\[4\] VGND VGND VPWR VPWR net4324 sky130_fd_sc_hd__buf_1
Xwire5131 net5132 VGND VGND VPWR VPWR net5131 sky130_fd_sc_hd__clkbuf_1
X_15021_ net4178 VGND VGND VPWR VPWR _07095_ sky130_fd_sc_hd__buf_1
Xwire5142 net5145 VGND VGND VPWR VPWR net5142 sky130_fd_sc_hd__buf_1
X_24219_ net4937 net4501 VGND VGND VPWR VPWR _04080_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5153 net5154 VGND VGND VPWR VPWR net5153 sky130_fd_sc_hd__clkbuf_1
X_25199_ clknet_leaf_62_clk _00088_ net8666 VGND VGND VPWR VPWR matmul0.b_in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout4368 net4376 VGND VGND VPWR VPWR net4368 sky130_fd_sc_hd__buf_1
Xwire5175 pid_q.curr_int\[12\] VGND VGND VPWR VPWR net5175 sky130_fd_sc_hd__clkbuf_2
Xfanout4379 net4388 VGND VGND VPWR VPWR net4379 sky130_fd_sc_hd__buf_1
Xwire5186 net5187 VGND VGND VPWR VPWR net5186 sky130_fd_sc_hd__clkbuf_1
Xwire4441 net4442 VGND VGND VPWR VPWR net4441 sky130_fd_sc_hd__clkbuf_1
Xwire4452 net4453 VGND VGND VPWR VPWR net4452 sky130_fd_sc_hd__clkbuf_1
Xwire4463 net4464 VGND VGND VPWR VPWR net4463 sky130_fd_sc_hd__clkbuf_1
Xwire4485 net4482 VGND VGND VPWR VPWR net4485 sky130_fd_sc_hd__buf_1
Xwire3740 _03771_ VGND VGND VPWR VPWR net3740 sky130_fd_sc_hd__clkbuf_1
Xwire4496 net4497 VGND VGND VPWR VPWR net4496 sky130_fd_sc_hd__buf_1
Xwire3751 net3752 VGND VGND VPWR VPWR net3751 sky130_fd_sc_hd__clkbuf_1
X_16972_ net2606 _08934_ VGND VGND VPWR VPWR _08935_ sky130_fd_sc_hd__xnor2_1
X_19760_ _11517_ _11524_ net1415 VGND VGND VPWR VPWR _11595_ sky130_fd_sc_hd__a21o_1
Xwire3762 _02716_ VGND VGND VPWR VPWR net3762 sky130_fd_sc_hd__buf_1
Xwire3773 _02545_ VGND VGND VPWR VPWR net3773 sky130_fd_sc_hd__clkbuf_1
Xwire3784 _01863_ VGND VGND VPWR VPWR net3784 sky130_fd_sc_hd__clkbuf_1
X_15923_ net2836 net2829 net2846 net1846 VGND VGND VPWR VPWR _07992_ sky130_fd_sc_hd__and4_1
X_18711_ _10464_ _10555_ _10556_ VGND VGND VPWR VPWR _10557_ sky130_fd_sc_hd__o21ai_1
X_19691_ _11458_ net2101 net1749 VGND VGND VPWR VPWR _11527_ sky130_fd_sc_hd__o21a_1
X_18642_ _10488_ VGND VGND VPWR VPWR _10489_ sky130_fd_sc_hd__inv_2
X_15854_ _07923_ VGND VGND VPWR VPWR _00219_ sky130_fd_sc_hd__clkbuf_1
X_14805_ net9002 net2871 _06919_ VGND VGND VPWR VPWR _00174_ sky130_fd_sc_hd__a21o_1
X_18573_ _10171_ net3960 _10364_ VGND VGND VPWR VPWR _10421_ sky130_fd_sc_hd__mux2_1
X_15785_ _07852_ _07854_ VGND VGND VPWR VPWR _07855_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12997_ net7803 net1619 _05178_ _05179_ VGND VGND VPWR VPWR _05270_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17524_ net6694 _09407_ _09408_ _09406_ VGND VGND VPWR VPWR _00404_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14736_ net7455 _06827_ VGND VGND VPWR VPWR _06871_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17455_ svm0.delta\[3\] _09349_ VGND VGND VPWR VPWR _09350_ sky130_fd_sc_hd__xnor2_1
X_14667_ net9024 net2872 _06819_ VGND VGND VPWR VPWR _00136_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16406_ net2625 net2623 net2213 VGND VGND VPWR VPWR _08468_ sky130_fd_sc_hd__or3_1
X_13618_ _05878_ _05887_ VGND VGND VPWR VPWR _05888_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17386_ _09291_ net614 _09292_ _09294_ VGND VGND VPWR VPWR _00380_ sky130_fd_sc_hd__a31o_1
X_14598_ _06770_ _06771_ net2882 VGND VGND VPWR VPWR _06772_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19125_ net6069 _10961_ VGND VGND VPWR VPWR _10962_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16337_ _08393_ _08398_ VGND VGND VPWR VPWR _08400_ sky130_fd_sc_hd__or2_1
X_13549_ _05818_ _05819_ VGND VGND VPWR VPWR _05820_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19056_ _10891_ _10892_ VGND VGND VPWR VPWR _10893_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16268_ _08325_ net1249 VGND VGND VPWR VPWR _08332_ sky130_fd_sc_hd__xnor2_1
X_18007_ net6990 net7035 VGND VGND VPWR VPWR _09858_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_51_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15219_ net1883 _07250_ VGND VGND VPWR VPWR _07293_ sky130_fd_sc_hd__xor2_1
XFILLER_0_112_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16199_ _08170_ _08172_ _08263_ net2815 VGND VGND VPWR VPWR _08264_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_168_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19958_ _11755_ net3199 _11758_ VGND VGND VPWR VPWR _11789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18909_ _10748_ _10749_ net1443 VGND VGND VPWR VPWR _10750_ sky130_fd_sc_hd__a21oi_1
X_19889_ _11667_ net708 VGND VGND VPWR VPWR _11722_ sky130_fd_sc_hd__or2_1
X_21920_ _00977_ net5649 VGND VGND VPWR VPWR _01928_ sky130_fd_sc_hd__nand2_1
XFILLER_0_184_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21851_ net2475 _01787_ _01859_ VGND VGND VPWR VPWR _01860_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20802_ _12536_ _12547_ _00815_ _00817_ VGND VGND VPWR VPWR _00818_ sky130_fd_sc_hd__o211a_1
X_24570_ net4843 net4487 VGND VGND VPWR VPWR _04426_ sky130_fd_sc_hd__nand2_1
X_21782_ _01780_ _01791_ VGND VGND VPWR VPWR _01792_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23521_ pid_q.curr_int\[1\] net3061 net2028 _03389_ VGND VGND VPWR VPWR _00666_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20733_ net5509 net5867 VGND VGND VPWR VPWR _12504_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8707 net8702 VGND VGND VPWR VPWR net8707 sky130_fd_sc_hd__buf_1
XFILLER_0_18_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8718 net8719 VGND VGND VPWR VPWR net8718 sky130_fd_sc_hd__buf_1
XFILLER_0_92_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8729 net8727 VGND VGND VPWR VPWR net8729 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_133_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23452_ _03282_ _03293_ _03320_ VGND VGND VPWR VPWR _03321_ sky130_fd_sc_hd__a21o_1
X_20664_ net4039 net6757 _12440_ VGND VGND VPWR VPWR _12441_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_190_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire408 net409 VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__buf_1
XFILLER_0_80_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22403_ _02403_ _02404_ VGND VGND VPWR VPWR _02405_ sky130_fd_sc_hd__or2b_1
XFILLER_0_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire419 _01533_ VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__clkbuf_1
X_23383_ _03251_ _03252_ VGND VGND VPWR VPWR _03253_ sky130_fd_sc_hd__and2b_1
X_20595_ _09069_ _12376_ _12315_ _09029_ VGND VGND VPWR VPWR _12377_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3748 _03456_ VGND VGND VPWR VPWR net3748 sky130_fd_sc_hd__buf_1
XFILLER_0_73_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25122_ pid_d.prev_int\[10\] net3033 _04852_ net9169 VGND VGND VPWR VPWR _00803_
+ sky130_fd_sc_hd__a22o_1
X_22334_ net336 _02324_ _02325_ VGND VGND VPWR VPWR _02337_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_115_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22265_ pid_d.prev_int\[11\] VGND VGND VPWR VPWR _02269_ sky130_fd_sc_hd__inv_2
X_25053_ net1628 _04802_ net2147 VGND VGND VPWR VPWR _04803_ sky130_fd_sc_hd__a21o_1
XFILLER_0_103_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24004_ net795 _03835_ VGND VGND VPWR VPWR _03867_ sky130_fd_sc_hd__nor2_1
X_21216_ _01027_ _01222_ _01231_ VGND VGND VPWR VPWR _01232_ sky130_fd_sc_hd__a21oi_1
X_22196_ _02200_ VGND VGND VPWR VPWR _02201_ sky130_fd_sc_hd__buf_1
Xwire3014 net3015 VGND VGND VPWR VPWR net3014 sky130_fd_sc_hd__clkbuf_1
Xwire3025 net3026 VGND VGND VPWR VPWR net3025 sky130_fd_sc_hd__clkbuf_1
Xwire3036 _04532_ VGND VGND VPWR VPWR net3036 sky130_fd_sc_hd__clkbuf_1
Xwire2302 _05419_ VGND VGND VPWR VPWR net2302 sky130_fd_sc_hd__buf_1
X_21147_ _01121_ _01162_ VGND VGND VPWR VPWR _01163_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3058 _03313_ VGND VGND VPWR VPWR net3058 sky130_fd_sc_hd__clkbuf_1
Xwire2313 net2314 VGND VGND VPWR VPWR net2313 sky130_fd_sc_hd__clkbuf_1
Xwire2324 _04974_ VGND VGND VPWR VPWR net2324 sky130_fd_sc_hd__buf_1
Xwire3069 _02682_ VGND VGND VPWR VPWR net3069 sky130_fd_sc_hd__clkbuf_1
Xwire2335 net2336 VGND VGND VPWR VPWR net2335 sky130_fd_sc_hd__buf_1
Xwire1601 net1602 VGND VGND VPWR VPWR net1601 sky130_fd_sc_hd__buf_1
Xwire2357 net2358 VGND VGND VPWR VPWR net2357 sky130_fd_sc_hd__buf_1
Xwire1612 net1613 VGND VGND VPWR VPWR net1612 sky130_fd_sc_hd__clkbuf_1
X_21078_ _01088_ _01090_ _01093_ VGND VGND VPWR VPWR _01094_ sky130_fd_sc_hd__a21o_1
Xwire2368 net2369 VGND VGND VPWR VPWR net2368 sky130_fd_sc_hd__buf_1
Xwire1623 net1624 VGND VGND VPWR VPWR net1623 sky130_fd_sc_hd__clkbuf_1
Xwire2379 net2380 VGND VGND VPWR VPWR net2379 sky130_fd_sc_hd__buf_1
X_24906_ net115 net118 net117 net120 VGND VGND VPWR VPWR _04696_ sky130_fd_sc_hd__or4_1
X_12920_ _05188_ _05192_ VGND VGND VPWR VPWR _05193_ sky130_fd_sc_hd__xnor2_1
X_20029_ net6134 net3132 net6077 VGND VGND VPWR VPWR _11859_ sky130_fd_sc_hd__or3_1
Xwire1656 _04093_ VGND VGND VPWR VPWR net1656 sky130_fd_sc_hd__buf_1
X_25886_ clknet_leaf_17_clk _00759_ net8632 VGND VGND VPWR VPWR pid_q.ki\[14\] sky130_fd_sc_hd__dfrtp_1
Xwire1667 net1668 VGND VGND VPWR VPWR net1667 sky130_fd_sc_hd__clkbuf_2
Xwire1678 _02931_ VGND VGND VPWR VPWR net1678 sky130_fd_sc_hd__buf_1
Xwire1689 net1690 VGND VGND VPWR VPWR net1689 sky130_fd_sc_hd__dlymetal6s2s_1
X_24837_ net4956 _04642_ net2001 net686 VGND VGND VPWR VPWR _00720_ sky130_fd_sc_hd__a22o_1
X_12851_ _05067_ _05068_ _05069_ VGND VGND VPWR VPWR _05124_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_68_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15570_ _07569_ _07635_ net674 VGND VGND VPWR VPWR _07642_ sky130_fd_sc_hd__a21oi_1
X_24768_ net7985 VGND VGND VPWR VPWR _04596_ sky130_fd_sc_hd__inv_2
X_12782_ _05053_ _05054_ VGND VGND VPWR VPWR _05055_ sky130_fd_sc_hd__and2_1
XFILLER_0_96_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14521_ _06692_ _06693_ _06700_ VGND VGND VPWR VPWR _06701_ sky130_fd_sc_hd__o21a_1
X_23719_ _03564_ net639 VGND VGND VPWR VPWR _03585_ sky130_fd_sc_hd__or2b_1
XFILLER_0_3_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24699_ net8034 net5307 VGND VGND VPWR VPWR _04536_ sky130_fd_sc_hd__or2b_1
X_17240_ svm0.state\[0\] VGND VGND VPWR VPWR _09187_ sky130_fd_sc_hd__inv_2
X_14452_ net8168 net4234 VGND VGND VPWR VPWR _06643_ sky130_fd_sc_hd__and2_1
X_13403_ _05674_ _05675_ VGND VGND VPWR VPWR _05676_ sky130_fd_sc_hd__nor2_1
XFILLER_0_187_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17171_ net1801 _09114_ _09113_ VGND VGND VPWR VPWR _09123_ sky130_fd_sc_hd__or3_1
Xwire920 net921 VGND VGND VPWR VPWR net920 sky130_fd_sc_hd__buf_1
X_14383_ _06590_ VGND VGND VPWR VPWR _00081_ sky130_fd_sc_hd__clkbuf_1
Xwire931 _04020_ VGND VGND VPWR VPWR net931 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire942 _02581_ VGND VGND VPWR VPWR net942 sky130_fd_sc_hd__clkbuf_1
Xwire953 net954 VGND VGND VPWR VPWR net953 sky130_fd_sc_hd__clkbuf_2
X_16122_ net3484 net3599 VGND VGND VPWR VPWR _08188_ sky130_fd_sc_hd__nor2_1
X_13334_ net7792 net2307 net1952 VGND VGND VPWR VPWR _05607_ sky130_fd_sc_hd__and3_1
Xwire964 _09570_ VGND VGND VPWR VPWR net964 sky130_fd_sc_hd__clkbuf_1
Xwire975 _08520_ VGND VGND VPWR VPWR net975 sky130_fd_sc_hd__buf_1
Xwire986 _07934_ VGND VGND VPWR VPWR net986 sky130_fd_sc_hd__clkbuf_1
Xwire997 _05739_ VGND VGND VPWR VPWR net997 sky130_fd_sc_hd__buf_1
X_16053_ _08019_ _08020_ _08119_ VGND VGND VPWR VPWR _08120_ sky130_fd_sc_hd__o21a_1
X_13265_ _05524_ _05537_ VGND VGND VPWR VPWR _05538_ sky130_fd_sc_hd__xor2_1
X_15004_ net4136 net4129 VGND VGND VPWR VPWR _07078_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13196_ _05467_ _05468_ VGND VGND VPWR VPWR _05469_ sky130_fd_sc_hd__or2_1
Xwire4260 net4261 VGND VGND VPWR VPWR net4260 sky130_fd_sc_hd__buf_1
Xwire4271 _04911_ VGND VGND VPWR VPWR net4271 sky130_fd_sc_hd__clkbuf_1
X_19812_ net6121 _11451_ VGND VGND VPWR VPWR _11646_ sky130_fd_sc_hd__nor2_1
Xwire4282 net4283 VGND VGND VPWR VPWR net4282 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4293 net4294 VGND VGND VPWR VPWR net4293 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3570 net3572 VGND VGND VPWR VPWR net3570 sky130_fd_sc_hd__buf_1
X_19743_ net3919 net3157 _11522_ net6275 VGND VGND VPWR VPWR _11578_ sky130_fd_sc_hd__o22a_1
Xwire3581 _07021_ VGND VGND VPWR VPWR net3581 sky130_fd_sc_hd__buf_1
X_16955_ _08856_ _08860_ net2176 net2174 _08903_ VGND VGND VPWR VPWR _08918_ sky130_fd_sc_hd__o221ai_1
Xwire3592 net3593 VGND VGND VPWR VPWR net3592 sky130_fd_sc_hd__buf_1
XFILLER_0_21_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15906_ _07973_ _07974_ VGND VGND VPWR VPWR _07975_ sky130_fd_sc_hd__and2_1
Xwire2880 _06801_ VGND VGND VPWR VPWR net2880 sky130_fd_sc_hd__buf_1
XFILLER_0_194_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19674_ _11505_ _11509_ VGND VGND VPWR VPWR _11510_ sky130_fd_sc_hd__xnor2_1
X_16886_ net6462 VGND VGND VPWR VPWR _08850_ sky130_fd_sc_hd__inv_2
Xwire2891 net2892 VGND VGND VPWR VPWR net2891 sky130_fd_sc_hd__buf_1
XFILLER_0_189_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15837_ _07892_ _07905_ VGND VGND VPWR VPWR _07907_ sky130_fd_sc_hd__nor2_1
X_18625_ net3988 net6893 net3232 VGND VGND VPWR VPWR _10472_ sky130_fd_sc_hd__or3_1
XFILLER_0_78_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18556_ _10333_ _10332_ _10397_ VGND VGND VPWR VPWR _10404_ sky130_fd_sc_hd__mux2_1
X_15768_ net3400 VGND VGND VPWR VPWR _07838_ sky130_fd_sc_hd__buf_1
X_17507_ _09311_ _09388_ net4016 VGND VGND VPWR VPWR _09394_ sky130_fd_sc_hd__o21a_1
X_14719_ net7457 _06858_ net7148 VGND VGND VPWR VPWR _06859_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_157_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18487_ _10249_ _10254_ _10252_ VGND VGND VPWR VPWR _10337_ sky130_fd_sc_hd__a21bo_1
X_15699_ _07518_ _07769_ _07697_ VGND VGND VPWR VPWR _07770_ sky130_fd_sc_hd__a21bo_1
X_17438_ net6741 net7376 VGND VGND VPWR VPWR _09335_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17369_ _09280_ VGND VGND VPWR VPWR _00377_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19108_ _10943_ _10944_ net6302 VGND VGND VPWR VPWR _10945_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20380_ net6374 _12159_ _12168_ net1054 VGND VGND VPWR VPWR _12179_ sky130_fd_sc_hd__a211o_1
XFILLER_0_63_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19039_ net6229 _10875_ VGND VGND VPWR VPWR _10876_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_24_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22050_ net5380 _02056_ VGND VGND VPWR VPWR _02057_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21001_ _00998_ _01002_ VGND VGND VPWR VPWR _01017_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25740_ clknet_leaf_13_clk _00613_ net8604 VGND VGND VPWR VPWR pid_d.ki\[14\] sky130_fd_sc_hd__dfrtp_1
X_22952_ _02839_ _02515_ _02838_ _02387_ VGND VGND VPWR VPWR _02840_ sky130_fd_sc_hd__o22a_1
XFILLER_0_179_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21903_ _01910_ _01911_ VGND VGND VPWR VPWR _01912_ sky130_fd_sc_hd__nand2_1
X_25671_ clknet_leaf_4_clk _00544_ net8568 VGND VGND VPWR VPWR pid_d.prev_error\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_22883_ _01917_ _02770_ net5360 VGND VGND VPWR VPWR _02778_ sky130_fd_sc_hd__o21ba_1
X_24622_ net3047 _04476_ VGND VGND VPWR VPWR _04477_ sky130_fd_sc_hd__or2_1
X_21834_ _01831_ _01842_ VGND VGND VPWR VPWR _01843_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_195_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24553_ _04405_ _04407_ VGND VGND VPWR VPWR _04409_ sky130_fd_sc_hd__nand2_1
XFILLER_0_194_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21765_ _01767_ _01774_ VGND VGND VPWR VPWR _01775_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_148_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8504 net8501 VGND VGND VPWR VPWR net8504 sky130_fd_sc_hd__buf_1
X_23504_ _03372_ VGND VGND VPWR VPWR _03373_ sky130_fd_sc_hd__buf_1
Xmax_length4202 net4203 VGND VGND VPWR VPWR net4202 sky130_fd_sc_hd__buf_1
Xwire8515 net8516 VGND VGND VPWR VPWR net8515 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20716_ net6764 net5998 VGND VGND VPWR VPWR _12488_ sky130_fd_sc_hd__xnor2_1
Xwire8526 net8527 VGND VGND VPWR VPWR net8526 sky130_fd_sc_hd__clkbuf_1
X_24484_ _04200_ _04202_ _04340_ net4515 VGND VGND VPWR VPWR _04341_ sky130_fd_sc_hd__a2bb2o_1
Xmax_length4224 _06826_ VGND VGND VPWR VPWR net4224 sky130_fd_sc_hd__clkbuf_1
Xmax_length4235 _06512_ VGND VGND VPWR VPWR net4235 sky130_fd_sc_hd__buf_1
X_21696_ net1173 _01706_ VGND VGND VPWR VPWR _01707_ sky130_fd_sc_hd__xor2_1
Xwire8548 net8549 VGND VGND VPWR VPWR net8548 sky130_fd_sc_hd__clkbuf_1
Xwire7814 net7815 VGND VGND VPWR VPWR net7814 sky130_fd_sc_hd__buf_1
Xwire8559 net8560 VGND VGND VPWR VPWR net8559 sky130_fd_sc_hd__clkbuf_2
Xwire205 _02459_ VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__buf_1
XFILLER_0_80_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23435_ _03299_ _03304_ VGND VGND VPWR VPWR _03305_ sky130_fd_sc_hd__xnor2_1
Xwire7825 net7826 VGND VGND VPWR VPWR net7825 sky130_fd_sc_hd__buf_1
Xwire216 _08489_ VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_1
Xwire227 net228 VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__buf_1
Xwire7836 net7843 VGND VGND VPWR VPWR net7836 sky130_fd_sc_hd__buf_1
X_20647_ net8058 net3147 _12424_ _12425_ VGND VGND VPWR VPWR _00511_ sky130_fd_sc_hd__a31o_1
XFILLER_0_34_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7847 net7848 VGND VGND VPWR VPWR net7847 sky130_fd_sc_hd__buf_1
Xmax_length3534 net3535 VGND VGND VPWR VPWR net3534 sky130_fd_sc_hd__buf_1
Xwire238 _04170_ VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__buf_1
XFILLER_0_191_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire7858 net7859 VGND VGND VPWR VPWR net7858 sky130_fd_sc_hd__clkbuf_1
Xwire249 net250 VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__clkbuf_1
Xwire7869 net7870 VGND VGND VPWR VPWR net7869 sky130_fd_sc_hd__clkbuf_1
X_23366_ _03231_ _03235_ VGND VGND VPWR VPWR _03236_ sky130_fd_sc_hd__and2_1
X_20578_ net3174 _12360_ _12361_ VGND VGND VPWR VPWR _00506_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25105_ net196 _04829_ VGND VGND VPWR VPWR _04848_ sky130_fd_sc_hd__nor2_1
X_22317_ net2058 net943 VGND VGND VPWR VPWR _02321_ sky130_fd_sc_hd__nor2_1
Xmax_length2866 _06824_ VGND VGND VPWR VPWR net2866 sky130_fd_sc_hd__buf_1
XFILLER_0_147_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23297_ _03154_ _03151_ VGND VGND VPWR VPWR _03167_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25036_ net405 net1630 _04786_ net9166 _04788_ VGND VGND VPWR VPWR _00782_ sky130_fd_sc_hd__a221o_1
X_13050_ net851 VGND VGND VPWR VPWR _05323_ sky130_fd_sc_hd__inv_2
X_22248_ _02251_ _02252_ VGND VGND VPWR VPWR _02253_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22179_ _02182_ _02111_ _02183_ VGND VGND VPWR VPWR _02184_ sky130_fd_sc_hd__o21a_1
Xwire2110 _10953_ VGND VGND VPWR VPWR net2110 sky130_fd_sc_hd__buf_1
Xwire2121 net2124 VGND VGND VPWR VPWR net2121 sky130_fd_sc_hd__buf_1
Xwire2132 net2133 VGND VGND VPWR VPWR net2132 sky130_fd_sc_hd__clkbuf_1
Xwire2143 net2144 VGND VGND VPWR VPWR net2143 sky130_fd_sc_hd__clkbuf_2
Xwire2165 _09185_ VGND VGND VPWR VPWR net2165 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1420 _11305_ VGND VGND VPWR VPWR net1420 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2176 _08883_ VGND VGND VPWR VPWR net2176 sky130_fd_sc_hd__buf_1
Xwire1431 net1432 VGND VGND VPWR VPWR net1431 sky130_fd_sc_hd__buf_1
X_16740_ _08758_ VGND VGND VPWR VPWR _00270_ sky130_fd_sc_hd__clkbuf_1
X_13952_ _06158_ _06213_ _06214_ VGND VGND VPWR VPWR _06217_ sky130_fd_sc_hd__o21a_1
X_25938_ clknet_4_4__leaf_clk net2997 net8556 VGND VGND VPWR VPWR pid_d.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire2187 _08841_ VGND VGND VPWR VPWR net2187 sky130_fd_sc_hd__buf_1
Xwire1442 _10274_ VGND VGND VPWR VPWR net1442 sky130_fd_sc_hd__clkbuf_1
Xwire1453 net1454 VGND VGND VPWR VPWR net1453 sky130_fd_sc_hd__buf_1
Xwire2198 net2199 VGND VGND VPWR VPWR net2198 sky130_fd_sc_hd__clkbuf_1
Xwire1464 net1465 VGND VGND VPWR VPWR net1464 sky130_fd_sc_hd__clkbuf_1
X_12903_ _05095_ _05096_ _05175_ VGND VGND VPWR VPWR _05176_ sky130_fd_sc_hd__o21a_1
Xwire1475 _09068_ VGND VGND VPWR VPWR net1475 sky130_fd_sc_hd__buf_1
Xwire1486 _08952_ VGND VGND VPWR VPWR net1486 sky130_fd_sc_hd__buf_1
X_16671_ matmul0.matmul_stage_inst.mult1\[7\] VGND VGND VPWR VPWR _08704_ sky130_fd_sc_hd__inv_2
X_25869_ clknet_leaf_18_clk _00742_ net8630 VGND VGND VPWR VPWR pid_q.mult0.a\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13883_ _06145_ _06147_ net449 VGND VGND VPWR VPWR _06150_ sky130_fd_sc_hd__mux2_1
Xwire1497 _08916_ VGND VGND VPWR VPWR net1497 sky130_fd_sc_hd__clkbuf_1
X_18410_ net1786 VGND VGND VPWR VPWR _10261_ sky130_fd_sc_hd__buf_1
X_15622_ _07692_ VGND VGND VPWR VPWR _07694_ sky130_fd_sc_hd__buf_1
X_12834_ _05103_ _05106_ VGND VGND VPWR VPWR _05107_ sky130_fd_sc_hd__xnor2_1
X_19390_ net2509 _11157_ _11220_ VGND VGND VPWR VPWR _11227_ sky130_fd_sc_hd__a21o_1
XFILLER_0_185_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18341_ _10186_ _10191_ VGND VGND VPWR VPWR _10192_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_189_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15553_ net889 _07625_ VGND VGND VPWR VPWR _07626_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12765_ _05033_ net1604 VGND VGND VPWR VPWR _05038_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_68_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14504_ net7313 net5269 VGND VGND VPWR VPWR _06686_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18272_ net6832 net6881 VGND VGND VPWR VPWR _10123_ sky130_fd_sc_hd__nand2_1
X_15484_ _07557_ net675 VGND VGND VPWR VPWR _07558_ sky130_fd_sc_hd__nand2_1
X_12696_ _04950_ _04951_ _04968_ VGND VGND VPWR VPWR _04969_ sky130_fd_sc_hd__o21ai_2
X_17223_ net6806 _09165_ VGND VGND VPWR VPWR _09171_ sky130_fd_sc_hd__nor2_1
X_14435_ _06630_ VGND VGND VPWR VPWR _00093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput13 angle_in[6] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_1
XFILLER_0_64_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput24 currA_in[1] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17154_ net2199 _09107_ net8048 VGND VGND VPWR VPWR _09108_ sky130_fd_sc_hd__o21a_1
Xwire750 net751 VGND VGND VPWR VPWR net750 sky130_fd_sc_hd__clkbuf_1
Xmax_length4791 net4792 VGND VGND VPWR VPWR net4791 sky130_fd_sc_hd__buf_1
Xinput35 currB_in[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_1
X_14366_ _06577_ matmul0.a_in\[10\] _06572_ VGND VGND VPWR VPWR _06578_ sky130_fd_sc_hd__mux2_1
Xwire761 net762 VGND VGND VPWR VPWR net761 sky130_fd_sc_hd__buf_1
Xinput46 currB_in[7] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_1
Xinput57 currT_in[2] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire772 _09046_ VGND VGND VPWR VPWR net772 sky130_fd_sc_hd__buf_1
XFILLER_0_13_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput68 periodTop[12] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_1
X_16105_ net3561 _07684_ net4075 net2840 VGND VGND VPWR VPWR _08171_ sky130_fd_sc_hd__o2bb2a_1
Xwire783 net784 VGND VGND VPWR VPWR net783 sky130_fd_sc_hd__buf_1
X_13317_ _05581_ _05589_ VGND VGND VPWR VPWR _05590_ sky130_fd_sc_hd__xor2_1
XFILLER_0_134_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire794 _04053_ VGND VGND VPWR VPWR net794 sky130_fd_sc_hd__clkbuf_1
Xinput79 periodTop[8] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_1
X_17085_ net3328 _09019_ _09041_ VGND VGND VPWR VPWR _09043_ sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_172_Right_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14297_ net71 net3649 net2915 net7614 VGND VGND VPWR VPWR _00066_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16036_ _08038_ _08039_ _08102_ VGND VGND VPWR VPWR _08103_ sky130_fd_sc_hd__o21a_1
X_13248_ net7821 net2304 net2964 VGND VGND VPWR VPWR _05521_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_196_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13179_ net7732 net1983 net2361 VGND VGND VPWR VPWR _05452_ sky130_fd_sc_hd__and3_1
Xwire4090 net4091 VGND VGND VPWR VPWR net4090 sky130_fd_sc_hd__clkbuf_1
X_17987_ _09826_ _09837_ net1447 VGND VGND VPWR VPWR _09838_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19726_ _11449_ _11508_ _11431_ VGND VGND VPWR VPWR _11561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16938_ _08854_ _08901_ _08852_ VGND VGND VPWR VPWR _08902_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19657_ _11454_ _11456_ VGND VGND VPWR VPWR _11493_ sky130_fd_sc_hd__nand2_1
X_16869_ net6020 net5997 net6523 VGND VGND VPWR VPWR _08834_ sky130_fd_sc_hd__mux2_1
X_18608_ net814 _10455_ VGND VGND VPWR VPWR _10456_ sky130_fd_sc_hd__xnor2_2
X_19588_ _11419_ _11422_ VGND VGND VPWR VPWR _11425_ sky130_fd_sc_hd__nor2_1
XFILLER_0_177_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18539_ _10387_ net2541 _10221_ VGND VGND VPWR VPWR _10388_ sky130_fd_sc_hd__o21a_1
XFILLER_0_176_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21550_ net5743 net5537 VGND VGND VPWR VPWR _01562_ sky130_fd_sc_hd__nand2_2
XFILLER_0_30_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20501_ net1484 _12287_ net3169 VGND VGND VPWR VPWR _12288_ sky130_fd_sc_hd__a21oi_1
X_21481_ _01489_ _01493_ VGND VGND VPWR VPWR _01494_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6409 cordic0.slte0.opB\[8\] VGND VGND VPWR VPWR net6409 sky130_fd_sc_hd__clkbuf_1
X_23220_ _03048_ _03069_ _03072_ _03089_ VGND VGND VPWR VPWR _03090_ sky130_fd_sc_hd__a2bb2o_1
X_20432_ _12205_ _12210_ net863 cordic0.slte0.opA\[11\] _12219_ VGND VGND VPWR VPWR
+ _12227_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5708 net5709 VGND VGND VPWR VPWR net5708 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire5719 net5718 VGND VGND VPWR VPWR net5719 sky130_fd_sc_hd__buf_1
X_23151_ net5064 net4716 VGND VGND VPWR VPWR _03021_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20363_ net6374 _12162_ _12163_ _12161_ VGND VGND VPWR VPWR _00489_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22102_ pid_d.prev_int\[9\] VGND VGND VPWR VPWR _02108_ sky130_fd_sc_hd__inv_2
X_23082_ _02950_ _02951_ VGND VGND VPWR VPWR _02952_ sky130_fd_sc_hd__xnor2_1
X_20294_ _12094_ _12099_ net2608 VGND VGND VPWR VPWR _12100_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22033_ net5763 net5410 VGND VGND VPWR VPWR _02040_ sky130_fd_sc_hd__nand2_1
X_23984_ _03847_ VGND VGND VPWR VPWR _03848_ sky130_fd_sc_hd__inv_2
X_25723_ clknet_leaf_13_clk _00596_ net8609 VGND VGND VPWR VPWR pid_d.mult0.a\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22935_ net5327 _02824_ net3064 VGND VGND VPWR VPWR _02825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25654_ clknet_leaf_2_clk _00527_ net8570 VGND VGND VPWR VPWR pid_d.curr_int\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22866_ net5363 net5979 VGND VGND VPWR VPWR _02763_ sky130_fd_sc_hd__xnor2_1
X_24605_ _04408_ _04438_ VGND VGND VPWR VPWR _04460_ sky130_fd_sc_hd__nand2_1
XFILLER_0_168_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21817_ _01804_ _01806_ VGND VGND VPWR VPWR _01826_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_196_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25585_ clknet_leaf_91_clk _00458_ net8428 VGND VGND VPWR VPWR cordic0.cos\[5\] sky130_fd_sc_hd__dfrtp_1
X_22797_ _02706_ VGND VGND VPWR VPWR _00625_ sky130_fd_sc_hd__clkbuf_1
Xwire8301 net8302 VGND VGND VPWR VPWR net8301 sky130_fd_sc_hd__clkbuf_1
X_24536_ _04390_ _04391_ VGND VGND VPWR VPWR _04392_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_159_Left_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21748_ net5725 net5515 VGND VGND VPWR VPWR _01758_ sky130_fd_sc_hd__nand2_1
Xwire8312 net8313 VGND VGND VPWR VPWR net8312 sky130_fd_sc_hd__clkbuf_1
Xwire8323 net8324 VGND VGND VPWR VPWR net8323 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7600 matmul0.a_in\[8\] VGND VGND VPWR VPWR net7600 sky130_fd_sc_hd__clkbuf_1
X_24467_ pid_q.prev_error\[11\] pid_q.curr_error\[11\] _04324_ VGND VGND VPWR VPWR
+ _04325_ sky130_fd_sc_hd__a21oi_1
Xwire7622 net7623 VGND VGND VPWR VPWR net7622 sky130_fd_sc_hd__clkbuf_1
Xfanout6815 net6822 VGND VGND VPWR VPWR net6815 sky130_fd_sc_hd__buf_1
XFILLER_0_65_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21679_ net5859 net5401 VGND VGND VPWR VPWR _01690_ sky130_fd_sc_hd__nand2_1
Xwire8367 net8368 VGND VGND VPWR VPWR net8367 sky130_fd_sc_hd__buf_1
XFILLER_0_0_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8378 net8379 VGND VGND VPWR VPWR net8378 sky130_fd_sc_hd__clkbuf_1
Xwire7644 net7645 VGND VGND VPWR VPWR net7644 sky130_fd_sc_hd__clkbuf_1
X_14220_ _06463_ _06478_ VGND VGND VPWR VPWR _06479_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_149_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8389 net8390 VGND VGND VPWR VPWR net8389 sky130_fd_sc_hd__buf_1
X_23418_ _03217_ _03218_ _03219_ VGND VGND VPWR VPWR _03288_ sky130_fd_sc_hd__o21a_1
Xwire7655 net7656 VGND VGND VPWR VPWR net7655 sky130_fd_sc_hd__buf_1
Xwire6910 net6911 VGND VGND VPWR VPWR net6910 sky130_fd_sc_hd__buf_1
XFILLER_0_184_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7666 net7667 VGND VGND VPWR VPWR net7666 sky130_fd_sc_hd__buf_1
Xwire6921 net6919 VGND VGND VPWR VPWR net6921 sky130_fd_sc_hd__buf_1
X_24398_ net7506 _04255_ _04256_ VGND VGND VPWR VPWR _04257_ sky130_fd_sc_hd__and3_1
Xwire7677 net7678 VGND VGND VPWR VPWR net7677 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6943 net6944 VGND VGND VPWR VPWR net6943 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire7699 net7691 VGND VGND VPWR VPWR net7699 sky130_fd_sc_hd__buf_1
X_14151_ _06378_ _06380_ VGND VGND VPWR VPWR _06412_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6954 net6955 VGND VGND VPWR VPWR net6954 sky130_fd_sc_hd__clkbuf_1
X_23349_ net4990 net4667 VGND VGND VPWR VPWR _03219_ sky130_fd_sc_hd__nand2_1
Xwire6965 net6969 VGND VGND VPWR VPWR net6965 sky130_fd_sc_hd__buf_1
Xwire6976 net6977 VGND VGND VPWR VPWR net6976 sky130_fd_sc_hd__clkbuf_2
Xwire6987 net6989 VGND VGND VPWR VPWR net6987 sky130_fd_sc_hd__clkbuf_1
X_13102_ net7735 _04904_ net2989 VGND VGND VPWR VPWR _05375_ sky130_fd_sc_hd__and3_1
Xmax_length1951 _05134_ VGND VGND VPWR VPWR net1951 sky130_fd_sc_hd__clkbuf_1
X_14082_ _06341_ _06344_ VGND VGND VPWR VPWR _06345_ sky130_fd_sc_hd__xnor2_1
X_25019_ _03578_ _04768_ net4462 VGND VGND VPWR VPWR _04773_ sky130_fd_sc_hd__o21ba_1
X_13033_ _05246_ _05248_ net684 VGND VGND VPWR VPWR _05306_ sky130_fd_sc_hd__a21o_1
X_17910_ _09747_ _09760_ VGND VGND VPWR VPWR _09761_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_168_Left_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18890_ net1437 _10731_ VGND VGND VPWR VPWR _10732_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17841_ _09690_ net2558 VGND VGND VPWR VPWR _09692_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17772_ net7116 net7092 VGND VGND VPWR VPWR _09623_ sky130_fd_sc_hd__or2b_1
X_14984_ _07056_ _07057_ VGND VGND VPWR VPWR _07058_ sky130_fd_sc_hd__xnor2_1
Xwire1250 _08262_ VGND VGND VPWR VPWR net1250 sky130_fd_sc_hd__buf_2
XFILLER_0_191_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19511_ net6067 net6103 VGND VGND VPWR VPWR _11348_ sky130_fd_sc_hd__nand2_2
Xwire1261 _08035_ VGND VGND VPWR VPWR net1261 sky130_fd_sc_hd__buf_1
X_13935_ _06098_ _06103_ _06200_ VGND VGND VPWR VPWR _06201_ sky130_fd_sc_hd__o21a_1
XFILLER_0_135_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1272 _07587_ VGND VGND VPWR VPWR net1272 sky130_fd_sc_hd__buf_1
XFILLER_0_92_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16723_ _08742_ _08747_ _08748_ VGND VGND VPWR VPWR _08749_ sky130_fd_sc_hd__o21a_1
Xwire1283 net1284 VGND VGND VPWR VPWR net1283 sky130_fd_sc_hd__buf_1
XFILLER_0_117_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1294 _06608_ VGND VGND VPWR VPWR net1294 sky130_fd_sc_hd__buf_1
XFILLER_0_159_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19442_ _11276_ _11277_ net3161 _11275_ VGND VGND VPWR VPWR _11279_ sky130_fd_sc_hd__o211ai_2
X_16654_ _08688_ _08689_ VGND VGND VPWR VPWR _08690_ sky130_fd_sc_hd__xnor2_1
X_13866_ net7788 net1930 VGND VGND VPWR VPWR _06133_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15605_ _07613_ _07615_ _07614_ VGND VGND VPWR VPWR _07677_ sky130_fd_sc_hd__a21o_1
X_12817_ net7824 net2370 net2367 VGND VGND VPWR VPWR _05090_ sky130_fd_sc_hd__and3_1
X_19373_ net3166 net2523 VGND VGND VPWR VPWR _11210_ sky130_fd_sc_hd__nand2_1
X_16585_ matmul0.matmul_stage_inst.mult2\[3\] net426 net2619 VGND VGND VPWR VPWR _08640_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_177_Left_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13797_ _05954_ _05957_ VGND VGND VPWR VPWR _06065_ sky130_fd_sc_hd__nor2_1
XFILLER_0_158_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15536_ net1857 _07608_ VGND VGND VPWR VPWR _07609_ sky130_fd_sc_hd__xnor2_1
X_18324_ net6872 _10102_ _10173_ net3947 _10174_ VGND VGND VPWR VPWR _10175_ sky130_fd_sc_hd__a221o_1
XFILLER_0_84_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12748_ net7907 VGND VGND VPWR VPWR _05021_ sky130_fd_sc_hd__inv_2
Xfanout8751 net8793 VGND VGND VPWR VPWR net8751 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8773 net8800 VGND VGND VPWR VPWR net8773 sky130_fd_sc_hd__buf_1
XFILLER_0_155_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18255_ _10100_ _10101_ _10105_ VGND VGND VPWR VPWR _10106_ sky130_fd_sc_hd__a21o_1
Xfanout8784 net8790 VGND VGND VPWR VPWR net8784 sky130_fd_sc_hd__buf_1
X_15467_ net1113 _07540_ VGND VGND VPWR VPWR _07541_ sky130_fd_sc_hd__xnor2_2
X_12679_ _04950_ _04951_ VGND VGND VPWR VPWR _04952_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17206_ net6810 VGND VGND VPWR VPWR _09156_ sky130_fd_sc_hd__inv_2
X_14418_ _06617_ matmul0.b_in\[6\] net896 VGND VGND VPWR VPWR _06618_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18186_ net7032 net7124 VGND VGND VPWR VPWR _10037_ sky130_fd_sc_hd__xnor2_4
X_15398_ _07342_ _07411_ VGND VGND VPWR VPWR _07472_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17137_ net6914 _09090_ _09091_ VGND VGND VPWR VPWR _00334_ sky130_fd_sc_hd__a21bo_1
Xwire580 _05769_ VGND VGND VPWR VPWR net580 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14349_ net7291 net1301 net2899 net5358 _06563_ VGND VGND VPWR VPWR _06564_ sky130_fd_sc_hd__a221o_1
XFILLER_0_170_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire591 _04025_ VGND VGND VPWR VPWR net591 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17068_ _09024_ _09025_ _09026_ VGND VGND VPWR VPWR _09027_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_186_Left_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16019_ matmul0.matmul_stage_inst.mult1\[6\] net359 net2679 VGND VGND VPWR VPWR _08087_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19709_ _11488_ _11542_ VGND VGND VPWR VPWR _11545_ sky130_fd_sc_hd__nor2_1
Xmax_length7608 net7609 VGND VGND VPWR VPWR net7608 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20981_ net5527 net5884 VGND VGND VPWR VPWR _00997_ sky130_fd_sc_hd__nand2_1
X_22720_ net8107 net8105 net84 net8103 VGND VGND VPWR VPWR _02656_ sky130_fd_sc_hd__or4_1
XFILLER_0_177_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_195_Left_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length6918 net6914 VGND VGND VPWR VPWR net6918 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_178_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22651_ net9154 net3086 _02610_ _02014_ net8901 VGND VGND VPWR VPWR _00575_ sky130_fd_sc_hd__o221a_1
XFILLER_0_75_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21602_ _01612_ _01613_ VGND VGND VPWR VPWR _01614_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25370_ clknet_leaf_81_clk _00253_ net8500 VGND VGND VPWR VPWR matmul0.alpha_pass\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_193_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22582_ pid_d.curr_error\[4\] net2040 net3087 VGND VGND VPWR VPWR _02562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24321_ pid_q.prev_error\[10\] pid_q.curr_error\[10\] VGND VGND VPWR VPWR _04181_
+ sky130_fd_sc_hd__xnor2_1
X_21533_ net860 net806 _01418_ VGND VGND VPWR VPWR _01545_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24252_ _04111_ _04112_ VGND VGND VPWR VPWR _04113_ sky130_fd_sc_hd__nand2_1
Xwire6217 net6215 VGND VGND VPWR VPWR net6217 sky130_fd_sc_hd__buf_1
XFILLER_0_7_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21464_ net1726 _01476_ VGND VGND VPWR VPWR _01477_ sky130_fd_sc_hd__nor2_1
Xwire6239 net6233 VGND VGND VPWR VPWR net6239 sky130_fd_sc_hd__buf_1
X_23203_ net5111 net4756 net4772 net5089 VGND VGND VPWR VPWR _03073_ sky130_fd_sc_hd__a22o_1
Xwire5516 net5517 VGND VGND VPWR VPWR net5516 sky130_fd_sc_hd__buf_1
X_20415_ _06506_ _12211_ net4239 VGND VGND VPWR VPWR _12212_ sky130_fd_sc_hd__a21o_1
XFILLER_0_161_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24183_ _04022_ net590 VGND VGND VPWR VPWR _04044_ sky130_fd_sc_hd__nor2_1
Xmax_length1214 net1215 VGND VGND VPWR VPWR net1214 sky130_fd_sc_hd__clkbuf_2
X_21395_ _01400_ _01408_ VGND VGND VPWR VPWR _01409_ sky130_fd_sc_hd__xnor2_1
Xwire5527 net5528 VGND VGND VPWR VPWR net5527 sky130_fd_sc_hd__buf_1
Xwire5538 net5539 VGND VGND VPWR VPWR net5538 sky130_fd_sc_hd__buf_1
XFILLER_0_4_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5549 net5550 VGND VGND VPWR VPWR net5549 sky130_fd_sc_hd__buf_1
X_23134_ _02917_ _03003_ VGND VGND VPWR VPWR _03004_ sky130_fd_sc_hd__xnor2_1
Xwire4815 net4816 VGND VGND VPWR VPWR net4815 sky130_fd_sc_hd__clkbuf_1
X_20346_ net1500 net1054 _12147_ VGND VGND VPWR VPWR _12148_ sky130_fd_sc_hd__mux2_1
Xwire4837 net4838 VGND VGND VPWR VPWR net4837 sky130_fd_sc_hd__buf_1
XFILLER_0_144_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4859 net4860 VGND VGND VPWR VPWR net4859 sky130_fd_sc_hd__clkbuf_1
X_23065_ net5118 net4574 VGND VGND VPWR VPWR _02935_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20277_ net4041 net6472 VGND VGND VPWR VPWR _12084_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22016_ _01928_ _01930_ _01929_ VGND VGND VPWR VPWR _02023_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length8810 net8811 VGND VGND VPWR VPWR net8810 sky130_fd_sc_hd__buf_1
X_23967_ net3048 _03830_ VGND VGND VPWR VPWR _03831_ sky130_fd_sc_hd__xnor2_1
X_13720_ _05987_ _05988_ VGND VGND VPWR VPWR _05989_ sky130_fd_sc_hd__xnor2_1
X_25706_ clknet_leaf_6_clk _00579_ net8562 VGND VGND VPWR VPWR pid_d.mult0.b\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_22918_ net5339 net3104 VGND VGND VPWR VPWR _02809_ sky130_fd_sc_hd__nor2_1
X_23898_ _03762_ _03664_ pid_q.prev_error\[4\] VGND VGND VPWR VPWR _03763_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_116_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13651_ _05803_ _05920_ VGND VGND VPWR VPWR _05921_ sky130_fd_sc_hd__nand2_2
X_25637_ clknet_leaf_103_clk _00510_ net8375 VGND VGND VPWR VPWR cordic0.vec\[0\]\[9\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_39_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22849_ pid_d.out\[4\] net5981 VGND VGND VPWR VPWR _02748_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12602_ net8864 net7530 pid_q.state\[0\] VGND VGND VPWR VPWR _04880_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16370_ matmul0.matmul_stage_inst.mult1\[11\] net276 net3478 VGND VGND VPWR VPWR
+ _08433_ sky130_fd_sc_hd__mux2_1
X_13582_ net504 _05773_ VGND VGND VPWR VPWR _05853_ sky130_fd_sc_hd__nor2_1
X_25568_ clknet_leaf_98_clk _00441_ net8383 VGND VGND VPWR VPWR cordic0.sin\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8058 net8074 VGND VGND VPWR VPWR net8058 sky130_fd_sc_hd__buf_1
X_15321_ _07011_ _07015_ _07024_ _07031_ VGND VGND VPWR VPWR _07395_ sky130_fd_sc_hd__a22o_1
X_24519_ net792 _04315_ _04314_ VGND VGND VPWR VPWR _04376_ sky130_fd_sc_hd__a21bo_1
Xwire8131 net47 VGND VGND VPWR VPWR net8131 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_186_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8142 net8143 VGND VGND VPWR VPWR net8142 sky130_fd_sc_hd__clkbuf_1
X_25499_ clknet_leaf_41_clk _00379_ net8782 VGND VGND VPWR VPWR svm0.delta\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8153 net8154 VGND VGND VPWR VPWR net8153 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8164 net8165 VGND VGND VPWR VPWR net8164 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8175 net8176 VGND VGND VPWR VPWR net8175 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18040_ net7050 _09888_ net3237 _09890_ VGND VGND VPWR VPWR _09891_ sky130_fd_sc_hd__o2bb2a_2
Xwire7430 net7431 VGND VGND VPWR VPWR net7430 sky130_fd_sc_hd__clkbuf_1
X_15252_ net1878 _07313_ _07325_ VGND VGND VPWR VPWR _07326_ sky130_fd_sc_hd__a21oi_1
Xwire7441 net7442 VGND VGND VPWR VPWR net7441 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_191_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8186 net8187 VGND VGND VPWR VPWR net8186 sky130_fd_sc_hd__clkbuf_1
Xfanout6656 net6671 VGND VGND VPWR VPWR net6656 sky130_fd_sc_hd__buf_1
Xwire8197 net34 VGND VGND VPWR VPWR net8197 sky130_fd_sc_hd__clkbuf_1
Xwire7452 matmul0.op\[1\] VGND VGND VPWR VPWR net7452 sky130_fd_sc_hd__buf_1
XFILLER_0_163_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7463 net7465 VGND VGND VPWR VPWR net7463 sky130_fd_sc_hd__buf_1
XFILLER_0_81_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14203_ net9126 _05779_ net160 net2373 VGND VGND VPWR VPWR _00029_ sky130_fd_sc_hd__a22o_1
Xwire7474 net7470 VGND VGND VPWR VPWR net7474 sky130_fd_sc_hd__clkbuf_1
Xwire6740 net6741 VGND VGND VPWR VPWR net6740 sky130_fd_sc_hd__buf_1
Xwire7485 net7486 VGND VGND VPWR VPWR net7485 sky130_fd_sc_hd__buf_1
Xwire6751 net6752 VGND VGND VPWR VPWR net6751 sky130_fd_sc_hd__clkbuf_1
X_15183_ _07235_ _07256_ VGND VGND VPWR VPWR _07257_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire6762 net6763 VGND VGND VPWR VPWR net6762 sky130_fd_sc_hd__buf_1
Xwire6773 net6774 VGND VGND VPWR VPWR net6773 sky130_fd_sc_hd__buf_1
X_14134_ _06394_ _06395_ VGND VGND VPWR VPWR _06396_ sky130_fd_sc_hd__nand2_1
Xfanout5988 net5991 VGND VGND VPWR VPWR net5988 sky130_fd_sc_hd__buf_1
Xwire6784 net6785 VGND VGND VPWR VPWR net6784 sky130_fd_sc_hd__buf_1
Xfanout5999 net6003 VGND VGND VPWR VPWR net5999 sky130_fd_sc_hd__buf_1
X_19991_ _11819_ _11821_ VGND VGND VPWR VPWR _11822_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14065_ net7680 net1122 _06301_ VGND VGND VPWR VPWR _06328_ sky130_fd_sc_hd__a21o_1
X_18942_ net6375 _10772_ net207 VGND VGND VPWR VPWR _10781_ sky130_fd_sc_hd__a21oi_1
X_13016_ net7908 _05189_ net2965 VGND VGND VPWR VPWR _05289_ sky130_fd_sc_hd__and3_1
X_18873_ net3934 _10714_ net6794 VGND VGND VPWR VPWR _10715_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17824_ net6943 _09674_ VGND VGND VPWR VPWR _09675_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_146_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2 matmul0.matmul_stage_inst.c\[6\] VGND VGND VPWR VPWR net8955 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14967_ net3584 net3577 VGND VGND VPWR VPWR _07041_ sky130_fd_sc_hd__nor2_1
X_17755_ net7030 net7022 VGND VGND VPWR VPWR _09606_ sky130_fd_sc_hd__nor2b_1
Xwire1080 _08410_ VGND VGND VPWR VPWR net1080 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1091 _08182_ VGND VGND VPWR VPWR net1091 sky130_fd_sc_hd__buf_1
X_16706_ matmul0.matmul_stage_inst.mult1\[12\] VGND VGND VPWR VPWR _08734_ sky130_fd_sc_hd__inv_2
X_13918_ net7641 _06176_ _06180_ net1961 _06183_ VGND VGND VPWR VPWR _06184_ sky130_fd_sc_hd__o221a_1
X_17686_ net3272 svm0.tA\[11\] _09536_ _09565_ VGND VGND VPWR VPWR _09566_ sky130_fd_sc_hd__a22o_1
X_14898_ net6631 matmul0.matmul_stage_inst.d\[9\] net7408 net6533 VGND VGND VPWR VPWR
+ _06972_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19425_ net6333 net6241 VGND VGND VPWR VPWR _11262_ sky130_fd_sc_hd__and2b_1
X_13849_ net7610 net1962 VGND VGND VPWR VPWR _06116_ sky130_fd_sc_hd__nand2_1
X_16637_ _08672_ _08674_ VGND VGND VPWR VPWR _08675_ sky130_fd_sc_hd__nand2_1
XFILLER_0_162_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19356_ net3204 _11192_ VGND VGND VPWR VPWR _11193_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16568_ _08554_ _08624_ VGND VGND VPWR VPWR _08627_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18307_ _09675_ net3331 _10108_ VGND VGND VPWR VPWR _10158_ sky130_fd_sc_hd__mux2_1
X_15519_ _07525_ _07539_ _07591_ VGND VGND VPWR VPWR _07592_ sky130_fd_sc_hd__o21a_1
Xfanout8581 net8585 VGND VGND VPWR VPWR net8581 sky130_fd_sc_hd__dlymetal6s2s_1
X_19287_ net3197 net2526 _11123_ net3176 VGND VGND VPWR VPWR _11124_ sky130_fd_sc_hd__a211oi_1
X_16499_ _08555_ _08558_ VGND VGND VPWR VPWR _08559_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_183_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18238_ _10037_ net2564 VGND VGND VPWR VPWR _10089_ sky130_fd_sc_hd__nand2_1
Xfanout7880 net7899 VGND VGND VPWR VPWR net7880 sky130_fd_sc_hd__buf_1
X_18169_ _09840_ _09839_ VGND VGND VPWR VPWR _10020_ sky130_fd_sc_hd__or2_1
XFILLER_0_187_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20200_ _12022_ _12024_ VGND VGND VPWR VPWR _12025_ sky130_fd_sc_hd__and2b_1
XFILLER_0_142_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21180_ _01191_ _01195_ VGND VGND VPWR VPWR _01196_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20131_ _11844_ _11873_ VGND VGND VPWR VPWR _11959_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2709 net2710 VGND VGND VPWR VPWR net2709 sky130_fd_sc_hd__clkbuf_1
X_20062_ net3294 _11890_ VGND VGND VPWR VPWR _11891_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24870_ _04671_ VGND VGND VPWR VPWR _00733_ sky130_fd_sc_hd__clkbuf_1
X_23821_ _03600_ _03602_ VGND VGND VPWR VPWR _03686_ sky130_fd_sc_hd__nand2_1
X_23752_ net4703 net4828 VGND VGND VPWR VPWR _03618_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length7438 net7439 VGND VGND VPWR VPWR net7438 sky130_fd_sc_hd__buf_1
X_20964_ net5528 net5930 VGND VGND VPWR VPWR _00980_ sky130_fd_sc_hd__nand2_1
X_22703_ _02643_ net5459 net3095 VGND VGND VPWR VPWR _02644_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23683_ _03433_ _03434_ _03549_ VGND VGND VPWR VPWR _03550_ sky130_fd_sc_hd__a21oi_1
X_20895_ _00906_ _00910_ VGND VGND VPWR VPWR _00911_ sky130_fd_sc_hd__nand2_1
X_25422_ clknet_leaf_99_clk _00305_ net8382 VGND VGND VPWR VPWR matmul0.cos\[9\] sky130_fd_sc_hd__dfrtp_1
X_22634_ net5958 net3083 net2456 net8891 VGND VGND VPWR VPWR _00567_ sky130_fd_sc_hd__o211a_1
XFILLER_0_177_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25353_ clknet_leaf_83_clk _00236_ net8507 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult2\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_181_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22565_ net8987 net2043 _02548_ net7368 VGND VGND VPWR VPWR _00551_ sky130_fd_sc_hd__a22o_1
XFILLER_0_192_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24304_ net1013 net1656 _04163_ VGND VGND VPWR VPWR _04164_ sky130_fd_sc_hd__a21o_1
XFILLER_0_111_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21516_ _01418_ _01525_ VGND VGND VPWR VPWR _01529_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25284_ clknet_leaf_77_clk _00167_ net8440 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.c\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_145_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22496_ _02494_ _02496_ VGND VGND VPWR VPWR _02497_ sky130_fd_sc_hd__xnor2_1
Xwire6025 net6026 VGND VGND VPWR VPWR net6025 sky130_fd_sc_hd__buf_1
XFILLER_0_90_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6036 net6037 VGND VGND VPWR VPWR net6036 sky130_fd_sc_hd__buf_1
XFILLER_0_160_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24235_ _04088_ _04095_ VGND VGND VPWR VPWR _04096_ sky130_fd_sc_hd__xnor2_1
Xwire5302 net5303 VGND VGND VPWR VPWR net5302 sky130_fd_sc_hd__clkbuf_1
X_21447_ _01454_ _01459_ VGND VGND VPWR VPWR _01460_ sky130_fd_sc_hd__xor2_1
XFILLER_0_82_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout4517 net4528 VGND VGND VPWR VPWR net4517 sky130_fd_sc_hd__clkbuf_1
Xwire5313 matmul0.beta_pass\[0\] VGND VGND VPWR VPWR net5313 sky130_fd_sc_hd__buf_1
Xwire5324 net5325 VGND VGND VPWR VPWR net5324 sky130_fd_sc_hd__clkbuf_1
Xwire6069 net6071 VGND VGND VPWR VPWR net6069 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire5335 net5336 VGND VGND VPWR VPWR net5335 sky130_fd_sc_hd__clkbuf_1
Xwire4601 pid_q.mult0.a\[9\] VGND VGND VPWR VPWR net4601 sky130_fd_sc_hd__clkbuf_1
Xwire5346 net5347 VGND VGND VPWR VPWR net5346 sky130_fd_sc_hd__clkbuf_1
X_24166_ _04027_ VGND VGND VPWR VPWR _04028_ sky130_fd_sc_hd__inv_2
X_21378_ _01386_ _01391_ VGND VGND VPWR VPWR _01392_ sky130_fd_sc_hd__xnor2_1
Xwire5368 net5369 VGND VGND VPWR VPWR net5368 sky130_fd_sc_hd__clkbuf_1
Xwire4634 net4630 VGND VGND VPWR VPWR net4634 sky130_fd_sc_hd__buf_1
Xwire5379 net5374 VGND VGND VPWR VPWR net5379 sky130_fd_sc_hd__clkbuf_1
X_23117_ _02968_ net1677 VGND VGND VPWR VPWR _02987_ sky130_fd_sc_hd__nand2_1
X_20329_ net6479 net6472 net6466 _12084_ net3314 VGND VGND VPWR VPWR _12132_ sky130_fd_sc_hd__a2111o_1
Xwire3911 net3912 VGND VGND VPWR VPWR net3911 sky130_fd_sc_hd__clkbuf_1
Xwire4667 net4668 VGND VGND VPWR VPWR net4667 sky130_fd_sc_hd__buf_1
X_24097_ _03957_ _03958_ VGND VGND VPWR VPWR _03959_ sky130_fd_sc_hd__xnor2_1
Xwire3922 _10479_ VGND VGND VPWR VPWR net3922 sky130_fd_sc_hd__buf_1
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3933 _10094_ VGND VGND VPWR VPWR net3933 sky130_fd_sc_hd__clkbuf_1
Xwire4678 net4679 VGND VGND VPWR VPWR net4678 sky130_fd_sc_hd__clkbuf_1
Xwire4689 net4690 VGND VGND VPWR VPWR net4689 sky130_fd_sc_hd__clkbuf_1
Xwire3944 net3946 VGND VGND VPWR VPWR net3944 sky130_fd_sc_hd__clkbuf_1
X_23048_ _02913_ _02915_ _02917_ VGND VGND VPWR VPWR _02918_ sky130_fd_sc_hd__o21ba_1
Xwire3966 net3967 VGND VGND VPWR VPWR net3966 sky130_fd_sc_hd__buf_1
Xwire3977 net3978 VGND VGND VPWR VPWR net3977 sky130_fd_sc_hd__clkbuf_2
Xwire3988 net3989 VGND VGND VPWR VPWR net3988 sky130_fd_sc_hd__buf_1
Xwire3999 net4000 VGND VGND VPWR VPWR net3999 sky130_fd_sc_hd__clkbuf_1
X_15870_ _07937_ _07938_ VGND VGND VPWR VPWR _07939_ sky130_fd_sc_hd__xnor2_1
X_14821_ net7183 matmul0.matmul_stage_inst.e\[0\] net3630 VGND VGND VPWR VPWR _06927_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24999_ pid_q.out\[1\] net5181 VGND VGND VPWR VPWR _04756_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17540_ net6687 svm0.tC\[14\] VGND VGND VPWR VPWR _09422_ sky130_fd_sc_hd__and2b_1
X_14752_ net7448 net7155 VGND VGND VPWR VPWR _06884_ sky130_fd_sc_hd__nand2_1
X_13703_ net7647 VGND VGND VPWR VPWR _05972_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17471_ net3273 _09363_ net6661 VGND VGND VPWR VPWR _09364_ sky130_fd_sc_hd__o21a_1
X_14683_ net7161 net7165 net7159 net7157 VGND VGND VPWR VPWR _06832_ sky130_fd_sc_hd__or4_2
XFILLER_0_6_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19210_ net6276 net6218 VGND VGND VPWR VPWR _11047_ sky130_fd_sc_hd__nand2_1
XFILLER_0_196_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13634_ _05825_ _05826_ _05903_ VGND VGND VPWR VPWR _05904_ sky130_fd_sc_hd__a21o_1
X_16422_ _08381_ _08483_ _08428_ VGND VGND VPWR VPWR _08484_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_157_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout7110 net7114 VGND VGND VPWR VPWR net7110 sky130_fd_sc_hd__buf_1
XFILLER_0_26_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19141_ net6153 _10939_ _10976_ net3915 _10977_ VGND VGND VPWR VPWR _10978_ sky130_fd_sc_hd__a221oi_1
X_16353_ net3522 net2222 _08312_ _07936_ _08329_ VGND VGND VPWR VPWR _08416_ sky130_fd_sc_hd__o221a_1
X_13565_ _05728_ _05759_ _05727_ VGND VGND VPWR VPWR _05836_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_82_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout7143 cordic0.vec\[1\]\[0\] VGND VGND VPWR VPWR net7143 sky130_fd_sc_hd__buf_1
X_15304_ net4216 net4214 VGND VGND VPWR VPWR _07378_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19072_ _10862_ _10907_ _10908_ VGND VGND VPWR VPWR _10909_ sky130_fd_sc_hd__and3_1
X_16284_ _08347_ VGND VGND VPWR VPWR _08348_ sky130_fd_sc_hd__inv_2
X_13496_ net628 _05767_ _05768_ VGND VGND VPWR VPWR _05769_ sky130_fd_sc_hd__o21a_1
Xwire7260 net7261 VGND VGND VPWR VPWR net7260 sky130_fd_sc_hd__buf_1
X_18023_ _09872_ _09873_ VGND VGND VPWR VPWR _09874_ sky130_fd_sc_hd__xor2_1
X_15235_ net3551 VGND VGND VPWR VPWR _07309_ sky130_fd_sc_hd__clkbuf_1
Xwire7271 net7274 VGND VGND VPWR VPWR net7271 sky130_fd_sc_hd__buf_1
Xfanout6475 net6481 VGND VGND VPWR VPWR net6475 sky130_fd_sc_hd__buf_1
Xwire7282 net7283 VGND VGND VPWR VPWR net7282 sky130_fd_sc_hd__buf_1
XFILLER_0_152_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7293 matmul0.alpha_pass\[7\] VGND VGND VPWR VPWR net7293 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15166_ net3502 VGND VGND VPWR VPWR _07240_ sky130_fd_sc_hd__clkbuf_1
Xwire6581 net6580 VGND VGND VPWR VPWR net6581 sky130_fd_sc_hd__buf_1
Xfanout5774 net5778 VGND VGND VPWR VPWR net5774 sky130_fd_sc_hd__buf_1
X_14117_ net7666 net1314 VGND VGND VPWR VPWR _06379_ sky130_fd_sc_hd__nand2_1
Xwire5880 net5881 VGND VGND VPWR VPWR net5880 sky130_fd_sc_hd__buf_1
Xwire5891 net5892 VGND VGND VPWR VPWR net5891 sky130_fd_sc_hd__clkbuf_1
X_19974_ net6021 net3125 _11803_ _11804_ VGND VGND VPWR VPWR _11805_ sky130_fd_sc_hd__a211o_1
X_15097_ _07169_ _07170_ VGND VGND VPWR VPWR _07171_ sky130_fd_sc_hd__xnor2_1
X_14048_ _06253_ _06254_ VGND VGND VPWR VPWR _06312_ sky130_fd_sc_hd__and2b_1
X_18925_ _10742_ _10745_ _10741_ VGND VGND VPWR VPWR _10765_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18856_ net9085 net2288 net1449 _10698_ VGND VGND VPWR VPWR _00447_ sky130_fd_sc_hd__a31o_1
X_17807_ _09656_ _09657_ net7132 VGND VGND VPWR VPWR _09658_ sky130_fd_sc_hd__a21bo_1
X_18787_ _10584_ _10630_ VGND VGND VPWR VPWR _10631_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15999_ _07979_ net1094 _07977_ VGND VGND VPWR VPWR _08067_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17738_ net6454 _06541_ _09592_ VGND VGND VPWR VPWR _09593_ sky130_fd_sc_hd__or3_1
XFILLER_0_159_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17669_ _09544_ _09546_ _09547_ _09548_ VGND VGND VPWR VPWR _09549_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_175_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19408_ _11094_ _11045_ VGND VGND VPWR VPWR _11245_ sky130_fd_sc_hd__or2_1
X_20680_ net6091 _12445_ VGND VGND VPWR VPWR _12456_ sky130_fd_sc_hd__or2_1
XFILLER_0_175_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19339_ net3883 _10989_ _11175_ net6320 VGND VGND VPWR VPWR _11176_ sky130_fd_sc_hd__o31a_1
XFILLER_0_45_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3919 _10787_ VGND VGND VPWR VPWR net3919 sky130_fd_sc_hd__buf_1
X_22350_ net5438 net5670 VGND VGND VPWR VPWR _02353_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21301_ net5473 _12515_ _12516_ _00862_ VGND VGND VPWR VPWR _01316_ sky130_fd_sc_hd__o31a_1
XFILLER_0_60_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22281_ net5707 net5409 VGND VGND VPWR VPWR _02285_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24020_ _03879_ _03882_ VGND VGND VPWR VPWR _03883_ sky130_fd_sc_hd__xnor2_1
Xhold210 pid_q.out\[0\] VGND VGND VPWR VPWR net9163 sky130_fd_sc_hd__dlygate4sd3_1
X_21232_ net5987 net4392 VGND VGND VPWR VPWR _01247_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold221 pid_q.out\[6\] VGND VGND VPWR VPWR net9174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 pid_q.prev_int\[12\] VGND VGND VPWR VPWR net9185 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold243 pid_d.curr_int\[6\] VGND VGND VPWR VPWR net9196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 pid_q.prev_int\[3\] VGND VGND VPWR VPWR net9207 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3207 net3208 VGND VGND VPWR VPWR net3207 sky130_fd_sc_hd__clkbuf_1
X_21163_ _01149_ _01177_ _01178_ VGND VGND VPWR VPWR _01179_ sky130_fd_sc_hd__a21o_1
Xhold265 cordic0.slte0.opA\[4\] VGND VGND VPWR VPWR net9218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 pid_q.out\[7\] VGND VGND VPWR VPWR net9229 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3218 net3219 VGND VGND VPWR VPWR net3218 sky130_fd_sc_hd__clkbuf_1
Xhold287 cordic0.cos\[1\] VGND VGND VPWR VPWR net9240 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3229 _10104_ VGND VGND VPWR VPWR net3229 sky130_fd_sc_hd__clkbuf_2
X_20114_ net6107 net6042 VGND VGND VPWR VPWR _11942_ sky130_fd_sc_hd__or2_1
X_21094_ _01095_ _01109_ VGND VGND VPWR VPWR _01110_ sky130_fd_sc_hd__xnor2_1
Xwire2517 net2518 VGND VGND VPWR VPWR net2517 sky130_fd_sc_hd__clkbuf_1
Xwire2528 _10826_ VGND VGND VPWR VPWR net2528 sky130_fd_sc_hd__buf_1
Xwire2539 _10435_ VGND VGND VPWR VPWR net2539 sky130_fd_sc_hd__clkbuf_2
X_24922_ pid_q.ki\[3\] _04708_ net1362 VGND VGND VPWR VPWR _04709_ sky130_fd_sc_hd__mux2_1
Xwire1805 _08974_ VGND VGND VPWR VPWR net1805 sky130_fd_sc_hd__buf_1
X_20045_ _11844_ _11874_ VGND VGND VPWR VPWR _11875_ sky130_fd_sc_hd__xnor2_1
Xwire1816 net1817 VGND VGND VPWR VPWR net1816 sky130_fd_sc_hd__clkbuf_1
Xwire1827 _08904_ VGND VGND VPWR VPWR net1827 sky130_fd_sc_hd__buf_1
Xwire1838 net1839 VGND VGND VPWR VPWR net1838 sky130_fd_sc_hd__clkbuf_1
Xwire1849 _07901_ VGND VGND VPWR VPWR net1849 sky130_fd_sc_hd__buf_1
X_24853_ net7488 _04540_ net175 _04659_ VGND VGND VPWR VPWR _00728_ sky130_fd_sc_hd__a31o_1
X_23804_ pid_q.curr_int\[4\] net3062 net2028 _03669_ VGND VGND VPWR VPWR _00669_ sky130_fd_sc_hd__a22o_1
X_24784_ _04607_ _04610_ VGND VGND VPWR VPWR _04611_ sky130_fd_sc_hd__xnor2_1
X_21996_ _01999_ _02002_ _01998_ VGND VGND VPWR VPWR _02004_ sky130_fd_sc_hd__a21oi_2
Xmax_length7224 matmul0.alpha_pass\[13\] VGND VGND VPWR VPWR net7224 sky130_fd_sc_hd__buf_1
X_23735_ net4527 net5051 VGND VGND VPWR VPWR _03601_ sky130_fd_sc_hd__nand2_1
Xmax_length6523 net6521 VGND VGND VPWR VPWR net6523 sky130_fd_sc_hd__buf_1
X_20947_ _00956_ net1734 _00962_ VGND VGND VPWR VPWR _00963_ sky130_fd_sc_hd__a21oi_2
Xmax_length7279 net7280 VGND VGND VPWR VPWR net7279 sky130_fd_sc_hd__buf_1
Xmax_length5800 net5801 VGND VGND VPWR VPWR net5800 sky130_fd_sc_hd__buf_1
X_23666_ _03400_ _03401_ _03402_ VGND VGND VPWR VPWR _03533_ sky130_fd_sc_hd__o21a_1
X_20878_ net2486 net2485 VGND VGND VPWR VPWR _00894_ sky130_fd_sc_hd__xor2_1
XFILLER_0_76_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25405_ clknet_leaf_72_clk _00288_ net8469 VGND VGND VPWR VPWR matmul0.a\[8\] sky130_fd_sc_hd__dfrtp_1
X_22617_ net8888 _02588_ VGND VGND VPWR VPWR _02589_ sky130_fd_sc_hd__and2_1
X_23597_ net934 _03464_ _03376_ VGND VGND VPWR VPWR _03465_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_181_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13350_ _05613_ _05614_ _05621_ _05622_ VGND VGND VPWR VPWR _05623_ sky130_fd_sc_hd__o211a_1
X_25336_ clknet_leaf_84_clk _00219_ net8507 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_22548_ net9181 _02521_ _02536_ VGND VGND VPWR VPWR _00546_ sky130_fd_sc_hd__a21o_1
Xmax_length700 _01914_ VGND VGND VPWR VPWR net700 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13281_ net918 _05429_ _05428_ VGND VGND VPWR VPWR _05554_ sky130_fd_sc_hd__a21oi_2
X_25267_ clknet_leaf_77_clk _00150_ net8440 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.b\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_22479_ net5377 _02479_ VGND VGND VPWR VPWR _02480_ sky130_fd_sc_hd__nand2_1
Xwire5110 net5103 VGND VGND VPWR VPWR net5110 sky130_fd_sc_hd__buf_1
Xwire5121 net5122 VGND VGND VPWR VPWR net5121 sky130_fd_sc_hd__buf_1
Xfanout4314 net4322 VGND VGND VPWR VPWR net4314 sky130_fd_sc_hd__clkbuf_1
X_15020_ _07085_ _07091_ _07093_ VGND VGND VPWR VPWR _07094_ sky130_fd_sc_hd__a21o_1
X_24218_ net4484 _04078_ VGND VGND VPWR VPWR _04079_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5132 net5133 VGND VGND VPWR VPWR net5132 sky130_fd_sc_hd__buf_1
XFILLER_0_20_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5143 net5144 VGND VGND VPWR VPWR net5143 sky130_fd_sc_hd__buf_1
XFILLER_0_20_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25198_ clknet_leaf_73_clk _00087_ net8474 VGND VGND VPWR VPWR matmul0.b_in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire5154 net5155 VGND VGND VPWR VPWR net5154 sky130_fd_sc_hd__buf_1
Xwire5165 net5156 VGND VGND VPWR VPWR net5165 sky130_fd_sc_hd__buf_1
Xwire4420 net4421 VGND VGND VPWR VPWR net4420 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4431 net4432 VGND VGND VPWR VPWR net4431 sky130_fd_sc_hd__clkbuf_1
X_24149_ _03903_ _04008_ net2023 VGND VGND VPWR VPWR _04011_ sky130_fd_sc_hd__o21a_1
Xwire5176 net5177 VGND VGND VPWR VPWR net5176 sky130_fd_sc_hd__buf_1
Xwire5187 net5188 VGND VGND VPWR VPWR net5187 sky130_fd_sc_hd__clkbuf_1
Xwire4442 pid_q.out\[7\] VGND VGND VPWR VPWR net4442 sky130_fd_sc_hd__clkbuf_1
Xwire5198 net5200 VGND VGND VPWR VPWR net5198 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4453 net4454 VGND VGND VPWR VPWR net4453 sky130_fd_sc_hd__clkbuf_1
Xwire4464 net4465 VGND VGND VPWR VPWR net4464 sky130_fd_sc_hd__clkbuf_1
Xwire4475 pid_q.kp\[15\] VGND VGND VPWR VPWR net4475 sky130_fd_sc_hd__clkbuf_1
Xwire3741 net3742 VGND VGND VPWR VPWR net3741 sky130_fd_sc_hd__buf_1
Xwire3752 _03065_ VGND VGND VPWR VPWR net3752 sky130_fd_sc_hd__buf_1
X_16971_ _08838_ net2612 net1808 VGND VGND VPWR VPWR _08934_ sky130_fd_sc_hd__o21a_1
Xwire4497 net4492 VGND VGND VPWR VPWR net4497 sky130_fd_sc_hd__clkbuf_1
Xwire3763 _02712_ VGND VGND VPWR VPWR net3763 sky130_fd_sc_hd__clkbuf_1
Xwire3774 _02541_ VGND VGND VPWR VPWR net3774 sky130_fd_sc_hd__buf_1
X_18710_ _10485_ _10491_ VGND VGND VPWR VPWR _10556_ sky130_fd_sc_hd__nand2_1
Xwire3785 net3787 VGND VGND VPWR VPWR net3785 sky130_fd_sc_hd__clkbuf_1
X_15922_ net2829 net2846 _07898_ net2212 net2836 VGND VGND VPWR VPWR _07991_ sky130_fd_sc_hd__a32o_1
X_19690_ net1415 _11525_ VGND VGND VPWR VPWR _11526_ sky130_fd_sc_hd__xnor2_1
Xwire3796 net3797 VGND VGND VPWR VPWR net3796 sky130_fd_sc_hd__buf_1
XFILLER_0_36_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18641_ net6792 net6769 net2539 VGND VGND VPWR VPWR _10488_ sky130_fd_sc_hd__mux2_1
X_15853_ matmul0.matmul_stage_inst.mult1\[4\] net396 net2680 VGND VGND VPWR VPWR _07923_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14804_ net3625 matmul0.cos\[6\] _06802_ net2855 VGND VGND VPWR VPWR _06919_ sky130_fd_sc_hd__o211a_1
X_18572_ net1197 _10377_ _10378_ VGND VGND VPWR VPWR _10420_ sky130_fd_sc_hd__o21ai_1
X_12996_ _05265_ _05268_ VGND VGND VPWR VPWR _05269_ sky130_fd_sc_hd__xnor2_2
X_15784_ _07752_ _07753_ _07853_ VGND VGND VPWR VPWR _07854_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17523_ net6694 _09272_ VGND VGND VPWR VPWR _09408_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14735_ net9071 net2860 _06867_ _06870_ VGND VGND VPWR VPWR _00153_ sky130_fd_sc_hd__a22o_1
X_17454_ _09347_ _09348_ VGND VGND VPWR VPWR _09349_ sky130_fd_sc_hd__nand2_1
X_14666_ net3625 net7166 net2876 VGND VGND VPWR VPWR _06819_ sky130_fd_sc_hd__o21a_1
XFILLER_0_86_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13617_ _05881_ _05886_ VGND VGND VPWR VPWR _05887_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16405_ net882 _08405_ _08406_ VGND VGND VPWR VPWR _08467_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_67_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17385_ net612 _09293_ _09291_ VGND VGND VPWR VPWR _09294_ sky130_fd_sc_hd__a21oi_1
X_14597_ net7214 net5200 _06769_ VGND VGND VPWR VPWR _06771_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_138_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19124_ net6119 net6155 VGND VGND VPWR VPWR _10961_ sky130_fd_sc_hd__nand2_1
X_13548_ _05814_ _05815_ _05816_ _05817_ VGND VGND VPWR VPWR _05819_ sky130_fd_sc_hd__o22a_1
XFILLER_0_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16336_ _08393_ _08398_ VGND VGND VPWR VPWR _08399_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6250 net6256 VGND VGND VPWR VPWR net6250 sky130_fd_sc_hd__clkbuf_1
Xfanout6261 net6282 VGND VGND VPWR VPWR net6261 sky130_fd_sc_hd__clkbuf_2
X_19055_ _10884_ _10886_ _10890_ VGND VGND VPWR VPWR _10892_ sky130_fd_sc_hd__and3_1
X_16267_ _08329_ _08330_ VGND VGND VPWR VPWR _08331_ sky130_fd_sc_hd__and2_1
X_13479_ net7640 net2350 net2346 VGND VGND VPWR VPWR _05752_ sky130_fd_sc_hd__and3_1
XFILLER_0_125_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18006_ net3257 _09615_ VGND VGND VPWR VPWR _09857_ sky130_fd_sc_hd__nand2_1
X_15218_ net1881 net1880 _07291_ VGND VGND VPWR VPWR _07292_ sky130_fd_sc_hd__a21o_1
X_16198_ net2840 net3394 _08170_ net2670 VGND VGND VPWR VPWR _08263_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15149_ _07221_ _07222_ VGND VGND VPWR VPWR _07223_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_11_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19957_ net1409 _11766_ _11787_ VGND VGND VPWR VPWR _11788_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_96_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18908_ net6376 _10747_ net275 VGND VGND VPWR VPWR _10749_ sky130_fd_sc_hd__a21bo_1
X_19888_ _11667_ net708 VGND VGND VPWR VPWR _11721_ sky130_fd_sc_hd__and2_1
XFILLER_0_184_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18839_ net1428 _10681_ VGND VGND VPWR VPWR _10682_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_171_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21850_ net2475 _01787_ net2064 VGND VGND VPWR VPWR _01859_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20801_ _00810_ _00816_ _12536_ VGND VGND VPWR VPWR _00817_ sky130_fd_sc_hd__o21ai_1
X_21781_ _01788_ _01790_ VGND VGND VPWR VPWR _01791_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23520_ net7526 _03317_ net540 net7466 net2417 VGND VGND VPWR VPWR _03389_ sky130_fd_sc_hd__a221o_1
X_20732_ net2487 VGND VGND VPWR VPWR _12503_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8719 net8720 VGND VGND VPWR VPWR net8719 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_186_Right_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23451_ _03282_ _03293_ net1385 VGND VGND VPWR VPWR _03320_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_122_Left_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20663_ net6502 net3325 net3850 VGND VGND VPWR VPWR _12440_ sky130_fd_sc_hd__or3_1
XFILLER_0_135_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire409 _03761_ VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__clkbuf_1
X_22402_ pid_d.prev_error\[14\] pid_d.curr_error\[14\] VGND VGND VPWR VPWR _02404_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_46_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length3716 _04869_ VGND VGND VPWR VPWR net3716 sky130_fd_sc_hd__clkbuf_1
X_23382_ _03247_ _03250_ VGND VGND VPWR VPWR _03252_ sky130_fd_sc_hd__nand2_1
X_20594_ net3124 _12314_ _09004_ VGND VGND VPWR VPWR _12376_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25121_ net9205 _04850_ _04853_ net5976 VGND VGND VPWR VPWR _00802_ sky130_fd_sc_hd__a22o_1
X_22333_ _02332_ _02335_ VGND VGND VPWR VPWR _02336_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_190_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25052_ net3737 net685 VGND VGND VPWR VPWR _04802_ sky130_fd_sc_hd__xnor2_1
X_22264_ _02264_ _02267_ VGND VGND VPWR VPWR _02268_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24003_ _03778_ _03847_ _03849_ VGND VGND VPWR VPWR _03866_ sky130_fd_sc_hd__a21oi_1
X_21215_ _01027_ _01222_ net861 VGND VGND VPWR VPWR _01231_ sky130_fd_sc_hd__o21a_1
X_22195_ net1712 _02152_ net1169 VGND VGND VPWR VPWR _02200_ sky130_fd_sc_hd__a21o_1
Xwire3004 net3005 VGND VGND VPWR VPWR net3004 sky130_fd_sc_hd__buf_1
Xwire3015 net3018 VGND VGND VPWR VPWR net3015 sky130_fd_sc_hd__clkbuf_1
Xwire3026 _04870_ VGND VGND VPWR VPWR net3026 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3037 net3038 VGND VGND VPWR VPWR net3037 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_131_Left_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21146_ net5605 net5880 VGND VGND VPWR VPWR _01162_ sky130_fd_sc_hd__nand2_1
Xwire3048 _03739_ VGND VGND VPWR VPWR net3048 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2303 _05348_ VGND VGND VPWR VPWR net2303 sky130_fd_sc_hd__buf_1
Xwire3059 _03198_ VGND VGND VPWR VPWR net3059 sky130_fd_sc_hd__buf_1
Xwire2314 net2315 VGND VGND VPWR VPWR net2314 sky130_fd_sc_hd__clkbuf_1
Xwire2325 net2326 VGND VGND VPWR VPWR net2325 sky130_fd_sc_hd__buf_1
Xwire2336 net2337 VGND VGND VPWR VPWR net2336 sky130_fd_sc_hd__buf_1
Xwire1602 net1603 VGND VGND VPWR VPWR net1602 sky130_fd_sc_hd__buf_1
Xwire2347 net2348 VGND VGND VPWR VPWR net2347 sky130_fd_sc_hd__buf_1
X_21077_ net5581 _01092_ VGND VGND VPWR VPWR _01093_ sky130_fd_sc_hd__and2_1
Xwire1613 net1614 VGND VGND VPWR VPWR net1613 sky130_fd_sc_hd__clkbuf_1
Xwire2358 _04910_ VGND VGND VPWR VPWR net2358 sky130_fd_sc_hd__clkbuf_1
Xwire1624 net1625 VGND VGND VPWR VPWR net1624 sky130_fd_sc_hd__buf_1
Xwire2369 net2370 VGND VGND VPWR VPWR net2369 sky130_fd_sc_hd__clkbuf_1
Xwire1635 _04734_ VGND VGND VPWR VPWR net1635 sky130_fd_sc_hd__buf_1
X_24905_ net129 net8885 net116 net119 VGND VGND VPWR VPWR _04695_ sky130_fd_sc_hd__or4_1
Xwire1646 _04509_ VGND VGND VPWR VPWR net1646 sky130_fd_sc_hd__buf_1
X_20028_ net3147 net6062 net3144 VGND VGND VPWR VPWR _11858_ sky130_fd_sc_hd__or3_1
X_25885_ clknet_leaf_18_clk _00758_ net8630 VGND VGND VPWR VPWR pid_q.ki\[13\] sky130_fd_sc_hd__dfrtp_1
Xwire1657 _04085_ VGND VGND VPWR VPWR net1657 sky130_fd_sc_hd__buf_1
Xwire1668 net1669 VGND VGND VPWR VPWR net1668 sky130_fd_sc_hd__clkbuf_1
Xwire1679 net1680 VGND VGND VPWR VPWR net1679 sky130_fd_sc_hd__dlymetal6s2s_1
X_12850_ _05102_ _05122_ VGND VGND VPWR VPWR _05123_ sky130_fd_sc_hd__xnor2_1
X_24836_ net7481 net737 _03952_ VGND VGND VPWR VPWR _04651_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length7021 net7022 VGND VGND VPWR VPWR net7021 sky130_fd_sc_hd__buf_1
XFILLER_0_68_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24767_ pid_q.curr_error\[9\] net1370 net1367 net629 VGND VGND VPWR VPWR _00706_
+ sky130_fd_sc_hd__a22o_1
X_12781_ svm0.vC\[8\] _04889_ VGND VGND VPWR VPWR _05054_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21979_ _01880_ _01881_ _01878_ VGND VGND VPWR VPWR _01987_ sky130_fd_sc_hd__mux2_1
X_14520_ _06692_ _06694_ net5262 VGND VGND VPWR VPWR _06700_ sky130_fd_sc_hd__a21o_1
X_23718_ net696 _03470_ _03472_ _03583_ VGND VGND VPWR VPWR _03584_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_140_Left_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24698_ pid_q.curr_error\[0\] net1370 _04533_ net2015 VGND VGND VPWR VPWR _00697_
+ sky130_fd_sc_hd__a22o_1
Xmax_length7098 net7099 VGND VGND VPWR VPWR net7098 sky130_fd_sc_hd__buf_1
XFILLER_0_127_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14451_ _06642_ VGND VGND VPWR VPWR _00097_ sky130_fd_sc_hd__clkbuf_1
Xmax_length5641 net5643 VGND VGND VPWR VPWR net5641 sky130_fd_sc_hd__buf_1
X_23649_ _03512_ _03515_ VGND VGND VPWR VPWR _03516_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_166_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_153_Right_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13402_ _05563_ _05486_ _05481_ _05405_ VGND VGND VPWR VPWR _05675_ sky130_fd_sc_hd__o2bb2a_1
Xmax_length5674 net5673 VGND VGND VPWR VPWR net5674 sky130_fd_sc_hd__buf_1
XFILLER_0_25_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17170_ net5997 net3361 _09096_ VGND VGND VPWR VPWR _09122_ sky130_fd_sc_hd__mux2_1
Xwire910 _05964_ VGND VGND VPWR VPWR net910 sky130_fd_sc_hd__clkbuf_1
X_14382_ _06589_ net7584 net899 VGND VGND VPWR VPWR _06590_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire921 _05299_ VGND VGND VPWR VPWR net921 sky130_fd_sc_hd__clkbuf_1
Xwire932 _03828_ VGND VGND VPWR VPWR net932 sky130_fd_sc_hd__buf_1
X_16121_ net2752 net3435 VGND VGND VPWR VPWR _08187_ sky130_fd_sc_hd__nor2_1
X_13333_ net7827 net1590 VGND VGND VPWR VPWR _05606_ sky130_fd_sc_hd__nand2_1
Xwire943 _02239_ VGND VGND VPWR VPWR net943 sky130_fd_sc_hd__buf_1
XFILLER_0_109_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25319_ clknet_leaf_78_clk _00202_ net8439 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.f\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire954 net955 VGND VGND VPWR VPWR net954 sky130_fd_sc_hd__clkbuf_1
Xwire965 _09464_ VGND VGND VPWR VPWR net965 sky130_fd_sc_hd__clkbuf_1
Xwire976 net977 VGND VGND VPWR VPWR net976 sky130_fd_sc_hd__buf_2
X_16052_ _08019_ _08020_ _08021_ VGND VGND VPWR VPWR _08119_ sky130_fd_sc_hd__a21o_1
Xwire987 _07833_ VGND VGND VPWR VPWR net987 sky130_fd_sc_hd__buf_1
Xwire998 _05735_ VGND VGND VPWR VPWR net998 sky130_fd_sc_hd__buf_1
X_13264_ net1330 _05536_ VGND VGND VPWR VPWR _05537_ sky130_fd_sc_hd__xor2_1
Xmax_length585 _05317_ VGND VGND VPWR VPWR net585 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15003_ net3584 net3577 VGND VGND VPWR VPWR _07077_ sky130_fd_sc_hd__or2_1
X_13195_ _05382_ net849 _05379_ VGND VGND VPWR VPWR _05468_ sky130_fd_sc_hd__a21oi_1
X_19811_ net6121 net3913 VGND VGND VPWR VPWR _11645_ sky130_fd_sc_hd__nand2_1
Xwire4261 net4262 VGND VGND VPWR VPWR net4261 sky130_fd_sc_hd__buf_1
Xwire4272 net4273 VGND VGND VPWR VPWR net4272 sky130_fd_sc_hd__buf_1
Xwire4283 net4284 VGND VGND VPWR VPWR net4283 sky130_fd_sc_hd__buf_1
Xwire4294 net4295 VGND VGND VPWR VPWR net4294 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19742_ _11518_ _11522_ net3157 VGND VGND VPWR VPWR _11577_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_21_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16954_ net1495 VGND VGND VPWR VPWR _08917_ sky130_fd_sc_hd__clkbuf_1
Xwire3582 net3583 VGND VGND VPWR VPWR net3582 sky130_fd_sc_hd__buf_1
Xwire3593 _06985_ VGND VGND VPWR VPWR net3593 sky130_fd_sc_hd__buf_1
XFILLER_0_194_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15905_ net3546 net3392 _07971_ _07972_ VGND VGND VPWR VPWR _07974_ sky130_fd_sc_hd__o211ai_1
Xwire2881 _06719_ VGND VGND VPWR VPWR net2881 sky130_fd_sc_hd__buf_1
X_19673_ net6030 _11508_ VGND VGND VPWR VPWR _11509_ sky130_fd_sc_hd__xnor2_1
X_16885_ net3362 _08845_ _08847_ net4056 _08825_ net4059 VGND VGND VPWR VPWR _08849_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_95_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18624_ net7016 _10467_ _10470_ VGND VGND VPWR VPWR _10471_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15836_ _07892_ _07905_ VGND VGND VPWR VPWR _07906_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18555_ net9088 net2289 _09598_ _10403_ VGND VGND VPWR VPWR _00441_ sky130_fd_sc_hd__a31o_1
X_12979_ _05250_ _05251_ VGND VGND VPWR VPWR _05252_ sky130_fd_sc_hd__xor2_1
X_15767_ _07834_ _07836_ VGND VGND VPWR VPWR _07837_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_86_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17506_ _09392_ VGND VGND VPWR VPWR _09393_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14718_ matmul0.sin\[12\] _06855_ VGND VGND VPWR VPWR _06858_ sky130_fd_sc_hd__or2_1
X_18486_ net3923 net607 VGND VGND VPWR VPWR _10336_ sky130_fd_sc_hd__nor2_1
X_15698_ net2720 net3414 VGND VGND VPWR VPWR _07769_ sky130_fd_sc_hd__nor2_1
X_17437_ net4035 net7376 net2570 _09334_ VGND VGND VPWR VPWR _00391_ sky130_fd_sc_hd__a31o_1
XFILLER_0_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14649_ net7437 matmul0.cos\[6\] net2875 VGND VGND VPWR VPWR _06809_ sky130_fd_sc_hd__and3_1
XFILLER_0_170_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_120_Right_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17368_ _09277_ _09279_ svm0.delta\[2\] VGND VGND VPWR VPWR _09280_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19107_ net6272 net6241 VGND VGND VPWR VPWR _10944_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16319_ net2815 net1250 net2648 VGND VGND VPWR VPWR _08382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_121_clk clknet_4_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_121_clk
+ sky130_fd_sc_hd__clkbuf_16
X_17299_ net7682 _09212_ VGND VGND VPWR VPWR _09213_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6080 cordic0.vec\[0\]\[13\] VGND VGND VPWR VPWR net6080 sky130_fd_sc_hd__buf_1
XFILLER_0_42_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19038_ net6260 net6245 VGND VGND VPWR VPWR _10875_ sky130_fd_sc_hd__and2b_1
Xfanout6091 net6104 VGND VGND VPWR VPWR net6091 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_113_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21000_ _00998_ _01002_ VGND VGND VPWR VPWR _01016_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22951_ net336 _02324_ VGND VGND VPWR VPWR _02839_ sky130_fd_sc_hd__nand2_1
XFILLER_0_173_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21902_ pid_d.prev_error\[7\] pid_d.curr_error\[7\] VGND VGND VPWR VPWR _01911_ sky130_fd_sc_hd__xnor2_1
X_25670_ clknet_leaf_5_clk _00543_ net8565 VGND VGND VPWR VPWR pid_d.prev_error\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_22882_ net5357 net3103 VGND VGND VPWR VPWR _02777_ sky130_fd_sc_hd__nor2_1
XFILLER_0_168_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24621_ net4539 _04475_ _04424_ net4514 VGND VGND VPWR VPWR _04476_ sky130_fd_sc_hd__o31a_1
X_21833_ _01836_ _01841_ VGND VGND VPWR VPWR _01842_ sky130_fd_sc_hd__xor2_1
XFILLER_0_195_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24552_ _04405_ _04407_ VGND VGND VPWR VPWR _04408_ sky130_fd_sc_hd__nor2_1
X_21764_ _01770_ _01773_ VGND VGND VPWR VPWR _01774_ sky130_fd_sc_hd__xor2_1
XFILLER_0_182_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23503_ net4842 net4827 VGND VGND VPWR VPWR _03372_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20715_ net6023 _12486_ _12487_ VGND VGND VPWR VPWR _00517_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_176_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24483_ net4485 _04202_ _04288_ VGND VGND VPWR VPWR _04340_ sky130_fd_sc_hd__o21ai_1
Xwire8516 net8510 VGND VGND VPWR VPWR net8516 sky130_fd_sc_hd__clkbuf_1
X_21695_ _01698_ _01705_ VGND VGND VPWR VPWR _01706_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_93_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8527 net8528 VGND VGND VPWR VPWR net8527 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8538 net8539 VGND VGND VPWR VPWR net8538 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7804 net7800 VGND VGND VPWR VPWR net7804 sky130_fd_sc_hd__clkbuf_2
Xwire8549 net8550 VGND VGND VPWR VPWR net8549 sky130_fd_sc_hd__clkbuf_1
X_23434_ net1166 net938 VGND VGND VPWR VPWR _03304_ sky130_fd_sc_hd__xnor2_1
Xwire7815 net7816 VGND VGND VPWR VPWR net7815 sky130_fd_sc_hd__buf_1
Xmax_length4247 _06499_ VGND VGND VPWR VPWR net4247 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4258 _05127_ VGND VGND VPWR VPWR net4258 sky130_fd_sc_hd__clkbuf_1
Xwire206 _02407_ VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_1
X_20646_ net1239 _12423_ net3147 VGND VGND VPWR VPWR _12425_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3513 _07095_ VGND VGND VPWR VPWR net3513 sky130_fd_sc_hd__buf_1
XFILLER_0_92_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire217 _06364_ VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__clkbuf_2
Xwire7826 net7820 VGND VGND VPWR VPWR net7826 sky130_fd_sc_hd__buf_1
Xwire7837 net7840 VGND VGND VPWR VPWR net7837 sky130_fd_sc_hd__clkbuf_1
Xwire228 net229 VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__clkbuf_1
Xwire239 net240 VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__clkbuf_1
Xwire7848 net7849 VGND VGND VPWR VPWR net7848 sky130_fd_sc_hd__buf_1
XFILLER_0_61_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7859 net7856 VGND VGND VPWR VPWR net7859 sky130_fd_sc_hd__clkbuf_1
X_23365_ _03232_ _03234_ VGND VGND VPWR VPWR _03235_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length2812 net2813 VGND VGND VPWR VPWR net2812 sky130_fd_sc_hd__buf_1
X_20577_ net6253 net1492 _12359_ VGND VGND VPWR VPWR _12361_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_112_clk clknet_4_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_112_clk
+ sky130_fd_sc_hd__clkbuf_16
X_25104_ _04845_ _04846_ VGND VGND VPWR VPWR _04847_ sky130_fd_sc_hd__xnor2_1
X_22316_ _02237_ _02240_ _02319_ VGND VGND VPWR VPWR _02320_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length2845 _07016_ VGND VGND VPWR VPWR net2845 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2856 _06869_ VGND VGND VPWR VPWR net2856 sky130_fd_sc_hd__clkbuf_1
X_23296_ _03145_ _03158_ _03159_ _03165_ VGND VGND VPWR VPWR _03166_ sky130_fd_sc_hd__a211o_1
XFILLER_0_108_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2878 _06802_ VGND VGND VPWR VPWR net2878 sky130_fd_sc_hd__buf_1
XFILLER_0_42_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25035_ pid_q.out\[5\] _04783_ net1995 VGND VGND VPWR VPWR _04788_ sky130_fd_sc_hd__nor3_1
X_22247_ _02115_ _02169_ _02170_ VGND VGND VPWR VPWR _02252_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_44_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22178_ pid_d.curr_int\[10\] VGND VGND VPWR VPWR _02183_ sky130_fd_sc_hd__inv_2
Xwire2100 _11586_ VGND VGND VPWR VPWR net2100 sky130_fd_sc_hd__clkbuf_2
Xwire2111 _10952_ VGND VGND VPWR VPWR net2111 sky130_fd_sc_hd__buf_1
X_21129_ _01104_ _01111_ _01110_ VGND VGND VPWR VPWR _01145_ sky130_fd_sc_hd__and3_1
Xwire2133 net2134 VGND VGND VPWR VPWR net2133 sky130_fd_sc_hd__buf_1
Xwire2144 _09698_ VGND VGND VPWR VPWR net2144 sky130_fd_sc_hd__clkbuf_1
Xwire2155 _09429_ VGND VGND VPWR VPWR net2155 sky130_fd_sc_hd__buf_1
XFILLER_0_108_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1410 net1411 VGND VGND VPWR VPWR net1410 sky130_fd_sc_hd__buf_1
Xwire2166 net2167 VGND VGND VPWR VPWR net2166 sky130_fd_sc_hd__buf_1
Xwire1421 _11173_ VGND VGND VPWR VPWR net1421 sky130_fd_sc_hd__buf_1
X_13951_ net9118 net1126 net220 net1926 VGND VGND VPWR VPWR _00023_ sky130_fd_sc_hd__a22o_1
X_25937_ clknet_leaf_25_clk _00002_ net8581 VGND VGND VPWR VPWR pid_d.state\[1\] sky130_fd_sc_hd__dfrtp_1
Xwire2177 _08851_ VGND VGND VPWR VPWR net2177 sky130_fd_sc_hd__clkbuf_2
Xwire1432 _10477_ VGND VGND VPWR VPWR net1432 sky130_fd_sc_hd__clkbuf_1
Xwire1443 _10261_ VGND VGND VPWR VPWR net1443 sky130_fd_sc_hd__buf_1
Xwire1454 _09584_ VGND VGND VPWR VPWR net1454 sky130_fd_sc_hd__buf_1
Xwire2199 net2200 VGND VGND VPWR VPWR net2199 sky130_fd_sc_hd__buf_1
X_12902_ net7759 net1617 _05095_ _05096_ VGND VGND VPWR VPWR _05175_ sky130_fd_sc_hd__a22o_1
Xwire1476 net1477 VGND VGND VPWR VPWR net1476 sky130_fd_sc_hd__dlymetal6s2s_1
X_13882_ net283 _06148_ VGND VGND VPWR VPWR _06149_ sky130_fd_sc_hd__nand2_1
X_16670_ _08703_ VGND VGND VPWR VPWR _00255_ sky130_fd_sc_hd__clkbuf_1
X_25868_ clknet_leaf_17_clk _00741_ net8624 VGND VGND VPWR VPWR pid_q.mult0.a\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1487 net1488 VGND VGND VPWR VPWR net1487 sky130_fd_sc_hd__clkbuf_1
X_12833_ _05104_ _05105_ VGND VGND VPWR VPWR _05106_ sky130_fd_sc_hd__xnor2_1
X_15621_ net2851 _07692_ _07605_ VGND VGND VPWR VPWR _07693_ sky130_fd_sc_hd__a21o_1
X_24819_ net2403 VGND VGND VPWR VPWR _04641_ sky130_fd_sc_hd__clkbuf_1
X_25799_ clknet_leaf_29_clk _00672_ net8678 VGND VGND VPWR VPWR pid_q.curr_int\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18340_ _10189_ _10190_ VGND VGND VPWR VPWR _10191_ sky130_fd_sc_hd__xor2_1
X_12764_ _05034_ _05036_ VGND VGND VPWR VPWR _05037_ sky130_fd_sc_hd__xor2_1
X_15552_ net1270 _07624_ VGND VGND VPWR VPWR _07625_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_84_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14503_ _06679_ _06681_ _06684_ VGND VGND VPWR VPWR _06685_ sky130_fd_sc_hd__a21o_1
X_15483_ _07341_ _07471_ _07472_ VGND VGND VPWR VPWR _07557_ sky130_fd_sc_hd__a21o_1
X_18271_ net6760 VGND VGND VPWR VPWR _10122_ sky130_fd_sc_hd__inv_2
XFILLER_0_166_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12695_ _04950_ _04951_ _04949_ VGND VGND VPWR VPWR _04968_ sky130_fd_sc_hd__a21o_1
Xmax_length6183 net6184 VGND VGND VPWR VPWR net6183 sky130_fd_sc_hd__buf_1
XFILLER_0_12_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length5460 net5461 VGND VGND VPWR VPWR net5460 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17222_ net3290 VGND VGND VPWR VPWR _09170_ sky130_fd_sc_hd__buf_1
X_14434_ _06629_ matmul0.b_in\[10\] net896 VGND VGND VPWR VPWR _06630_ sky130_fd_sc_hd__mux2_1
Xinput14 angle_in[7] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_1
Xwire740 _04018_ VGND VGND VPWR VPWR net740 sky130_fd_sc_hd__clkbuf_1
X_14365_ net7259 _06574_ _06569_ net5346 _06576_ VGND VGND VPWR VPWR _06577_ sky130_fd_sc_hd__a221o_1
Xinput25 currA_in[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
X_17153_ _09102_ net527 VGND VGND VPWR VPWR _09107_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_103_clk clknet_4_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_103_clk
+ sky130_fd_sc_hd__clkbuf_16
Xinput36 currB_in[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
Xwire751 net752 VGND VGND VPWR VPWR net751 sky130_fd_sc_hd__clkbuf_1
Xinput47 currB_in[8] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_1
Xwire762 _01216_ VGND VGND VPWR VPWR net762 sky130_fd_sc_hd__clkbuf_1
Xinput58 currT_in[3] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_1
X_13316_ net1131 _05588_ VGND VGND VPWR VPWR _05589_ sky130_fd_sc_hd__xnor2_1
X_16104_ net2648 net3418 VGND VGND VPWR VPWR _08170_ sky130_fd_sc_hd__nor2_2
Xwire773 _08426_ VGND VGND VPWR VPWR net773 sky130_fd_sc_hd__buf_1
Xwire784 _05844_ VGND VGND VPWR VPWR net784 sky130_fd_sc_hd__clkbuf_1
Xinput69 periodTop[13] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_1
X_17084_ _09040_ _09041_ VGND VGND VPWR VPWR _09042_ sky130_fd_sc_hd__nand2b_1
Xwire795 _03781_ VGND VGND VPWR VPWR net795 sky130_fd_sc_hd__buf_1
X_14296_ net70 net3649 net2915 net7634 VGND VGND VPWR VPWR _00065_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13247_ _05519_ VGND VGND VPWR VPWR _05520_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16035_ _08038_ _08039_ _08041_ VGND VGND VPWR VPWR _08102_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13178_ net7714 net1976 net2312 VGND VGND VPWR VPWR _05451_ sky130_fd_sc_hd__and3_1
Xwire4080 _07572_ VGND VGND VPWR VPWR net4080 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_196_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4091 _07370_ VGND VGND VPWR VPWR net4091 sky130_fd_sc_hd__clkbuf_1
X_17986_ _09834_ _09836_ net1215 VGND VGND VPWR VPWR _09837_ sky130_fd_sc_hd__a21boi_1
Xwire3390 net3391 VGND VGND VPWR VPWR net3390 sky130_fd_sc_hd__dlymetal6s2s_1
X_19725_ net3856 VGND VGND VPWR VPWR _11560_ sky130_fd_sc_hd__inv_2
X_16937_ net6393 cordic0.slte0.opA\[14\] VGND VGND VPWR VPWR _08901_ sky130_fd_sc_hd__and2b_1
XFILLER_0_74_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19656_ _11454_ _11456_ VGND VGND VPWR VPWR _11492_ sky130_fd_sc_hd__nor2_1
X_16868_ net3364 _08831_ net4059 VGND VGND VPWR VPWR _08833_ sky130_fd_sc_hd__mux2_1
X_18607_ _10453_ _10454_ VGND VGND VPWR VPWR _10455_ sky130_fd_sc_hd__or2_1
X_15819_ _07862_ _07888_ VGND VGND VPWR VPWR _07889_ sky130_fd_sc_hd__xnor2_1
X_19587_ _11363_ _11370_ _11371_ _11423_ VGND VGND VPWR VPWR _11424_ sky130_fd_sc_hd__o31a_1
X_16799_ _08789_ VGND VGND VPWR VPWR _00298_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18538_ net3225 VGND VGND VPWR VPWR _10387_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18469_ net3284 net3225 VGND VGND VPWR VPWR _10319_ sky130_fd_sc_hd__nand2_1
XFILLER_0_185_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20500_ net2086 VGND VGND VPWR VPWR _12287_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21480_ _01491_ _01492_ VGND VGND VPWR VPWR _01493_ sky130_fd_sc_hd__xor2_2
XFILLER_0_28_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20431_ net950 _12224_ _12225_ VGND VGND VPWR VPWR _12226_ sky130_fd_sc_hd__mux2_2
XFILLER_0_172_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5709 net5710 VGND VGND VPWR VPWR net5709 sky130_fd_sc_hd__buf_1
X_23150_ net5012 net4754 VGND VGND VPWR VPWR _03020_ sky130_fd_sc_hd__nand2_2
XFILLER_0_130_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20362_ net6374 net1558 VGND VGND VPWR VPWR _12163_ sky130_fd_sc_hd__nor2_1
X_22101_ net9018 _12500_ _12503_ _02107_ VGND VGND VPWR VPWR _00528_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23081_ net4969 net4712 VGND VGND VPWR VPWR _02951_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20293_ net6516 _12097_ _12098_ net6494 VGND VGND VPWR VPWR _12099_ sky130_fd_sc_hd__o22ai_1
X_22032_ net5799 net5375 VGND VGND VPWR VPWR _02039_ sky130_fd_sc_hd__nand2_2
XFILLER_0_11_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23983_ _03753_ _03779_ net511 VGND VGND VPWR VPWR _03847_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25722_ clknet_4_5__leaf_clk _00595_ net8609 VGND VGND VPWR VPWR pid_d.mult0.a\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_22934_ net4331 _02822_ _02823_ net271 net4362 VGND VGND VPWR VPWR _02824_ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22865_ net5364 _02760_ _02761_ VGND VGND VPWR VPWR _02762_ sky130_fd_sc_hd__a21oi_2
X_25653_ clknet_leaf_2_clk _00526_ net8570 VGND VGND VPWR VPWR pid_d.curr_int\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24604_ _04455_ _04458_ VGND VGND VPWR VPWR _04459_ sky130_fd_sc_hd__xnor2_1
X_21816_ _01804_ _01806_ _01824_ _01725_ VGND VGND VPWR VPWR _01825_ sky130_fd_sc_hd__a22o_1
X_25584_ clknet_leaf_86_clk _00457_ net8532 VGND VGND VPWR VPWR cordic0.cos\[4\] sky130_fd_sc_hd__dfrtp_1
X_22796_ pid_d.kp\[10\] net3069 net2035 VGND VGND VPWR VPWR _02706_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24535_ net5170 pid_q.prev_int\[14\] VGND VGND VPWR VPWR _04391_ sky130_fd_sc_hd__xnor2_1
X_21747_ net5703 net5538 VGND VGND VPWR VPWR _01757_ sky130_fd_sc_hd__nand2_1
Xwire8302 net8303 VGND VGND VPWR VPWR net8302 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8313 net8314 VGND VGND VPWR VPWR net8313 sky130_fd_sc_hd__clkbuf_1
Xmax_length4011 _09358_ VGND VGND VPWR VPWR net4011 sky130_fd_sc_hd__buf_1
Xwire8324 net8325 VGND VGND VPWR VPWR net8324 sky130_fd_sc_hd__clkbuf_1
X_24466_ pid_q.prev_error\[11\] pid_q.curr_error\[11\] _04253_ VGND VGND VPWR VPWR
+ _04324_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_19_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8346 net8343 VGND VGND VPWR VPWR net8346 sky130_fd_sc_hd__buf_1
XFILLER_0_0_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire7612 net7613 VGND VGND VPWR VPWR net7612 sky130_fd_sc_hd__clkbuf_1
X_21678_ _01586_ _01587_ _01688_ VGND VGND VPWR VPWR _01689_ sky130_fd_sc_hd__a21bo_1
Xwire7623 net7624 VGND VGND VPWR VPWR net7623 sky130_fd_sc_hd__clkbuf_1
Xwire8368 net8362 VGND VGND VPWR VPWR net8368 sky130_fd_sc_hd__buf_1
XFILLER_0_81_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23417_ _03283_ _03286_ VGND VGND VPWR VPWR _03287_ sky130_fd_sc_hd__xnor2_2
Xwire7645 net7641 VGND VGND VPWR VPWR net7645 sky130_fd_sc_hd__buf_1
X_20629_ net1395 _12397_ _08992_ VGND VGND VPWR VPWR _12409_ sky130_fd_sc_hd__o21a_1
Xmax_length3343 _08946_ VGND VGND VPWR VPWR net3343 sky130_fd_sc_hd__buf_1
Xwire7656 net7649 VGND VGND VPWR VPWR net7656 sky130_fd_sc_hd__clkbuf_1
X_24397_ _04253_ _04254_ VGND VGND VPWR VPWR _04256_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6911 net6912 VGND VGND VPWR VPWR net6911 sky130_fd_sc_hd__buf_1
Xwire7667 net7668 VGND VGND VPWR VPWR net7667 sky130_fd_sc_hd__clkbuf_1
Xmax_length3354 net3355 VGND VGND VPWR VPWR net3354 sky130_fd_sc_hd__buf_1
Xwire6922 net6919 VGND VGND VPWR VPWR net6922 sky130_fd_sc_hd__clkbuf_1
Xwire7678 svm0.periodTop\[12\] VGND VGND VPWR VPWR net7678 sky130_fd_sc_hd__clkbuf_1
Xmax_length3365 net3366 VGND VGND VPWR VPWR net3365 sky130_fd_sc_hd__clkbuf_2
Xmax_length2620 _08636_ VGND VGND VPWR VPWR net2620 sky130_fd_sc_hd__buf_1
X_14150_ _06409_ net833 VGND VGND VPWR VPWR _06411_ sky130_fd_sc_hd__xor2_2
Xwire7689 net7690 VGND VGND VPWR VPWR net7689 sky130_fd_sc_hd__clkbuf_1
Xwire6944 net6939 VGND VGND VPWR VPWR net6944 sky130_fd_sc_hd__buf_1
X_23348_ net4957 net4673 VGND VGND VPWR VPWR _03218_ sky130_fd_sc_hd__nand2_1
Xmax_length3387 net3388 VGND VGND VPWR VPWR net3387 sky130_fd_sc_hd__buf_1
Xwire6955 net6956 VGND VGND VPWR VPWR net6955 sky130_fd_sc_hd__clkbuf_2
Xwire6966 net6968 VGND VGND VPWR VPWR net6966 sky130_fd_sc_hd__buf_1
X_13101_ net7725 net2355 _05035_ VGND VGND VPWR VPWR _05374_ sky130_fd_sc_hd__and3_1
Xwire6977 net6973 VGND VGND VPWR VPWR net6977 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14081_ _06342_ _06343_ VGND VGND VPWR VPWR _06344_ sky130_fd_sc_hd__xnor2_1
Xwire6999 net6998 VGND VGND VPWR VPWR net6999 sky130_fd_sc_hd__clkbuf_1
X_23279_ net1676 _03148_ VGND VGND VPWR VPWR _03149_ sky130_fd_sc_hd__xnor2_2
X_25018_ net4462 net1631 net2394 _04772_ VGND VGND VPWR VPWR _00780_ sky130_fd_sc_hd__a22o_1
X_13032_ _05279_ _05304_ VGND VGND VPWR VPWR _05305_ sky130_fd_sc_hd__xnor2_1
Xmax_length1985 net1986 VGND VGND VPWR VPWR net1985 sky130_fd_sc_hd__clkbuf_1
X_17840_ _09648_ net3261 VGND VGND VPWR VPWR _09691_ sky130_fd_sc_hd__xnor2_1
X_17771_ net7092 net7116 VGND VGND VPWR VPWR _09622_ sky130_fd_sc_hd__or2b_1
X_14983_ _06981_ _06986_ VGND VGND VPWR VPWR _07057_ sky130_fd_sc_hd__xnor2_1
Xwire1240 net1241 VGND VGND VPWR VPWR net1240 sky130_fd_sc_hd__buf_1
X_19510_ net3866 _11290_ VGND VGND VPWR VPWR _11347_ sky130_fd_sc_hd__or2_1
Xwire1251 _08252_ VGND VGND VPWR VPWR net1251 sky130_fd_sc_hd__buf_1
XFILLER_0_92_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16722_ matmul0.matmul_stage_inst.mult2\[14\] matmul0.matmul_stage_inst.mult1\[14\]
+ VGND VGND VPWR VPWR _08748_ sky130_fd_sc_hd__nand2_1
X_13934_ _06098_ _06103_ _06096_ VGND VGND VPWR VPWR _06200_ sky130_fd_sc_hd__a21o_1
Xwire1262 _07993_ VGND VGND VPWR VPWR net1262 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_156_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1273 _07498_ VGND VGND VPWR VPWR net1273 sky130_fd_sc_hd__buf_1
Xwire1284 _07122_ VGND VGND VPWR VPWR net1284 sky130_fd_sc_hd__clkbuf_1
Xwire1295 _06608_ VGND VGND VPWR VPWR net1295 sky130_fd_sc_hd__buf_1
X_19441_ net3161 _11275_ _11276_ _11277_ VGND VGND VPWR VPWR _11278_ sky130_fd_sc_hd__a211o_1
XFILLER_0_44_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16653_ matmul0.matmul_stage_inst.mult2\[5\] matmul0.matmul_stage_inst.mult1\[5\]
+ VGND VGND VPWR VPWR _08689_ sky130_fd_sc_hd__xor2_1
X_13865_ _06129_ _06130_ _06131_ VGND VGND VPWR VPWR _06132_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15604_ _07594_ _07595_ _07675_ VGND VGND VPWR VPWR _07676_ sky130_fd_sc_hd__o21a_1
X_12816_ net7804 net1610 VGND VGND VPWR VPWR _05089_ sky130_fd_sc_hd__nand2_1
X_19372_ net6152 _11207_ VGND VGND VPWR VPWR _11209_ sky130_fd_sc_hd__nor2_1
X_16584_ _08639_ VGND VGND VPWR VPWR _00233_ sky130_fd_sc_hd__clkbuf_1
X_13796_ _06050_ _06063_ VGND VGND VPWR VPWR _06064_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_84_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18323_ net6892 net6872 VGND VGND VPWR VPWR _10174_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8730 net8733 VGND VGND VPWR VPWR net8730 sky130_fd_sc_hd__buf_2
X_15535_ _07604_ net2227 VGND VGND VPWR VPWR _07608_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12747_ _05004_ net851 VGND VGND VPWR VPWR _05020_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8763 net8798 VGND VGND VPWR VPWR net8763 sky130_fd_sc_hd__buf_1
XFILLER_0_155_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18254_ _10102_ _10104_ VGND VGND VPWR VPWR _10105_ sky130_fd_sc_hd__xor2_1
XFILLER_0_127_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12678_ net7881 net1981 net2359 VGND VGND VPWR VPWR _04951_ sky130_fd_sc_hd__and3_1
X_15466_ _07525_ _07539_ VGND VGND VPWR VPWR _07540_ sky130_fd_sc_hd__xor2_1
XFILLER_0_155_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17205_ net1922 _09153_ VGND VGND VPWR VPWR _09155_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14417_ matmul0.beta_pass\[6\] net1294 net2890 net4443 _06616_ VGND VGND VPWR VPWR
+ _06617_ sky130_fd_sc_hd__a221o_1
Xwire8880 net8873 VGND VGND VPWR VPWR net8880 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18185_ _10030_ _09630_ _10033_ net3254 _10035_ VGND VGND VPWR VPWR _10036_ sky130_fd_sc_hd__o221a_1
X_15397_ _07342_ _07411_ _07469_ _07470_ VGND VGND VPWR VPWR _07471_ sky130_fd_sc_hd__a22oi_2
Xwire8891 net8892 VGND VGND VPWR VPWR net8891 sky130_fd_sc_hd__buf_1
XFILLER_0_142_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17136_ net6914 net1819 _09089_ VGND VGND VPWR VPWR _09091_ sky130_fd_sc_hd__or3_1
Xwire570 _11485_ VGND VGND VPWR VPWR net570 sky130_fd_sc_hd__clkbuf_1
X_14348_ net8217 net3646 VGND VGND VPWR VPWR _06563_ sky130_fd_sc_hd__and2_1
Xwire581 net582 VGND VGND VPWR VPWR net581 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire592 net593 VGND VGND VPWR VPWR net592 sky130_fd_sc_hd__buf_1
X_14279_ net55 net2914 _06517_ net7954 VGND VGND VPWR VPWR _00050_ sky130_fd_sc_hd__a22o_1
X_17067_ net7004 VGND VGND VPWR VPWR _09026_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16018_ _08083_ _08085_ VGND VGND VPWR VPWR _08086_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17969_ _09818_ _09819_ net6909 net6946 net6845 VGND VGND VPWR VPWR _09820_ sky130_fd_sc_hd__o2111a_1
X_19708_ _11543_ VGND VGND VPWR VPWR _11544_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20980_ _00993_ _00976_ VGND VGND VPWR VPWR _00996_ sky130_fd_sc_hd__or2b_1
XFILLER_0_192_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19639_ _11413_ _11415_ VGND VGND VPWR VPWR _11476_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22650_ _02553_ _02574_ _02575_ net3081 VGND VGND VPWR VPWR _02610_ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21601_ net5416 net5893 _01513_ VGND VGND VPWR VPWR _01613_ sky130_fd_sc_hd__and3_1
XFILLER_0_164_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22581_ net4367 net3767 VGND VGND VPWR VPWR _02561_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24320_ _04178_ _04111_ _04179_ VGND VGND VPWR VPWR _04180_ sky130_fd_sc_hd__a21o_1
X_21532_ _01542_ _01543_ VGND VGND VPWR VPWR _01544_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24251_ pid_q.prev_error\[9\] pid_q.curr_error\[9\] VGND VGND VPWR VPWR _04112_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21463_ _01470_ _01475_ VGND VGND VPWR VPWR _01476_ sky130_fd_sc_hd__xnor2_1
Xwire6207 net6208 VGND VGND VPWR VPWR net6207 sky130_fd_sc_hd__clkbuf_1
Xwire6218 net6219 VGND VGND VPWR VPWR net6218 sky130_fd_sc_hd__buf_1
Xwire6229 net6230 VGND VGND VPWR VPWR net6229 sky130_fd_sc_hd__clkbuf_2
X_23202_ _03067_ _03048_ _03070_ _03071_ VGND VGND VPWR VPWR _03072_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_105_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20414_ _12205_ _12210_ VGND VGND VPWR VPWR _12211_ sky130_fd_sc_hd__xnor2_1
X_24182_ _04022_ net590 VGND VGND VPWR VPWR _04043_ sky130_fd_sc_hd__nand2_1
Xwire5506 net5507 VGND VGND VPWR VPWR net5506 sky130_fd_sc_hd__clkbuf_1
Xwire5517 net5518 VGND VGND VPWR VPWR net5517 sky130_fd_sc_hd__clkbuf_1
Xmax_length1204 _10343_ VGND VGND VPWR VPWR net1204 sky130_fd_sc_hd__clkbuf_1
X_21394_ _01403_ _01407_ VGND VGND VPWR VPWR _01408_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5528 net5523 VGND VGND VPWR VPWR net5528 sky130_fd_sc_hd__buf_1
Xwire5539 net5540 VGND VGND VPWR VPWR net5539 sky130_fd_sc_hd__buf_1
X_23133_ _02913_ _02915_ VGND VGND VPWR VPWR _03003_ sky130_fd_sc_hd__xor2_1
Xwire4805 net4798 VGND VGND VPWR VPWR net4805 sky130_fd_sc_hd__buf_1
Xwire4816 net4817 VGND VGND VPWR VPWR net4816 sky130_fd_sc_hd__buf_1
X_20345_ net6516 net6466 _08836_ _12146_ VGND VGND VPWR VPWR _12147_ sky130_fd_sc_hd__or4_1
Xwire4827 net4828 VGND VGND VPWR VPWR net4827 sky130_fd_sc_hd__buf_1
XFILLER_0_141_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4838 net4839 VGND VGND VPWR VPWR net4838 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23064_ net5147 net4561 VGND VGND VPWR VPWR _02934_ sky130_fd_sc_hd__nand2_1
X_20276_ _12083_ VGND VGND VPWR VPWR _00482_ sky130_fd_sc_hd__clkbuf_1
X_22015_ net471 _02003_ _02004_ VGND VGND VPWR VPWR _02022_ sky130_fd_sc_hd__a21oi_1
X_23966_ net4663 net4688 _03373_ VGND VGND VPWR VPWR _03830_ sky130_fd_sc_hd__and3_1
XFILLER_0_187_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length8855 net8856 VGND VGND VPWR VPWR net8855 sky130_fd_sc_hd__clkbuf_1
X_25705_ clknet_leaf_3_clk _00578_ net8580 VGND VGND VPWR VPWR pid_d.mult0.b\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_169_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22917_ _02808_ VGND VGND VPWR VPWR _00643_ sky130_fd_sc_hd__clkbuf_1
X_23897_ pid_q.curr_error\[4\] VGND VGND VPWR VPWR _03762_ sky130_fd_sc_hd__inv_2
Xmax_length8888 net8889 VGND VGND VPWR VPWR net8888 sky130_fd_sc_hd__buf_1
X_13650_ _05798_ _05804_ VGND VGND VPWR VPWR _05920_ sky130_fd_sc_hd__nand2_1
X_25636_ clknet_leaf_104_clk _00509_ net8359 VGND VGND VPWR VPWR cordic0.vec\[0\]\[8\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_39_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22848_ _02744_ _02737_ _02746_ VGND VGND VPWR VPWR _02747_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12601_ _04879_ VGND VGND VPWR VPWR _00007_ sky130_fd_sc_hd__clkbuf_1
X_13581_ _05850_ _05851_ VGND VGND VPWR VPWR _05852_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22779_ _02697_ VGND VGND VPWR VPWR _00616_ sky130_fd_sc_hd__clkbuf_1
X_25567_ clknet_leaf_98_clk _00440_ net8381 VGND VGND VPWR VPWR cordic0.sin\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8110 net8111 VGND VGND VPWR VPWR net8110 sky130_fd_sc_hd__clkbuf_1
X_15320_ _06996_ _07001_ _07393_ VGND VGND VPWR VPWR _07394_ sky130_fd_sc_hd__o21a_1
X_24518_ _04268_ net792 VGND VGND VPWR VPWR _04375_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8132 net8133 VGND VGND VPWR VPWR net8132 sky130_fd_sc_hd__clkbuf_1
X_25498_ clknet_leaf_42_clk _00378_ net8782 VGND VGND VPWR VPWR svm0.delta\[3\] sky130_fd_sc_hd__dfrtp_2
Xwire8143 net8144 VGND VGND VPWR VPWR net8143 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6613 net6625 VGND VGND VPWR VPWR net6613 sky130_fd_sc_hd__buf_1
Xwire8154 net8155 VGND VGND VPWR VPWR net8154 sky130_fd_sc_hd__clkbuf_1
Xwire8165 net8166 VGND VGND VPWR VPWR net8165 sky130_fd_sc_hd__clkbuf_1
Xwire7420 matmul0.matmul_stage_inst.b\[10\] VGND VGND VPWR VPWR net7420 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8176 net8177 VGND VGND VPWR VPWR net8176 sky130_fd_sc_hd__clkbuf_1
X_15251_ net1878 _07313_ net1275 VGND VGND VPWR VPWR _07325_ sky130_fd_sc_hd__o21a_1
XFILLER_0_81_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24449_ _04284_ _04306_ VGND VGND VPWR VPWR _04307_ sky130_fd_sc_hd__xor2_2
Xwire7442 net7440 VGND VGND VPWR VPWR net7442 sky130_fd_sc_hd__buf_1
Xwire8187 net8188 VGND VGND VPWR VPWR net8187 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout5912 net5918 VGND VGND VPWR VPWR net5912 sky130_fd_sc_hd__buf_1
Xwire8198 net8199 VGND VGND VPWR VPWR net8198 sky130_fd_sc_hd__clkbuf_1
Xwire6730 net6731 VGND VGND VPWR VPWR net6730 sky130_fd_sc_hd__clkbuf_1
X_14202_ _06438_ _06461_ VGND VGND VPWR VPWR _06462_ sky130_fd_sc_hd__xnor2_1
Xwire7475 net7476 VGND VGND VPWR VPWR net7475 sky130_fd_sc_hd__clkbuf_1
X_15182_ net1886 _07234_ VGND VGND VPWR VPWR _07256_ sky130_fd_sc_hd__nand2_1
Xwire6741 svm0.counter\[0\] VGND VGND VPWR VPWR net6741 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire7486 net7483 VGND VGND VPWR VPWR net7486 sky130_fd_sc_hd__buf_1
Xwire6752 net6753 VGND VGND VPWR VPWR net6752 sky130_fd_sc_hd__clkbuf_1
X_14133_ _06371_ _06393_ VGND VGND VPWR VPWR _06395_ sky130_fd_sc_hd__nand2_2
Xmax_length2461 _02523_ VGND VGND VPWR VPWR net2461 sky130_fd_sc_hd__buf_1
Xwire6774 net6775 VGND VGND VPWR VPWR net6774 sky130_fd_sc_hd__clkbuf_2
X_19990_ _11772_ _11777_ _11820_ VGND VGND VPWR VPWR _11821_ sky130_fd_sc_hd__a21o_1
Xwire6785 net6782 VGND VGND VPWR VPWR net6785 sky130_fd_sc_hd__buf_1
Xwire6796 net6795 VGND VGND VPWR VPWR net6796 sky130_fd_sc_hd__clkbuf_4
X_14064_ net7680 net1122 _06301_ net1315 net7706 VGND VGND VPWR VPWR _06327_ sky130_fd_sc_hd__a32o_1
X_18941_ _10764_ _10765_ _10778_ _10779_ VGND VGND VPWR VPWR _10780_ sky130_fd_sc_hd__a31oi_1
X_13015_ net7878 _05287_ VGND VGND VPWR VPWR _05288_ sky130_fd_sc_hd__xnor2_1
X_18872_ net6881 net6814 VGND VGND VPWR VPWR _10714_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17823_ net6989 net6965 VGND VGND VPWR VPWR _09674_ sky130_fd_sc_hd__nor2b_1
Xhold3 matmul0.matmul_stage_inst.a\[10\] VGND VGND VPWR VPWR net8956 sky130_fd_sc_hd__dlygate4sd3_1
X_17754_ net7105 net3998 VGND VGND VPWR VPWR _09605_ sky130_fd_sc_hd__nand2_1
X_14966_ net3567 net3562 net3560 net3558 VGND VGND VPWR VPWR _07040_ sky130_fd_sc_hd__o2bb2a_1
Xwire1070 _10420_ VGND VGND VPWR VPWR net1070 sky130_fd_sc_hd__buf_1
X_16705_ _08733_ VGND VGND VPWR VPWR _00260_ sky130_fd_sc_hd__clkbuf_1
Xwire1081 net1082 VGND VGND VPWR VPWR net1081 sky130_fd_sc_hd__dlymetal6s2s_1
X_13917_ net1311 net1583 _06181_ net7633 _06182_ VGND VGND VPWR VPWR _06183_ sky130_fd_sc_hd__o221a_1
XFILLER_0_18_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1092 _08129_ VGND VGND VPWR VPWR net1092 sky130_fd_sc_hd__dlymetal6s2s_1
X_17685_ net4015 svm0.tA\[10\] net6746 _09526_ _09564_ VGND VGND VPWR VPWR _09565_
+ sky130_fd_sc_hd__a221o_1
X_14897_ net6612 net7421 matmul0.matmul_stage_inst.a\[9\] net6580 VGND VGND VPWR VPWR
+ _06971_ sky130_fd_sc_hd__a22o_1
XFILLER_0_159_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19424_ net6299 _11258_ _11260_ VGND VGND VPWR VPWR _11261_ sky130_fd_sc_hd__a21o_1
XFILLER_0_162_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16636_ _08671_ _08665_ _08666_ _08673_ VGND VGND VPWR VPWR _08674_ sky130_fd_sc_hd__a31o_1
X_13848_ net7641 net1311 VGND VGND VPWR VPWR _06115_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19355_ _11120_ _11190_ _11191_ net3213 VGND VGND VPWR VPWR _11192_ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16567_ _08550_ _08625_ VGND VGND VPWR VPWR _08626_ sky130_fd_sc_hd__nor2_1
X_13779_ _05943_ _05944_ _05950_ _05951_ VGND VGND VPWR VPWR _06047_ sky130_fd_sc_hd__and4_1
XFILLER_0_73_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18306_ net1775 _10156_ VGND VGND VPWR VPWR _10157_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15518_ _07525_ _07539_ net1113 VGND VGND VPWR VPWR _07591_ sky130_fd_sc_hd__a21o_1
XFILLER_0_183_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19286_ net6258 _11119_ _11121_ net3173 VGND VGND VPWR VPWR _11123_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16498_ _08556_ _08557_ VGND VGND VPWR VPWR _08558_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18237_ net7142 net2554 net7095 VGND VGND VPWR VPWR _10088_ sky130_fd_sc_hd__a21oi_1
X_15449_ _07510_ _07522_ VGND VGND VPWR VPWR _07523_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_111_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18168_ net1212 _10006_ _10018_ _10012_ VGND VGND VPWR VPWR _10019_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_20_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17119_ _09072_ _09074_ VGND VGND VPWR VPWR _09075_ sky130_fd_sc_hd__xnor2_2
X_18099_ _09943_ _09947_ net962 VGND VGND VPWR VPWR _09950_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20130_ _11927_ _11932_ _11957_ VGND VGND VPWR VPWR _11958_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20061_ net6095 net6021 VGND VGND VPWR VPWR _11890_ sky130_fd_sc_hd__xor2_2
XFILLER_0_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23820_ _03681_ _03684_ VGND VGND VPWR VPWR _03685_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_174_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23751_ net4674 net4859 VGND VGND VPWR VPWR _03617_ sky130_fd_sc_hd__nand2_1
X_20963_ net3823 net3808 VGND VGND VPWR VPWR _00979_ sky130_fd_sc_hd__nor2_1
Xmax_length7428 matmul0.matmul_stage_inst.b\[5\] VGND VGND VPWR VPWR net7428 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_92_clk clknet_4_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_92_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22702_ pid_d.ki\[11\] net2446 net3696 pid_d.kp\[11\] VGND VGND VPWR VPWR _02643_
+ sky130_fd_sc_hd__a22o_1
X_23682_ _03433_ _03434_ _03435_ VGND VGND VPWR VPWR _03549_ sky130_fd_sc_hd__o21a_1
XFILLER_0_36_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20894_ _00900_ net2481 _00909_ VGND VGND VPWR VPWR _00910_ sky130_fd_sc_hd__a21o_1
X_25421_ clknet_leaf_99_clk _00304_ net8382 VGND VGND VPWR VPWR matmul0.cos\[8\] sky130_fd_sc_hd__dfrtp_1
X_22633_ net7368 net3090 net3080 _01245_ VGND VGND VPWR VPWR _02601_ sky130_fd_sc_hd__a211o_1
XFILLER_0_165_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25352_ clknet_leaf_84_clk _00235_ net8507 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult2\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_22564_ _02547_ VGND VGND VPWR VPWR _02548_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_134_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24303_ net1013 net1656 net2022 VGND VGND VPWR VPWR _04163_ sky130_fd_sc_hd__o21a_1
X_21515_ net860 _01522_ VGND VGND VPWR VPWR _01528_ sky130_fd_sc_hd__nor2_1
XFILLER_0_133_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25283_ clknet_leaf_77_clk _00166_ net8440 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.c\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_22495_ _02429_ _02436_ _02495_ VGND VGND VPWR VPWR _02496_ sky130_fd_sc_hd__o21a_1
Xwire6004 net6006 VGND VGND VPWR VPWR net6004 sky130_fd_sc_hd__buf_1
XFILLER_0_185_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout5219 matmul0.beta_pass\[10\] VGND VGND VPWR VPWR net5219 sky130_fd_sc_hd__buf_1
Xwire6015 net6014 VGND VGND VPWR VPWR net6015 sky130_fd_sc_hd__clkbuf_1
X_24234_ net1013 _04094_ VGND VGND VPWR VPWR _04095_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_106_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6026 net6024 VGND VGND VPWR VPWR net6026 sky130_fd_sc_hd__buf_1
X_21446_ _01455_ _01458_ VGND VGND VPWR VPWR _01459_ sky130_fd_sc_hd__xnor2_2
Xwire6037 net6038 VGND VGND VPWR VPWR net6037 sky130_fd_sc_hd__buf_1
Xfanout4507 pid_q.mult0.a\[14\] VGND VGND VPWR VPWR net4507 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5303 net5305 VGND VGND VPWR VPWR net5303 sky130_fd_sc_hd__clkbuf_1
Xwire6048 net6049 VGND VGND VPWR VPWR net6048 sky130_fd_sc_hd__buf_1
XFILLER_0_44_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5314 pid_d.out\[15\] VGND VGND VPWR VPWR net5314 sky130_fd_sc_hd__buf_1
Xwire6059 net6060 VGND VGND VPWR VPWR net6059 sky130_fd_sc_hd__clkbuf_1
Xwire5325 net5326 VGND VGND VPWR VPWR net5325 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24165_ _03961_ _04026_ VGND VGND VPWR VPWR _04027_ sky130_fd_sc_hd__xnor2_1
Xwire5336 net5337 VGND VGND VPWR VPWR net5336 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5347 net5348 VGND VGND VPWR VPWR net5347 sky130_fd_sc_hd__clkbuf_1
X_21377_ net1728 _01390_ VGND VGND VPWR VPWR _01391_ sky130_fd_sc_hd__xnor2_1
Xwire4613 net4609 VGND VGND VPWR VPWR net4613 sky130_fd_sc_hd__buf_1
XFILLER_0_160_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5358 net5359 VGND VGND VPWR VPWR net5358 sky130_fd_sc_hd__clkbuf_1
Xwire4624 net4625 VGND VGND VPWR VPWR net4624 sky130_fd_sc_hd__buf_1
Xwire5369 pid_d.out\[0\] VGND VGND VPWR VPWR net5369 sky130_fd_sc_hd__clkbuf_1
X_23116_ _02889_ _02985_ VGND VGND VPWR VPWR _02986_ sky130_fd_sc_hd__xnor2_1
Xwire4635 net4638 VGND VGND VPWR VPWR net4635 sky130_fd_sc_hd__clkbuf_1
Xwire3901 _10822_ VGND VGND VPWR VPWR net3901 sky130_fd_sc_hd__buf_1
X_20328_ _12131_ VGND VGND VPWR VPWR _00486_ sky130_fd_sc_hd__clkbuf_1
X_24096_ pid_q.curr_int\[8\] pid_q.prev_int\[8\] VGND VGND VPWR VPWR _03958_ sky130_fd_sc_hd__xor2_1
Xwire4657 net4658 VGND VGND VPWR VPWR net4657 sky130_fd_sc_hd__clkbuf_1
Xwire3912 net3913 VGND VGND VPWR VPWR net3912 sky130_fd_sc_hd__clkbuf_1
Xwire4668 net4656 VGND VGND VPWR VPWR net4668 sky130_fd_sc_hd__buf_1
Xwire3923 _10335_ VGND VGND VPWR VPWR net3923 sky130_fd_sc_hd__buf_1
Xwire3934 net3935 VGND VGND VPWR VPWR net3934 sky130_fd_sc_hd__buf_1
XFILLER_0_102_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23047_ _02895_ _02916_ VGND VGND VPWR VPWR _02917_ sky130_fd_sc_hd__xnor2_1
Xwire3945 _09879_ VGND VGND VPWR VPWR net3945 sky130_fd_sc_hd__clkbuf_1
X_20259_ _12071_ VGND VGND VPWR VPWR _00477_ sky130_fd_sc_hd__clkbuf_1
Xwire3956 net3961 VGND VGND VPWR VPWR net3956 sky130_fd_sc_hd__buf_1
Xwire3967 net3968 VGND VGND VPWR VPWR net3967 sky130_fd_sc_hd__buf_1
Xwire3978 net3979 VGND VGND VPWR VPWR net3978 sky130_fd_sc_hd__clkbuf_1
Xwire3989 _09660_ VGND VGND VPWR VPWR net3989 sky130_fd_sc_hd__buf_1
X_14820_ net8984 net2872 _06926_ VGND VGND VPWR VPWR _00182_ sky130_fd_sc_hd__a21o_1
X_24998_ net9163 net1632 net2395 _04755_ VGND VGND VPWR VPWR _00777_ sky130_fd_sc_hd__a22o_1
X_14751_ _06839_ _06882_ VGND VGND VPWR VPWR _06883_ sky130_fd_sc_hd__nand2_1
X_23949_ _03694_ _03696_ _03812_ VGND VGND VPWR VPWR _03813_ sky130_fd_sc_hd__a21oi_2
Xmax_length8652 net8649 VGND VGND VPWR VPWR net8652 sky130_fd_sc_hd__buf_1
XFILLER_0_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_83_clk clknet_4_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_83_clk sky130_fd_sc_hd__clkbuf_16
X_13702_ _05967_ _05970_ VGND VGND VPWR VPWR _05971_ sky130_fd_sc_hd__xnor2_1
X_17470_ _09361_ _09362_ VGND VGND VPWR VPWR _09363_ sky130_fd_sc_hd__nor2_1
X_14682_ net9033 net2868 _06825_ net3617 VGND VGND VPWR VPWR _00139_ sky130_fd_sc_hd__a22o_1
XFILLER_0_168_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16421_ _08427_ VGND VGND VPWR VPWR _08483_ sky130_fd_sc_hd__inv_2
Xmax_length7995 pid_q.target\[8\] VGND VGND VPWR VPWR net7995 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13633_ _05825_ _05826_ net7671 net1150 VGND VGND VPWR VPWR _05903_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_17_Left_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25619_ clknet_leaf_110_clk _00492_ net8347 VGND VGND VPWR VPWR cordic0.slte0.opA\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19140_ net6180 net6158 VGND VGND VPWR VPWR _10977_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16352_ net978 _08337_ _08414_ VGND VGND VPWR VPWR _08415_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_82_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13564_ _05806_ _05834_ VGND VGND VPWR VPWR _05835_ sky130_fd_sc_hd__xnor2_1
Xfanout7122 net7126 VGND VGND VPWR VPWR net7122 sky130_fd_sc_hd__clkbuf_1
X_15303_ net2852 VGND VGND VPWR VPWR _07377_ sky130_fd_sc_hd__buf_1
X_19071_ _10869_ _10889_ VGND VGND VPWR VPWR _10908_ sky130_fd_sc_hd__or2_1
X_13495_ _05636_ _05650_ VGND VGND VPWR VPWR _05768_ sky130_fd_sc_hd__or2_1
X_16283_ net1253 _08340_ _08346_ VGND VGND VPWR VPWR _08347_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_180_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout6443 net6444 VGND VGND VPWR VPWR net6443 sky130_fd_sc_hd__buf_2
Xwire7250 net7251 VGND VGND VPWR VPWR net7250 sky130_fd_sc_hd__clkbuf_2
X_18022_ net7107 _09624_ VGND VGND VPWR VPWR _09873_ sky130_fd_sc_hd__xnor2_2
Xwire7261 net7262 VGND VGND VPWR VPWR net7261 sky130_fd_sc_hd__clkbuf_1
X_15234_ _07302_ net3443 _07307_ VGND VGND VPWR VPWR _07308_ sky130_fd_sc_hd__o21a_1
Xwire7272 net7273 VGND VGND VPWR VPWR net7272 sky130_fd_sc_hd__clkbuf_1
Xwire7283 net7284 VGND VGND VPWR VPWR net7283 sky130_fd_sc_hd__buf_1
XFILLER_0_34_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout6498 net6504 VGND VGND VPWR VPWR net6498 sky130_fd_sc_hd__buf_2
Xwire7294 net7295 VGND VGND VPWR VPWR net7294 sky130_fd_sc_hd__buf_1
XFILLER_0_23_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6560 net6561 VGND VGND VPWR VPWR net6560 sky130_fd_sc_hd__clkbuf_1
X_15165_ net1893 _07238_ VGND VGND VPWR VPWR _07239_ sky130_fd_sc_hd__xnor2_2
Xwire6582 net6583 VGND VGND VPWR VPWR net6582 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire6593 net6595 VGND VGND VPWR VPWR net6593 sky130_fd_sc_hd__clkbuf_1
X_14116_ net7647 net1123 VGND VGND VPWR VPWR _06378_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5870 net5871 VGND VGND VPWR VPWR net5870 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_26_Left_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19973_ net6052 net6021 VGND VGND VPWR VPWR _11804_ sky130_fd_sc_hd__nor2_1
X_15096_ _07085_ _07090_ VGND VGND VPWR VPWR _07170_ sky130_fd_sc_hd__xnor2_1
Xwire5881 net5878 VGND VGND VPWR VPWR net5881 sky130_fd_sc_hd__buf_1
Xwire5892 net5893 VGND VGND VPWR VPWR net5892 sky130_fd_sc_hd__buf_1
XFILLER_0_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18924_ net1427 _10762_ _10763_ VGND VGND VPWR VPWR _10764_ sky130_fd_sc_hd__o21ba_1
X_14047_ _06290_ _06310_ VGND VGND VPWR VPWR _06311_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18855_ _10696_ _10697_ net1443 VGND VGND VPWR VPWR _10698_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17806_ net7060 net7090 _09620_ VGND VGND VPWR VPWR _09657_ sky130_fd_sc_hd__or3_1
X_18786_ net6862 _10579_ net3967 VGND VGND VPWR VPWR _10630_ sky130_fd_sc_hd__mux2_1
X_15998_ net826 _08065_ _07984_ VGND VGND VPWR VPWR _08066_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_167_Right_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17737_ net6445 net2881 net6447 VGND VGND VPWR VPWR _09592_ sky130_fd_sc_hd__o21a_1
X_14949_ net6543 net6588 net7391 VGND VGND VPWR VPWR _07023_ sky130_fd_sc_hd__o21a_1
XFILLER_0_82_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_74_clk clknet_4_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_74_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_159_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17668_ net6735 svm0.tA\[2\] VGND VGND VPWR VPWR _09548_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_35_Left_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19407_ _11107_ VGND VGND VPWR VPWR _11244_ sky130_fd_sc_hd__inv_2
X_16619_ net7373 net4063 net6558 VGND VGND VPWR VPWR _08660_ sky130_fd_sc_hd__mux2_1
X_17599_ net4006 svm0.tB\[7\] svm0.tB\[5\] net4023 _09479_ VGND VGND VPWR VPWR _09480_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_134_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19338_ net6287 net6334 net6270 VGND VGND VPWR VPWR _11175_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_17_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19269_ _11097_ _11105_ VGND VGND VPWR VPWR _11106_ sky130_fd_sc_hd__nand2_1
X_21300_ _01256_ _01314_ VGND VGND VPWR VPWR _01315_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22280_ net5752 net5378 VGND VGND VPWR VPWR _02284_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold200 cordic0.slte0.opA\[16\] VGND VGND VPWR VPWR net9153 sky130_fd_sc_hd__dlygate4sd3_1
X_21231_ net5987 net3122 net2077 _01246_ VGND VGND VPWR VPWR _00519_ sky130_fd_sc_hd__a22o_1
Xhold211 pid_q.curr_error\[15\] VGND VGND VPWR VPWR net9164 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_44_Left_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold222 pid_q.prev_error\[3\] VGND VGND VPWR VPWR net9175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 svm0.tA\[4\] VGND VGND VPWR VPWR net9186 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 _00799_ VGND VGND VPWR VPWR net9197 sky130_fd_sc_hd__dlygate4sd3_1
X_21162_ _01174_ _12556_ VGND VGND VPWR VPWR _01178_ sky130_fd_sc_hd__nand2_1
Xhold255 cordic0.slte0.opA\[0\] VGND VGND VPWR VPWR net9208 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3208 _10836_ VGND VGND VPWR VPWR net3208 sky130_fd_sc_hd__buf_1
Xhold266 svm0.tB\[7\] VGND VGND VPWR VPWR net9219 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3219 net3220 VGND VGND VPWR VPWR net3219 sky130_fd_sc_hd__clkbuf_1
Xhold277 matmul0.b\[12\] VGND VGND VPWR VPWR net9230 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20113_ net6112 _11937_ _11940_ VGND VGND VPWR VPWR _11941_ sky130_fd_sc_hd__a21oi_2
Xhold288 cordic0.cos\[5\] VGND VGND VPWR VPWR net9241 sky130_fd_sc_hd__dlygate4sd3_1
X_21093_ _01068_ _01108_ VGND VGND VPWR VPWR _01109_ sky130_fd_sc_hd__xnor2_1
Xwire2507 _11270_ VGND VGND VPWR VPWR net2507 sky130_fd_sc_hd__buf_1
XFILLER_0_102_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2518 _11127_ VGND VGND VPWR VPWR net2518 sky130_fd_sc_hd__buf_1
Xwire2529 _10816_ VGND VGND VPWR VPWR net2529 sky130_fd_sc_hd__clkbuf_1
X_24921_ net8866 net139 VGND VGND VPWR VPWR _04708_ sky130_fd_sc_hd__and2b_1
Xwire1806 _08957_ VGND VGND VPWR VPWR net1806 sky130_fd_sc_hd__buf_1
X_20044_ _11846_ _11873_ VGND VGND VPWR VPWR _11874_ sky130_fd_sc_hd__xnor2_1
Xwire1817 _08911_ VGND VGND VPWR VPWR net1817 sky130_fd_sc_hd__buf_1
Xwire1828 _08838_ VGND VGND VPWR VPWR net1828 sky130_fd_sc_hd__buf_1
Xwire1839 _08684_ VGND VGND VPWR VPWR net1839 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24852_ net7502 _04504_ _04540_ net2007 net4787 VGND VGND VPWR VPWR _04659_ sky130_fd_sc_hd__a32o_1
XFILLER_0_99_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23803_ net7527 _03582_ net463 net7468 net1381 VGND VGND VPWR VPWR _03669_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_134_Right_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_53_Left_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24783_ _04608_ _04609_ VGND VGND VPWR VPWR _04610_ sky130_fd_sc_hd__xnor2_1
X_21995_ _01998_ _01999_ _02002_ VGND VGND VPWR VPWR _02003_ sky130_fd_sc_hd__nand3_1
Xclkbuf_leaf_65_clk clknet_4_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_16
X_23734_ net5077 net4508 VGND VGND VPWR VPWR _03600_ sky130_fd_sc_hd__nand2_1
Xmax_length7247 net7248 VGND VGND VPWR VPWR net7247 sky130_fd_sc_hd__clkbuf_1
X_20946_ _00956_ net1734 net3111 VGND VGND VPWR VPWR _00962_ sky130_fd_sc_hd__o21ba_1
Xmax_length6513 net6514 VGND VGND VPWR VPWR net6513 sky130_fd_sc_hd__buf_1
XFILLER_0_95_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23665_ _03411_ _03412_ _03531_ VGND VGND VPWR VPWR _03532_ sky130_fd_sc_hd__a21oi_2
X_20877_ _00889_ _00892_ VGND VGND VPWR VPWR _00893_ sky130_fd_sc_hd__and2_1
X_25404_ clknet_leaf_72_clk _00287_ net8468 VGND VGND VPWR VPWR matmul0.a\[7\] sky130_fd_sc_hd__dfrtp_1
X_22616_ pid_d.curr_error\[12\] net939 net3088 VGND VGND VPWR VPWR _02588_ sky130_fd_sc_hd__mux2_1
X_23596_ _03370_ net1024 VGND VGND VPWR VPWR _03464_ sky130_fd_sc_hd__nor2_1
XFILLER_0_165_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22547_ net5966 net3017 net2461 VGND VGND VPWR VPWR _02536_ sky130_fd_sc_hd__and3_1
X_25335_ clknet_leaf_83_clk _00218_ net8502 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult1\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_11_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13280_ net732 _05552_ VGND VGND VPWR VPWR _05553_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22478_ _02228_ _02433_ _02478_ net5765 VGND VGND VPWR VPWR _02479_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25266_ clknet_leaf_88_clk _00149_ net8430 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.b\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5100 net5101 VGND VGND VPWR VPWR net5100 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5122 net5123 VGND VGND VPWR VPWR net5122 sky130_fd_sc_hd__buf_1
X_24217_ net4993 net4959 VGND VGND VPWR VPWR _04078_ sky130_fd_sc_hd__xor2_1
X_21429_ _01396_ _01409_ _01441_ VGND VGND VPWR VPWR _01442_ sky130_fd_sc_hd__a21o_1
Xwire5133 net5134 VGND VGND VPWR VPWR net5133 sky130_fd_sc_hd__buf_1
X_25197_ clknet_leaf_63_clk _00086_ net8665 VGND VGND VPWR VPWR matmul0.b_in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5155 net5146 VGND VGND VPWR VPWR net5155 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4410 net4411 VGND VGND VPWR VPWR net4410 sky130_fd_sc_hd__clkbuf_1
Xfanout4359 net4371 VGND VGND VPWR VPWR net4359 sky130_fd_sc_hd__buf_1
X_24148_ net4651 _04009_ net4605 net4625 VGND VGND VPWR VPWR _04010_ sky130_fd_sc_hd__or4bb_1
Xwire4421 net4422 VGND VGND VPWR VPWR net4421 sky130_fd_sc_hd__clkbuf_1
Xwire5177 pid_q.curr_int\[11\] VGND VGND VPWR VPWR net5177 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_47_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4432 net4433 VGND VGND VPWR VPWR net4432 sky130_fd_sc_hd__clkbuf_1
Xwire5188 svm0.in_valid VGND VGND VPWR VPWR net5188 sky130_fd_sc_hd__clkbuf_1
Xwire4443 net4444 VGND VGND VPWR VPWR net4443 sky130_fd_sc_hd__clkbuf_1
Xwire4454 net4455 VGND VGND VPWR VPWR net4454 sky130_fd_sc_hd__clkbuf_1
Xwire5199 net5200 VGND VGND VPWR VPWR net5199 sky130_fd_sc_hd__clkbuf_1
Xwire3720 net3721 VGND VGND VPWR VPWR net3720 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4465 pid_q.out\[2\] VGND VGND VPWR VPWR net4465 sky130_fd_sc_hd__clkbuf_1
Xwire4476 net4477 VGND VGND VPWR VPWR net4476 sky130_fd_sc_hd__clkbuf_1
Xwire3731 _04502_ VGND VGND VPWR VPWR net3731 sky130_fd_sc_hd__buf_1
X_24079_ net595 net592 VGND VGND VPWR VPWR _03942_ sky130_fd_sc_hd__nor2_1
X_16970_ _08927_ _08929_ _08931_ net4053 _08825_ net4059 VGND VGND VPWR VPWR _08933_
+ sky130_fd_sc_hd__mux4_1
Xwire3753 net3754 VGND VGND VPWR VPWR net3753 sky130_fd_sc_hd__buf_1
Xwire3764 net3765 VGND VGND VPWR VPWR net3764 sky130_fd_sc_hd__buf_1
X_15921_ net2666 VGND VGND VPWR VPWR _07990_ sky130_fd_sc_hd__clkbuf_1
Xwire3786 net3788 VGND VGND VPWR VPWR net3786 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3797 net3798 VGND VGND VPWR VPWR net3797 sky130_fd_sc_hd__clkbuf_1
X_18640_ net2538 net2539 VGND VGND VPWR VPWR _10487_ sky130_fd_sc_hd__nand2_1
X_15852_ _07831_ _07921_ VGND VGND VPWR VPWR _07922_ sky130_fd_sc_hd__xnor2_1
X_14803_ net9020 net3004 _06918_ VGND VGND VPWR VPWR _00173_ sky130_fd_sc_hd__o21a_1
X_18571_ net6769 net1435 VGND VGND VPWR VPWR _10419_ sky130_fd_sc_hd__nand2_1
X_15783_ _07752_ _07753_ _07754_ VGND VGND VPWR VPWR _07853_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12995_ _05266_ _05267_ VGND VGND VPWR VPWR _05268_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_56_clk clknet_4_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_8_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17522_ _09332_ _09406_ net6657 VGND VGND VPWR VPWR _09407_ sky130_fd_sc_hd__o21ai_1
X_14734_ net7455 _06868_ net2859 VGND VGND VPWR VPWR _06870_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17453_ _09341_ _09342_ net6743 VGND VGND VPWR VPWR _09348_ sky130_fd_sc_hd__a21o_1
XFILLER_0_129_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14665_ _06817_ VGND VGND VPWR VPWR _06818_ sky130_fd_sc_hd__buf_1
XFILLER_0_15_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16404_ _08446_ _08465_ VGND VGND VPWR VPWR _08466_ sky130_fd_sc_hd__xnor2_1
X_13616_ _05882_ _05885_ VGND VGND VPWR VPWR _05886_ sky130_fd_sc_hd__xnor2_1
X_17384_ net2572 _09292_ VGND VGND VPWR VPWR _09293_ sky130_fd_sc_hd__or2_1
XFILLER_0_184_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14596_ net7214 net5200 _06769_ VGND VGND VPWR VPWR _06770_ sky130_fd_sc_hd__or3_1
X_19123_ _10958_ _10959_ VGND VGND VPWR VPWR _10960_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16335_ net1840 _08397_ VGND VGND VPWR VPWR _08398_ sky130_fd_sc_hd__xnor2_1
X_13547_ _05814_ _05815_ _05816_ _05817_ VGND VGND VPWR VPWR _05818_ sky130_fd_sc_hd__nor4_1
XFILLER_0_137_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout6240 net6250 VGND VGND VPWR VPWR net6240 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_82_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19054_ _10884_ _10886_ _10890_ VGND VGND VPWR VPWR _10891_ sky130_fd_sc_hd__a21oi_1
X_16266_ net2651 net2220 _08328_ VGND VGND VPWR VPWR _08330_ sky130_fd_sc_hd__o21ai_1
X_13478_ net7619 net1972 net1969 VGND VGND VPWR VPWR _05751_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18005_ net7004 _09844_ _09853_ _09855_ VGND VGND VPWR VPWR _09856_ sky130_fd_sc_hd__o22a_1
Xwire7091 net7089 VGND VGND VPWR VPWR net7091 sky130_fd_sc_hd__dlymetal6s2s_1
X_15217_ net1881 net1880 net1879 VGND VGND VPWR VPWR _07291_ sky130_fd_sc_hd__o21a_1
Xfanout6295 net6303 VGND VGND VPWR VPWR net6295 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_26_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16197_ _08180_ VGND VGND VPWR VPWR _08262_ sky130_fd_sc_hd__buf_1
XFILLER_0_140_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6390 net6391 VGND VGND VPWR VPWR net6390 sky130_fd_sc_hd__clkbuf_1
X_15148_ _07177_ _07178_ VGND VGND VPWR VPWR _07222_ sky130_fd_sc_hd__xnor2_1
Xfanout4871 net4878 VGND VGND VPWR VPWR net4871 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_168_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19956_ net1409 _11766_ net1410 VGND VGND VPWR VPWR _11787_ sky130_fd_sc_hd__o21a_1
X_15079_ matmul0.matmul_stage_inst.e\[11\] _07151_ _07152_ net7382 VGND VGND VPWR
+ VPWR _07153_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_120_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18907_ _10335_ net275 _10747_ VGND VGND VPWR VPWR _10748_ sky130_fd_sc_hd__or3b_1
X_19887_ net569 _11719_ VGND VGND VPWR VPWR _11720_ sky130_fd_sc_hd__nand2_2
XFILLER_0_93_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_0__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_4_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_18838_ _10679_ _10680_ VGND VGND VPWR VPWR _10681_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18769_ _10607_ _10613_ _10335_ VGND VGND VPWR VPWR _10614_ sky130_fd_sc_hd__mux2_1
XFILLER_0_179_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_47_clk clknet_4_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_179_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20800_ _12547_ _00814_ VGND VGND VPWR VPWR _00816_ sky130_fd_sc_hd__and2_1
XFILLER_0_132_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21780_ _01680_ _01683_ _01789_ VGND VGND VPWR VPWR _01790_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_78_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20731_ _04873_ _00005_ _00002_ _12501_ VGND VGND VPWR VPWR _12502_ sky130_fd_sc_hd__o31a_1
XFILLER_0_65_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8709 net8710 VGND VGND VPWR VPWR net8709 sky130_fd_sc_hd__buf_1
X_23450_ _03262_ _03297_ _03296_ VGND VGND VPWR VPWR _03319_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_46_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20662_ net6109 _12438_ _12439_ VGND VGND VPWR VPWR _00512_ sky130_fd_sc_hd__o21a_1
XFILLER_0_163_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length4418 pid_q.out\[11\] VGND VGND VPWR VPWR net4418 sky130_fd_sc_hd__buf_1
XFILLER_0_58_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22401_ pid_d.prev_error\[14\] pid_d.curr_error\[14\] VGND VGND VPWR VPWR _02403_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_147_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23381_ _03247_ _03250_ VGND VGND VPWR VPWR _03251_ sky130_fd_sc_hd__nor2_1
XFILLER_0_162_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20593_ net1740 _12367_ net1226 VGND VGND VPWR VPWR _12375_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22332_ _02333_ _02334_ VGND VGND VPWR VPWR _02335_ sky130_fd_sc_hd__or2_1
X_25120_ net9217 _04850_ _04853_ net5977 VGND VGND VPWR VPWR _00801_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25051_ _03955_ _04795_ _04800_ VGND VGND VPWR VPWR _04801_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22263_ _02256_ _02265_ _02266_ VGND VGND VPWR VPWR _02267_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24002_ net743 _03864_ VGND VGND VPWR VPWR _03865_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21214_ _01022_ _01226_ _01228_ _01229_ VGND VGND VPWR VPWR _01230_ sky130_fd_sc_hd__o211a_1
XFILLER_0_143_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22194_ net2062 _02192_ _02198_ VGND VGND VPWR VPWR _02199_ sky130_fd_sc_hd__a21bo_1
Xwire3005 net3006 VGND VGND VPWR VPWR net3005 sky130_fd_sc_hd__buf_1
Xwire3016 net3017 VGND VGND VPWR VPWR net3016 sky130_fd_sc_hd__buf_1
X_21145_ _01158_ _01159_ _01160_ VGND VGND VPWR VPWR _01161_ sky130_fd_sc_hd__o21ba_1
Xwire3038 net3039 VGND VGND VPWR VPWR net3038 sky130_fd_sc_hd__clkbuf_1
Xwire3049 _03644_ VGND VGND VPWR VPWR net3049 sky130_fd_sc_hd__buf_1
Xwire2304 _05189_ VGND VGND VPWR VPWR net2304 sky130_fd_sc_hd__buf_1
Xwire2315 net2316 VGND VGND VPWR VPWR net2315 sky130_fd_sc_hd__buf_1
Xwire2326 net2327 VGND VGND VPWR VPWR net2326 sky130_fd_sc_hd__buf_1
Xwire2337 _04931_ VGND VGND VPWR VPWR net2337 sky130_fd_sc_hd__clkbuf_1
X_21076_ _01080_ _01081_ _01091_ VGND VGND VPWR VPWR _01092_ sky130_fd_sc_hd__a21oi_2
Xwire2348 net2349 VGND VGND VPWR VPWR net2348 sky130_fd_sc_hd__buf_1
Xwire1614 _04977_ VGND VGND VPWR VPWR net1614 sky130_fd_sc_hd__clkbuf_1
Xwire2359 net2363 VGND VGND VPWR VPWR net2359 sky130_fd_sc_hd__clkbuf_1
Xwire1625 _04860_ VGND VGND VPWR VPWR net1625 sky130_fd_sc_hd__buf_1
X_24904_ net8871 net130 VGND VGND VPWR VPWR _04694_ sky130_fd_sc_hd__and2b_1
X_20027_ net6168 _11853_ _11856_ VGND VGND VPWR VPWR _11857_ sky130_fd_sc_hd__a21o_1
Xwire1636 net1637 VGND VGND VPWR VPWR net1636 sky130_fd_sc_hd__clkbuf_2
X_25884_ clknet_leaf_17_clk _00757_ net8626 VGND VGND VPWR VPWR pid_q.ki\[12\] sky130_fd_sc_hd__dfrtp_1
Xwire1647 _04507_ VGND VGND VPWR VPWR net1647 sky130_fd_sc_hd__buf_1
Xwire1658 _04011_ VGND VGND VPWR VPWR net1658 sky130_fd_sc_hd__buf_1
Xwire1669 _03366_ VGND VGND VPWR VPWR net1669 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24835_ net4988 _04642_ net2001 net688 VGND VGND VPWR VPWR _00719_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_38_clk clknet_4_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length7022 net7023 VGND VGND VPWR VPWR net7022 sky130_fd_sc_hd__clkbuf_2
Xmax_length7033 net7030 VGND VGND VPWR VPWR net7033 sky130_fd_sc_hd__buf_1
X_24766_ _04593_ _04594_ VGND VGND VPWR VPWR _04595_ sky130_fd_sc_hd__xnor2_1
X_12780_ _05050_ _05051_ _05052_ VGND VGND VPWR VPWR _05053_ sky130_fd_sc_hd__o21ai_1
X_21978_ _01985_ VGND VGND VPWR VPWR _01986_ sky130_fd_sc_hd__inv_2
Xmax_length6321 net6322 VGND VGND VPWR VPWR net6321 sky130_fd_sc_hd__buf_1
X_23717_ net639 _03564_ VGND VGND VPWR VPWR _03583_ sky130_fd_sc_hd__and2b_1
Xmax_length6332 cordic0.vec\[0\]\[2\] VGND VGND VPWR VPWR net6332 sky130_fd_sc_hd__clkbuf_1
X_20929_ net5601 net5832 VGND VGND VPWR VPWR _00945_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24697_ net7501 _04534_ VGND VGND VPWR VPWR _04535_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14450_ _06641_ matmul0.b_in\[14\] net994 VGND VGND VPWR VPWR _06642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23648_ _03513_ _03514_ VGND VGND VPWR VPWR _03515_ sky130_fd_sc_hd__xor2_1
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13401_ _05486_ _05563_ VGND VGND VPWR VPWR _05674_ sky130_fd_sc_hd__nor2_1
Xmax_length4952 net4953 VGND VGND VPWR VPWR net4952 sky130_fd_sc_hd__buf_1
X_14381_ net7210 net1296 net2893 net5320 _06588_ VGND VGND VPWR VPWR _06589_ sky130_fd_sc_hd__a221o_1
Xwire900 net901 VGND VGND VPWR VPWR net900 sky130_fd_sc_hd__buf_1
XFILLER_0_14_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23579_ _03425_ _03445_ VGND VGND VPWR VPWR _03447_ sky130_fd_sc_hd__nand2_1
Xwire911 _05890_ VGND VGND VPWR VPWR net911 sky130_fd_sc_hd__clkbuf_1
Xwire922 net923 VGND VGND VPWR VPWR net922 sky130_fd_sc_hd__clkbuf_1
Xwire933 _03543_ VGND VGND VPWR VPWR net933 sky130_fd_sc_hd__buf_1
X_16120_ net1091 _08185_ VGND VGND VPWR VPWR _08186_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_187_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13332_ net845 _05604_ VGND VGND VPWR VPWR _05605_ sky130_fd_sc_hd__xnor2_1
Xwire944 _02201_ VGND VGND VPWR VPWR net944 sky130_fd_sc_hd__clkbuf_4
X_25318_ clknet_leaf_75_clk _00201_ net8463 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.f\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire955 _11623_ VGND VGND VPWR VPWR net955 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire966 _08993_ VGND VGND VPWR VPWR net966 sky130_fd_sc_hd__buf_1
Xwire977 _08444_ VGND VGND VPWR VPWR net977 sky130_fd_sc_hd__clkbuf_1
Xwire988 net989 VGND VGND VPWR VPWR net988 sky130_fd_sc_hd__buf_1
X_16051_ _08114_ _08117_ VGND VGND VPWR VPWR _08118_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_161_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13263_ _05528_ _05535_ VGND VGND VPWR VPWR _05536_ sky130_fd_sc_hd__xnor2_2
X_25249_ clknet_leaf_87_clk _00132_ net8442 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.a\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire999 _05447_ VGND VGND VPWR VPWR net999 sky130_fd_sc_hd__buf_1
XFILLER_0_122_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15002_ _07038_ net3558 VGND VGND VPWR VPWR _07076_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13194_ _05382_ net849 VGND VGND VPWR VPWR _05467_ sky130_fd_sc_hd__nor2_1
Xwire4251 net4252 VGND VGND VPWR VPWR net4251 sky130_fd_sc_hd__clkbuf_1
X_19810_ net2506 _11643_ VGND VGND VPWR VPWR _11644_ sky130_fd_sc_hd__xnor2_1
Xwire4262 net4263 VGND VGND VPWR VPWR net4262 sky130_fd_sc_hd__clkbuf_1
Xwire4273 net4274 VGND VGND VPWR VPWR net4273 sky130_fd_sc_hd__clkbuf_1
Xwire4284 net4285 VGND VGND VPWR VPWR net4284 sky130_fd_sc_hd__buf_1
Xwire3550 net3551 VGND VGND VPWR VPWR net3550 sky130_fd_sc_hd__buf_1
Xwire4295 net4296 VGND VGND VPWR VPWR net4295 sky130_fd_sc_hd__clkbuf_1
X_19741_ net3157 _11522_ _11575_ VGND VGND VPWR VPWR _11576_ sky130_fd_sc_hd__o21a_1
X_16953_ net1814 VGND VGND VPWR VPWR _08916_ sky130_fd_sc_hd__buf_1
Xwire3561 _07035_ VGND VGND VPWR VPWR net3561 sky130_fd_sc_hd__buf_1
XFILLER_0_194_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3572 _07028_ VGND VGND VPWR VPWR net3572 sky130_fd_sc_hd__buf_1
Xwire3583 _07019_ VGND VGND VPWR VPWR net3583 sky130_fd_sc_hd__buf_1
Xwire3594 net3595 VGND VGND VPWR VPWR net3594 sky130_fd_sc_hd__buf_1
XFILLER_0_159_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15904_ _07971_ _07972_ net3546 net3392 VGND VGND VPWR VPWR _07973_ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19672_ net6156 _11506_ _11507_ _11336_ VGND VGND VPWR VPWR _11508_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_95_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16884_ net6344 net6325 net6309 net6277 net6518 net6498 VGND VGND VPWR VPWR _08848_
+ sky130_fd_sc_hd__mux4_1
Xwire2871 _06814_ VGND VGND VPWR VPWR net2871 sky130_fd_sc_hd__buf_1
XFILLER_0_155_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2893 _06569_ VGND VGND VPWR VPWR net2893 sky130_fd_sc_hd__buf_1
XFILLER_0_21_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18623_ net6929 _10431_ _10468_ _10469_ VGND VGND VPWR VPWR _10470_ sky130_fd_sc_hd__a31o_1
X_15835_ _07894_ _07904_ VGND VGND VPWR VPWR _07905_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_29_clk clknet_4_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_189_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18554_ net1438 net382 VGND VGND VPWR VPWR _10403_ sky130_fd_sc_hd__nor2_1
X_15766_ _07769_ _07835_ VGND VGND VPWR VPWR _07836_ sky130_fd_sc_hd__xnor2_1
X_12978_ net7748 _05012_ VGND VGND VPWR VPWR _05251_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17505_ net6703 VGND VGND VPWR VPWR _09392_ sky130_fd_sc_hd__inv_2
X_14717_ net9092 net2861 net2865 net1118 VGND VGND VPWR VPWR _00148_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18485_ net6378 VGND VGND VPWR VPWR _10335_ sky130_fd_sc_hd__inv_2
X_15697_ net2676 _07672_ _07767_ VGND VGND VPWR VPWR _07768_ sky130_fd_sc_hd__o21a_1
X_17436_ net4035 _09333_ VGND VGND VPWR VPWR _09334_ sky130_fd_sc_hd__nor2_1
XFILLER_0_170_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14648_ net8961 _06801_ _06808_ VGND VGND VPWR VPWR _00128_ sky130_fd_sc_hd__a21o_1
XFILLER_0_184_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17367_ net7377 svm0.delta\[1\] net2573 net667 VGND VGND VPWR VPWR _09279_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_16_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14579_ _06753_ _06754_ VGND VGND VPWR VPWR _06755_ sky130_fd_sc_hd__xor2_1
X_19106_ net6336 net6359 VGND VGND VPWR VPWR _10943_ sky130_fd_sc_hd__and2_1
X_16318_ net571 VGND VGND VPWR VPWR _08381_ sky130_fd_sc_hd__inv_2
X_17298_ net7702 _09211_ VGND VGND VPWR VPWR _09212_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19037_ _10872_ _10873_ net6178 net6220 net6115 VGND VGND VPWR VPWR _10874_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16249_ net2651 _08312_ VGND VGND VPWR VPWR _08313_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout5380 net5381 VGND VGND VPWR VPWR net5380 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout5391 net5398 VGND VGND VPWR VPWR net5391 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19939_ _11768_ net1408 VGND VGND VPWR VPWR _11771_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_195_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22950_ _02279_ net552 _02514_ net336 VGND VGND VPWR VPWR _02838_ sky130_fd_sc_hd__a211o_1
X_21901_ _01908_ _01812_ _01909_ VGND VGND VPWR VPWR _01910_ sky130_fd_sc_hd__a21o_1
X_22881_ _02776_ VGND VGND VPWR VPWR _00639_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24620_ net4843 VGND VGND VPWR VPWR _04475_ sky130_fd_sc_hd__inv_2
X_21832_ _01837_ _01840_ VGND VGND VPWR VPWR _01841_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24551_ _04357_ _04361_ _04406_ VGND VGND VPWR VPWR _04407_ sky130_fd_sc_hd__a21o_1
X_21763_ net5768 net5502 _01771_ _01772_ VGND VGND VPWR VPWR _01773_ sky130_fd_sc_hd__a31o_1
XFILLER_0_144_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23502_ _03254_ _03259_ _03260_ VGND VGND VPWR VPWR _03371_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_175_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20714_ net6023 net2284 _12485_ VGND VGND VPWR VPWR _12487_ sky130_fd_sc_hd__or3_1
XFILLER_0_77_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8506 net8507 VGND VGND VPWR VPWR net8506 sky130_fd_sc_hd__buf_1
X_24482_ net1651 _04338_ net2018 VGND VGND VPWR VPWR _04339_ sky130_fd_sc_hd__o21ai_2
X_21694_ _01703_ _01704_ VGND VGND VPWR VPWR _01705_ sky130_fd_sc_hd__and2b_1
XFILLER_0_19_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8528 net8518 VGND VGND VPWR VPWR net8528 sky130_fd_sc_hd__clkbuf_1
Xwire8539 net8540 VGND VGND VPWR VPWR net8539 sky130_fd_sc_hd__buf_1
X_23433_ _03200_ _03229_ _03302_ VGND VGND VPWR VPWR _03303_ sky130_fd_sc_hd__o21a_1
Xmax_length4237 _06503_ VGND VGND VPWR VPWR net4237 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20645_ net2190 _12423_ VGND VGND VPWR VPWR _12424_ sky130_fd_sc_hd__or2_1
Xwire7816 net7817 VGND VGND VPWR VPWR net7816 sky130_fd_sc_hd__clkbuf_1
Xmax_length3503 _07101_ VGND VGND VPWR VPWR net3503 sky130_fd_sc_hd__buf_1
Xwire207 _10780_ VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__buf_1
Xwire7838 net7839 VGND VGND VPWR VPWR net7838 sky130_fd_sc_hd__clkbuf_1
Xwire229 _04632_ VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__clkbuf_1
X_23364_ _02932_ _02963_ _03233_ VGND VGND VPWR VPWR _03234_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7849 net7850 VGND VGND VPWR VPWR net7849 sky130_fd_sc_hd__buf_1
XFILLER_0_116_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2802 net2803 VGND VGND VPWR VPWR net2802 sky130_fd_sc_hd__buf_1
X_20576_ net1398 _12359_ net8056 VGND VGND VPWR VPWR _12360_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25103_ net4393 net5169 VGND VGND VPWR VPWR _04846_ sky130_fd_sc_hd__xor2_1
X_22315_ _02237_ _02240_ net756 VGND VGND VPWR VPWR _02319_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_15_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23295_ _03163_ _03164_ VGND VGND VPWR VPWR _03165_ sky130_fd_sc_hd__and2_1
XFILLER_0_61_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2879 net2880 VGND VGND VPWR VPWR net2879 sky130_fd_sc_hd__buf_1
X_22246_ _02248_ _02250_ VGND VGND VPWR VPWR _02251_ sky130_fd_sc_hd__nand2_1
X_25034_ net7473 net2396 VGND VGND VPWR VPWR _04787_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22177_ pid_d.prev_int\[10\] VGND VGND VPWR VPWR _02182_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2101 net2102 VGND VGND VPWR VPWR net2101 sky130_fd_sc_hd__buf_1
X_21128_ _01122_ _01124_ _01140_ _01142_ _01143_ VGND VGND VPWR VPWR _01144_ sky130_fd_sc_hd__a221o_1
Xwire2112 _10951_ VGND VGND VPWR VPWR net2112 sky130_fd_sc_hd__buf_1
Xwire2123 net2124 VGND VGND VPWR VPWR net2123 sky130_fd_sc_hd__buf_1
Xwire2134 net2135 VGND VGND VPWR VPWR net2134 sky130_fd_sc_hd__buf_1
Xwire1400 net1401 VGND VGND VPWR VPWR net1400 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2145 _09692_ VGND VGND VPWR VPWR net2145 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2156 net2158 VGND VGND VPWR VPWR net2156 sky130_fd_sc_hd__buf_1
Xwire1411 _11753_ VGND VGND VPWR VPWR net1411 sky130_fd_sc_hd__clkbuf_1
X_13950_ _06158_ _06215_ VGND VGND VPWR VPWR _06216_ sky130_fd_sc_hd__xnor2_1
X_25936_ clknet_4_7__leaf_clk _00015_ net8581 VGND VGND VPWR VPWR pid_d.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
Xwire1422 net1423 VGND VGND VPWR VPWR net1422 sky130_fd_sc_hd__buf_1
Xwire2167 net2168 VGND VGND VPWR VPWR net2167 sky130_fd_sc_hd__clkbuf_1
X_21059_ _01029_ _01065_ _01074_ VGND VGND VPWR VPWR _01075_ sky130_fd_sc_hd__a21o_1
Xwire2178 net2179 VGND VGND VPWR VPWR net2178 sky130_fd_sc_hd__buf_1
Xwire1433 net1434 VGND VGND VPWR VPWR net1433 sky130_fd_sc_hd__buf_1
Xwire1444 net1445 VGND VGND VPWR VPWR net1444 sky130_fd_sc_hd__buf_1
Xwire2189 _08833_ VGND VGND VPWR VPWR net2189 sky130_fd_sc_hd__buf_1
Xwire1455 _09579_ VGND VGND VPWR VPWR net1455 sky130_fd_sc_hd__buf_1
X_12901_ _05170_ _05173_ VGND VGND VPWR VPWR _05174_ sky130_fd_sc_hd__xnor2_1
Xwire1466 net1467 VGND VGND VPWR VPWR net1466 sky130_fd_sc_hd__clkbuf_1
X_13881_ net449 _06144_ _06147_ VGND VGND VPWR VPWR _06148_ sky130_fd_sc_hd__a21bo_1
X_25867_ clknet_leaf_16_clk _00740_ net8625 VGND VGND VPWR VPWR pid_q.mult0.a\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1477 _09057_ VGND VGND VPWR VPWR net1477 sky130_fd_sc_hd__clkbuf_1
Xwire1488 net1489 VGND VGND VPWR VPWR net1488 sky130_fd_sc_hd__clkbuf_1
Xwire1499 net1500 VGND VGND VPWR VPWR net1499 sky130_fd_sc_hd__clkbuf_1
X_15620_ net4075 net4074 VGND VGND VPWR VPWR _07692_ sky130_fd_sc_hd__or2_1
X_24818_ net9164 net1644 _04542_ net175 VGND VGND VPWR VPWR _00712_ sky130_fd_sc_hd__a22o_1
X_12832_ net7848 _04962_ net2971 VGND VGND VPWR VPWR _05105_ sky130_fd_sc_hd__and3_1
X_25798_ clknet_leaf_32_clk _00671_ net8683 VGND VGND VPWR VPWR pid_q.curr_int\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_97_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15551_ net1109 _07623_ VGND VGND VPWR VPWR _07624_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24749_ _04578_ _04579_ net4232 VGND VGND VPWR VPWR _04580_ sky130_fd_sc_hd__a21o_1
X_12763_ net7804 net2354 net2316 VGND VGND VPWR VPWR _05036_ sky130_fd_sc_hd__and3_2
XFILLER_0_16_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14502_ _06679_ _06681_ _06680_ VGND VGND VPWR VPWR _06684_ sky130_fd_sc_hd__o21ba_1
X_18270_ _09176_ _10065_ VGND VGND VPWR VPWR _10121_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15482_ _07341_ _07471_ _07472_ net675 VGND VGND VPWR VPWR _07556_ sky130_fd_sc_hd__a211o_1
X_12694_ _04961_ _04966_ VGND VGND VPWR VPWR _04967_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17221_ net6788 _09168_ _09169_ VGND VGND VPWR VPWR _00340_ sky130_fd_sc_hd__a21bo_1
X_14433_ net5219 net1294 net2890 net4419 _06628_ VGND VGND VPWR VPWR _06629_ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17152_ net6914 _09086_ _09104_ _09105_ VGND VGND VPWR VPWR _09106_ sky130_fd_sc_hd__o211a_1
Xwire730 _05697_ VGND VGND VPWR VPWR net730 sky130_fd_sc_hd__clkbuf_1
X_14364_ net8305 net3636 VGND VGND VPWR VPWR _06576_ sky130_fd_sc_hd__and2_1
Xinput15 angle_in[8] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_1
Xwire741 net742 VGND VGND VPWR VPWR net741 sky130_fd_sc_hd__clkbuf_1
Xinput26 currA_in[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
Xwire752 net753 VGND VGND VPWR VPWR net752 sky130_fd_sc_hd__clkbuf_1
Xmax_length4793 net4794 VGND VGND VPWR VPWR net4793 sky130_fd_sc_hd__buf_1
Xinput37 currB_in[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
Xwire763 _11117_ VGND VGND VPWR VPWR net763 sky130_fd_sc_hd__clkbuf_1
X_16103_ net1526 net1515 _08166_ _08168_ net2640 VGND VGND VPWR VPWR _08169_ sky130_fd_sc_hd__a32o_1
Xinput48 currB_in[9] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_1
Xinput59 currT_in[4] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_1
X_13315_ _05584_ _05587_ VGND VGND VPWR VPWR _05588_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17083_ net7008 _09012_ VGND VGND VPWR VPWR _09041_ sky130_fd_sc_hd__nand2_1
Xmax_length350 net351 VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__buf_1
Xwire774 net775 VGND VGND VPWR VPWR net774 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire785 net786 VGND VGND VPWR VPWR net785 sky130_fd_sc_hd__clkbuf_1
X_14295_ net69 net2901 net2264 net7649 VGND VGND VPWR VPWR _00064_ sky130_fd_sc_hd__a22o_1
Xwire796 net797 VGND VGND VPWR VPWR net796 sky130_fd_sc_hd__buf_1
X_16034_ _08099_ _08100_ _07932_ VGND VGND VPWR VPWR _08101_ sky130_fd_sc_hd__a21oi_1
X_13246_ net7808 net2309 net1954 VGND VGND VPWR VPWR _05519_ sky130_fd_sc_hd__and3_1
XFILLER_0_161_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13177_ net7740 net1353 VGND VGND VPWR VPWR _05450_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4070 _07683_ VGND VGND VPWR VPWR net4070 sky130_fd_sc_hd__clkbuf_1
Xwire4081 net4082 VGND VGND VPWR VPWR net4081 sky130_fd_sc_hd__buf_1
Xwire4092 net4093 VGND VGND VPWR VPWR net4092 sky130_fd_sc_hd__buf_1
X_17985_ net3245 _09835_ VGND VGND VPWR VPWR _09836_ sky130_fd_sc_hd__nand2_1
Xwire3380 net3381 VGND VGND VPWR VPWR net3380 sky130_fd_sc_hd__clkbuf_2
X_16936_ cordic0.slte0.opA\[16\] VGND VGND VPWR VPWR _08900_ sky130_fd_sc_hd__inv_2
X_19724_ net6080 net6062 VGND VGND VPWR VPWR _11559_ sky130_fd_sc_hd__nor2b_1
Xwire3391 _07847_ VGND VGND VPWR VPWR net3391 sky130_fd_sc_hd__clkbuf_1
Xwire2690 _07505_ VGND VGND VPWR VPWR net2690 sky130_fd_sc_hd__clkbuf_1
X_16867_ net6483 VGND VGND VPWR VPWR _08832_ sky130_fd_sc_hd__inv_2
X_19655_ net3133 net3863 VGND VGND VPWR VPWR _11491_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_9_Left_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15818_ _07878_ _07887_ VGND VGND VPWR VPWR _07888_ sky130_fd_sc_hd__xnor2_2
X_18606_ net1196 _10452_ VGND VGND VPWR VPWR _10454_ sky130_fd_sc_hd__nor2_1
X_19586_ _11419_ _11422_ VGND VGND VPWR VPWR _11423_ sky130_fd_sc_hd__nand2_1
X_16798_ cordic0.cos\[2\] matmul0.cos\[2\] net3370 VGND VGND VPWR VPWR _08789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18537_ _10322_ net1205 _10385_ VGND VGND VPWR VPWR _10386_ sky130_fd_sc_hd__a21oi_1
X_15749_ _07712_ _07732_ _07710_ VGND VGND VPWR VPWR _07820_ sky130_fd_sc_hd__o21a_1
X_18468_ net3284 net3225 VGND VGND VPWR VPWR _10318_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17419_ net3276 _09320_ VGND VGND VPWR VPWR _09321_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18399_ net6854 net6811 net6774 net1775 VGND VGND VPWR VPWR _10250_ sky130_fd_sc_hd__a31o_1
XFILLER_0_133_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20430_ net2596 net2166 VGND VGND VPWR VPWR _12225_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20361_ net1399 _12161_ net8041 VGND VGND VPWR VPWR _12162_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_9_clk clknet_4_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22100_ net4383 _02021_ net343 net4319 net522 VGND VGND VPWR VPWR _02107_ sky130_fd_sc_hd__a221o_1
XFILLER_0_67_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23080_ net5001 net4685 VGND VGND VPWR VPWR _02950_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20292_ net6468 net1486 VGND VGND VPWR VPWR _12098_ sky130_fd_sc_hd__nand2_2
X_22031_ _01932_ _01937_ _02037_ VGND VGND VPWR VPWR _02038_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23982_ _03837_ _03845_ VGND VGND VPWR VPWR _03846_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25721_ clknet_leaf_13_clk _00594_ net8603 VGND VGND VPWR VPWR pid_d.mult0.a\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_22933_ _02813_ _02820_ _02821_ VGND VGND VPWR VPWR _02823_ sky130_fd_sc_hd__nand3_1
XFILLER_0_155_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25652_ clknet_leaf_1_clk _00525_ net8401 VGND VGND VPWR VPWR pid_d.curr_int\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_196_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22864_ net5981 _02747_ _02751_ net5980 VGND VGND VPWR VPWR _02761_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24603_ _04390_ _04456_ _04457_ VGND VGND VPWR VPWR _04458_ sky130_fd_sc_hd__o21a_1
X_21815_ net600 _01631_ _01632_ _01724_ VGND VGND VPWR VPWR _01824_ sky130_fd_sc_hd__a211o_1
XFILLER_0_196_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25583_ clknet_leaf_90_clk _00456_ net8422 VGND VGND VPWR VPWR cordic0.cos\[3\] sky130_fd_sc_hd__dfrtp_1
X_22795_ _02705_ VGND VGND VPWR VPWR _00624_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24534_ _04331_ _04336_ _04332_ VGND VGND VPWR VPWR _04390_ sky130_fd_sc_hd__a21boi_1
X_21746_ net5742 net5500 VGND VGND VPWR VPWR _01756_ sky130_fd_sc_hd__nand2_1
Xfanout7507 net7516 VGND VGND VPWR VPWR net7507 sky130_fd_sc_hd__buf_1
Xmax_length4001 _09581_ VGND VGND VPWR VPWR net4001 sky130_fd_sc_hd__buf_1
Xwire8303 net8304 VGND VGND VPWR VPWR net8303 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8314 net8315 VGND VGND VPWR VPWR net8314 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8325 net8326 VGND VGND VPWR VPWR net8325 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8336 net8337 VGND VGND VPWR VPWR net8336 sky130_fd_sc_hd__buf_1
XFILLER_0_53_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7602 net7603 VGND VGND VPWR VPWR net7602 sky130_fd_sc_hd__buf_1
X_24465_ _04321_ _04322_ VGND VGND VPWR VPWR _04323_ sky130_fd_sc_hd__nand2_1
XFILLER_0_191_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7613 net7611 VGND VGND VPWR VPWR net7613 sky130_fd_sc_hd__buf_1
XFILLER_0_149_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21677_ _01586_ _01587_ _01585_ VGND VGND VPWR VPWR _01688_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4045 net4046 VGND VGND VPWR VPWR net4045 sky130_fd_sc_hd__buf_1
Xwire8358 net8357 VGND VGND VPWR VPWR net8358 sky130_fd_sc_hd__buf_1
Xmax_length3311 net3312 VGND VGND VPWR VPWR net3311 sky130_fd_sc_hd__buf_1
Xwire7624 svm0.periodTop\[15\] VGND VGND VPWR VPWR net7624 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout6828 net6832 VGND VGND VPWR VPWR net6828 sky130_fd_sc_hd__clkbuf_2
X_23416_ _03284_ _03285_ VGND VGND VPWR VPWR _03286_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout6839 net6843 VGND VGND VPWR VPWR net6839 sky130_fd_sc_hd__buf_1
Xmax_length3333 _08971_ VGND VGND VPWR VPWR net3333 sky130_fd_sc_hd__buf_1
X_20628_ net6755 _12407_ net3305 VGND VGND VPWR VPWR _12408_ sky130_fd_sc_hd__mux2_1
Xwire7657 net7658 VGND VGND VPWR VPWR net7657 sky130_fd_sc_hd__clkbuf_1
X_24396_ _04253_ _04254_ VGND VGND VPWR VPWR _04255_ sky130_fd_sc_hd__nand2_1
Xwire6912 net6913 VGND VGND VPWR VPWR net6912 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_190_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2610 _08925_ VGND VGND VPWR VPWR net2610 sky130_fd_sc_hd__buf_1
Xwire7668 net7669 VGND VGND VPWR VPWR net7668 sky130_fd_sc_hd__clkbuf_1
Xmax_length3366 _08803_ VGND VGND VPWR VPWR net3366 sky130_fd_sc_hd__clkbuf_2
Xwire6934 net6932 VGND VGND VPWR VPWR net6934 sky130_fd_sc_hd__buf_1
XFILLER_0_85_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23347_ net4941 net4707 VGND VGND VPWR VPWR _03217_ sky130_fd_sc_hd__nand2_2
X_20559_ net1745 _12343_ VGND VGND VPWR VPWR _12344_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_34_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3377 _08781_ VGND VGND VPWR VPWR net3377 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6956 net6957 VGND VGND VPWR VPWR net6956 sky130_fd_sc_hd__buf_1
Xmax_length2643 net2644 VGND VGND VPWR VPWR net2643 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13100_ net7757 net1620 VGND VGND VPWR VPWR _05373_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14080_ net4250 _05351_ VGND VGND VPWR VPWR _06343_ sky130_fd_sc_hd__nor2_1
Xwire6989 net6992 VGND VGND VPWR VPWR net6989 sky130_fd_sc_hd__buf_2
X_23278_ _02990_ _03002_ VGND VGND VPWR VPWR _03148_ sky130_fd_sc_hd__xor2_1
Xmax_length2698 _07489_ VGND VGND VPWR VPWR net2698 sky130_fd_sc_hd__clkbuf_1
Xmax_length1964 net1965 VGND VGND VPWR VPWR net1964 sky130_fd_sc_hd__clkbuf_1
X_25017_ net7471 _04770_ _04771_ net7497 net467 VGND VGND VPWR VPWR _04772_ sky130_fd_sc_hd__a32o_1
X_13031_ _05284_ _05303_ VGND VGND VPWR VPWR _05304_ sky130_fd_sc_hd__xor2_1
X_22229_ net1389 _02145_ _02135_ VGND VGND VPWR VPWR _02234_ sky130_fd_sc_hd__a21bo_1
Xmax_length1997 net1998 VGND VGND VPWR VPWR net1997 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17770_ net7140 _09618_ net3261 VGND VGND VPWR VPWR _09621_ sky130_fd_sc_hd__a21boi_1
X_14982_ net3603 _07055_ VGND VGND VPWR VPWR _07056_ sky130_fd_sc_hd__nor2_1
Xwire1230 net1231 VGND VGND VPWR VPWR net1230 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1241 _08690_ VGND VGND VPWR VPWR net1241 sky130_fd_sc_hd__clkbuf_1
X_16721_ matmul0.matmul_stage_inst.mult2\[14\] matmul0.matmul_stage_inst.mult1\[14\]
+ VGND VGND VPWR VPWR _08747_ sky130_fd_sc_hd__nor2_1
X_13933_ _06120_ _06122_ VGND VGND VPWR VPWR _06199_ sky130_fd_sc_hd__nand2_1
X_25919_ clknet_leaf_28_clk _00792_ net8656 VGND VGND VPWR VPWR pid_q.out\[15\] sky130_fd_sc_hd__dfrtp_1
Xwire1263 _07903_ VGND VGND VPWR VPWR net1263 sky130_fd_sc_hd__buf_1
XFILLER_0_191_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1274 _07356_ VGND VGND VPWR VPWR net1274 sky130_fd_sc_hd__clkbuf_2
X_19440_ _10983_ _10796_ net6209 VGND VGND VPWR VPWR _11277_ sky130_fd_sc_hd__o21a_1
Xwire1285 _07105_ VGND VGND VPWR VPWR net1285 sky130_fd_sc_hd__buf_1
XFILLER_0_92_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1296 net1297 VGND VGND VPWR VPWR net1296 sky130_fd_sc_hd__buf_1
X_16652_ _08686_ _08682_ _08687_ VGND VGND VPWR VPWR _08688_ sky130_fd_sc_hd__a21o_1
X_13864_ net7788 net1318 _06129_ _06130_ VGND VGND VPWR VPWR _06131_ sky130_fd_sc_hd__a22o_1
X_15603_ net2687 _07670_ _07593_ VGND VGND VPWR VPWR _07675_ sky130_fd_sc_hd__a21o_1
X_12815_ _05072_ _05087_ _05077_ VGND VGND VPWR VPWR _05088_ sky130_fd_sc_hd__a21oi_1
X_19371_ net6152 _11207_ VGND VGND VPWR VPWR _11208_ sky130_fd_sc_hd__nand2_1
X_16583_ matmul0.matmul_stage_inst.mult2\[2\] net433 net2619 VGND VGND VPWR VPWR _08639_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13795_ _06051_ net840 VGND VGND VPWR VPWR _06063_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18322_ net6892 net6872 _10102_ VGND VGND VPWR VPWR _10173_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15534_ _07605_ _07606_ VGND VGND VPWR VPWR _07607_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12746_ _05008_ _05010_ _05018_ VGND VGND VPWR VPWR _05019_ sky130_fd_sc_hd__o21ba_1
Xfanout8731 net8827 VGND VGND VPWR VPWR net8731 sky130_fd_sc_hd__buf_1
XFILLER_0_56_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18253_ net6872 net3932 VGND VGND VPWR VPWR _10104_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_166_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15465_ net1538 _07538_ VGND VGND VPWR VPWR _07539_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_72_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12677_ net7915 net2368 net2365 VGND VGND VPWR VPWR _04950_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout8786 net8791 VGND VGND VPWR VPWR net8786 sky130_fd_sc_hd__buf_1
X_17204_ net1815 _09153_ net4245 VGND VGND VPWR VPWR _09154_ sky130_fd_sc_hd__a21o_1
X_14416_ net8136 net3632 VGND VGND VPWR VPWR _06616_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8870 net8871 VGND VGND VPWR VPWR net8870 sky130_fd_sc_hd__buf_1
XFILLER_0_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18184_ net7142 _10034_ _09630_ VGND VGND VPWR VPWR _10035_ sky130_fd_sc_hd__or3b_1
Xwire8881 net134 VGND VGND VPWR VPWR net8881 sky130_fd_sc_hd__clkbuf_1
X_15396_ _07219_ _07265_ VGND VGND VPWR VPWR _07470_ sky130_fd_sc_hd__xor2_1
Xwire8892 net8894 VGND VGND VPWR VPWR net8892 sky130_fd_sc_hd__buf_1
X_17135_ net2181 _09089_ net3322 VGND VGND VPWR VPWR _09090_ sky130_fd_sc_hd__a21o_1
XFILLER_0_163_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire560 net561 VGND VGND VPWR VPWR net560 sky130_fd_sc_hd__clkbuf_1
X_14347_ _06562_ VGND VGND VPWR VPWR _00073_ sky130_fd_sc_hd__clkbuf_1
Xwire571 _08380_ VGND VGND VPWR VPWR net571 sky130_fd_sc_hd__clkbuf_2
Xwire582 _05666_ VGND VGND VPWR VPWR net582 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire593 net594 VGND VGND VPWR VPWR net593 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17066_ net1918 _09022_ VGND VGND VPWR VPWR _09025_ sky130_fd_sc_hd__nor2_1
X_14278_ net54 net2914 _06517_ net8990 VGND VGND VPWR VPWR _00049_ sky130_fd_sc_hd__a22o_1
X_16017_ net425 _08084_ _08008_ VGND VGND VPWR VPWR _08085_ sky130_fd_sc_hd__a21o_1
X_13229_ _05456_ _05461_ _05454_ VGND VGND VPWR VPWR _05502_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17968_ net6924 net6884 net4036 VGND VGND VPWR VPWR _09819_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19707_ _11488_ _11542_ VGND VGND VPWR VPWR _11543_ sky130_fd_sc_hd__nand2_1
X_16919_ _08864_ _08870_ _08878_ net2611 VGND VGND VPWR VPWR _08883_ sky130_fd_sc_hd__a211o_1
X_17899_ net7060 _09749_ VGND VGND VPWR VPWR _09750_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_178_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19638_ net3291 _11439_ _11473_ net1416 _11474_ VGND VGND VPWR VPWR _11475_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_178_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19569_ _11332_ _11338_ _11335_ VGND VGND VPWR VPWR _11406_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21600_ net5383 net3803 _01606_ _01611_ net5400 VGND VGND VPWR VPWR _01612_ sky130_fd_sc_hd__a32o_1
X_22580_ net4390 pid_d.state\[1\] net4315 net4326 VGND VGND VPWR VPWR _02560_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21531_ pid_d.curr_int\[4\] pid_d.prev_int\[4\] VGND VGND VPWR VPWR _01543_ sky130_fd_sc_hd__xor2_1
X_24250_ _04109_ _04031_ _04110_ VGND VGND VPWR VPWR _04111_ sky130_fd_sc_hd__o21a_1
XFILLER_0_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21462_ _01472_ _01474_ VGND VGND VPWR VPWR _01475_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6208 net6209 VGND VGND VPWR VPWR net6208 sky130_fd_sc_hd__buf_1
XFILLER_0_172_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6219 net6215 VGND VGND VPWR VPWR net6219 sky130_fd_sc_hd__buf_1
X_23201_ _03046_ _03047_ _03068_ VGND VGND VPWR VPWR _03071_ sky130_fd_sc_hd__or3b_1
X_20413_ cordic0.slte0.opA\[9\] _12198_ _12208_ _12209_ VGND VGND VPWR VPWR _12210_
+ sky130_fd_sc_hd__o211a_1
X_24181_ _04040_ _04041_ VGND VGND VPWR VPWR _04042_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21393_ _01404_ _01406_ net3117 VGND VGND VPWR VPWR _01407_ sky130_fd_sc_hd__a21o_1
Xwire5507 net5508 VGND VGND VPWR VPWR net5507 sky130_fd_sc_hd__buf_1
Xwire5518 net5512 VGND VGND VPWR VPWR net5518 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5529 net5530 VGND VGND VPWR VPWR net5529 sky130_fd_sc_hd__clkbuf_1
X_23132_ _02993_ net2431 _03001_ VGND VGND VPWR VPWR _03002_ sky130_fd_sc_hd__a21o_1
Xmax_length1227 _08991_ VGND VGND VPWR VPWR net1227 sky130_fd_sc_hd__clkbuf_1
X_20344_ net2591 _12090_ VGND VGND VPWR VPWR _12146_ sky130_fd_sc_hd__nor2_1
Xwire4817 net4818 VGND VGND VPWR VPWR net4817 sky130_fd_sc_hd__buf_1
Xwire4828 net4826 VGND VGND VPWR VPWR net4828 sky130_fd_sc_hd__buf_1
Xwire4839 net4829 VGND VGND VPWR VPWR net4839 sky130_fd_sc_hd__clkbuf_1
X_23063_ net5092 net4588 VGND VGND VPWR VPWR _02933_ sky130_fd_sc_hd__nand2_1
X_20275_ net7 cordic0.domain\[1\] net2533 VGND VGND VPWR VPWR _12083_ sky130_fd_sc_hd__mux2_1
X_22014_ _02019_ _02020_ VGND VGND VPWR VPWR _02021_ sky130_fd_sc_hd__xnor2_1
X_23965_ _03722_ _03727_ _03728_ VGND VGND VPWR VPWR _03829_ sky130_fd_sc_hd__a21oi_1
X_25704_ clknet_leaf_5_clk _00577_ net8567 VGND VGND VPWR VPWR pid_d.mult0.b\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_22916_ net8903 _02807_ VGND VGND VPWR VPWR _02808_ sky130_fd_sc_hd__and2_1
X_23896_ _03678_ _03760_ VGND VGND VPWR VPWR _03761_ sky130_fd_sc_hd__xor2_1
X_25635_ clknet_leaf_104_clk _00508_ net8361 VGND VGND VPWR VPWR cordic0.vec\[0\]\[7\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22847_ _02744_ _02734_ _02736_ _02745_ VGND VGND VPWR VPWR _02746_ sky130_fd_sc_hd__a31o_1
XFILLER_0_190_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12600_ net8864 net7463 VGND VGND VPWR VPWR _04879_ sky130_fd_sc_hd__and2_1
XFILLER_0_195_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13580_ _05849_ _05781_ VGND VGND VPWR VPWR _05851_ sky130_fd_sc_hd__or2b_1
XFILLER_0_38_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25566_ clknet_leaf_98_clk _00439_ net8387 VGND VGND VPWR VPWR cordic0.sin\[0\] sky130_fd_sc_hd__dfrtp_1
X_22778_ pid_d.kp\[1\] _02664_ net1679 VGND VGND VPWR VPWR _02697_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8100 net9 VGND VGND VPWR VPWR net8100 sky130_fd_sc_hd__buf_1
Xwire8111 net8112 VGND VGND VPWR VPWR net8111 sky130_fd_sc_hd__clkbuf_1
X_24517_ _04268_ net792 VGND VGND VPWR VPWR _04374_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21729_ pid_d.curr_int\[6\] pid_d.prev_int\[6\] VGND VGND VPWR VPWR _01739_ sky130_fd_sc_hd__xor2_1
X_25497_ clknet_leaf_42_clk _00377_ net8768 VGND VGND VPWR VPWR svm0.delta\[2\] sky130_fd_sc_hd__dfrtp_1
Xwire8133 net8134 VGND VGND VPWR VPWR net8133 sky130_fd_sc_hd__clkbuf_1
Xwire8144 net8145 VGND VGND VPWR VPWR net8144 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7410 matmul0.matmul_stage_inst.c\[8\] VGND VGND VPWR VPWR net7410 sky130_fd_sc_hd__clkbuf_1
Xwire8155 net8156 VGND VGND VPWR VPWR net8155 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8166 net8167 VGND VGND VPWR VPWR net8166 sky130_fd_sc_hd__clkbuf_1
X_15250_ _07315_ _07318_ _07323_ VGND VGND VPWR VPWR _07324_ sky130_fd_sc_hd__o21a_1
Xwire7421 net7422 VGND VGND VPWR VPWR net7421 sky130_fd_sc_hd__clkbuf_1
X_24448_ _04286_ _04305_ VGND VGND VPWR VPWR _04306_ sky130_fd_sc_hd__xor2_2
XFILLER_0_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7432 net7433 VGND VGND VPWR VPWR net7432 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8177 net8178 VGND VGND VPWR VPWR net8177 sky130_fd_sc_hd__clkbuf_1
Xmax_length3130 net3131 VGND VGND VPWR VPWR net3130 sky130_fd_sc_hd__buf_1
Xwire8188 net8189 VGND VGND VPWR VPWR net8188 sky130_fd_sc_hd__clkbuf_1
X_14201_ _06459_ _06460_ VGND VGND VPWR VPWR _06461_ sky130_fd_sc_hd__or2b_1
Xwire8199 net8200 VGND VGND VPWR VPWR net8199 sky130_fd_sc_hd__clkbuf_1
Xwire7454 net7453 VGND VGND VPWR VPWR net7454 sky130_fd_sc_hd__clkbuf_2
Xwire6720 net6721 VGND VGND VPWR VPWR net6720 sky130_fd_sc_hd__buf_1
Xwire7465 net7462 VGND VGND VPWR VPWR net7465 sky130_fd_sc_hd__clkbuf_2
Xwire6731 net6732 VGND VGND VPWR VPWR net6731 sky130_fd_sc_hd__clkbuf_1
Xwire7476 net7470 VGND VGND VPWR VPWR net7476 sky130_fd_sc_hd__clkbuf_1
X_15181_ _07237_ _07239_ _07254_ VGND VGND VPWR VPWR _07255_ sky130_fd_sc_hd__o21ai_2
Xwire6742 svm0.delta\[13\] VGND VGND VPWR VPWR net6742 sky130_fd_sc_hd__clkbuf_2
Xwire7487 net7488 VGND VGND VPWR VPWR net7487 sky130_fd_sc_hd__clkbuf_1
X_24379_ _04199_ _04237_ VGND VGND VPWR VPWR _04238_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7498 net7499 VGND VGND VPWR VPWR net7498 sky130_fd_sc_hd__buf_1
Xwire6753 net6754 VGND VGND VPWR VPWR net6753 sky130_fd_sc_hd__clkbuf_1
X_14132_ _06371_ _06393_ VGND VGND VPWR VPWR _06394_ sky130_fd_sc_hd__or2_2
Xmax_length3196 net3197 VGND VGND VPWR VPWR net3196 sky130_fd_sc_hd__clkbuf_1
Xwire6764 net6759 VGND VGND VPWR VPWR net6764 sky130_fd_sc_hd__buf_1
Xwire6775 net6776 VGND VGND VPWR VPWR net6775 sky130_fd_sc_hd__clkbuf_1
Xwire6786 net6787 VGND VGND VPWR VPWR net6786 sky130_fd_sc_hd__buf_1
XFILLER_0_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14063_ net1322 VGND VGND VPWR VPWR _06326_ sky130_fd_sc_hd__clkbuf_1
X_18940_ _10764_ _10765_ _10778_ VGND VGND VPWR VPWR _10779_ sky130_fd_sc_hd__a21oi_1
Xmax_length1772 _10264_ VGND VGND VPWR VPWR net1772 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_148_Right_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13014_ net5215 net3029 _05285_ _05286_ VGND VGND VPWR VPWR _05287_ sky130_fd_sc_hd__a31oi_4
X_18871_ _10369_ _10677_ _10708_ net6898 _10712_ VGND VGND VPWR VPWR _10713_ sky130_fd_sc_hd__a221o_1
X_17822_ _09629_ _09659_ _09672_ VGND VGND VPWR VPWR _09673_ sky130_fd_sc_hd__o21a_1
Xhold4 pid_d.curr_error\[5\] VGND VGND VPWR VPWR net8957 sky130_fd_sc_hd__dlygate4sd3_1
X_14965_ net4143 net4140 VGND VGND VPWR VPWR _07039_ sky130_fd_sc_hd__nor2_1
X_17753_ net7068 net7094 VGND VGND VPWR VPWR _09604_ sky130_fd_sc_hd__and2b_1
Xwire1060 _11316_ VGND VGND VPWR VPWR net1060 sky130_fd_sc_hd__clkbuf_2
Xwire1071 net1072 VGND VGND VPWR VPWR net1071 sky130_fd_sc_hd__clkbuf_2
X_13916_ _06173_ _06054_ net7610 VGND VGND VPWR VPWR _06182_ sky130_fd_sc_hd__o21bai_1
X_16704_ matmul0.alpha_pass\[12\] net353 net6557 VGND VGND VPWR VPWR _08733_ sky130_fd_sc_hd__mux2_1
Xwire1082 _08345_ VGND VGND VPWR VPWR net1082 sky130_fd_sc_hd__clkbuf_1
X_17684_ net6746 _09526_ net6710 VGND VGND VPWR VPWR _09564_ sky130_fd_sc_hd__o21ba_1
Xwire1093 _08113_ VGND VGND VPWR VPWR net1093 sky130_fd_sc_hd__dlymetal6s2s_1
X_14896_ net6543 net6588 net7396 VGND VGND VPWR VPWR _06970_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19423_ _11257_ _11259_ _10797_ VGND VGND VPWR VPWR _11260_ sky130_fd_sc_hd__mux2_1
X_16635_ matmul0.matmul_stage_inst.mult2\[2\] VGND VGND VPWR VPWR _08673_ sky130_fd_sc_hd__inv_2
XFILLER_0_187_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13847_ _06061_ _06113_ _06060_ VGND VGND VPWR VPWR _06114_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19354_ net6202 net6288 VGND VGND VPWR VPWR _11191_ sky130_fd_sc_hd__or2b_1
X_16566_ _08554_ _08623_ _08624_ VGND VGND VPWR VPWR _08625_ sky130_fd_sc_hd__o21a_1
X_13778_ _05943_ _05944_ _05950_ _05951_ VGND VGND VPWR VPWR _06046_ sky130_fd_sc_hd__a22o_1
XFILLER_0_186_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15517_ _07584_ _07589_ VGND VGND VPWR VPWR _07590_ sky130_fd_sc_hd__xnor2_2
X_18305_ _10154_ _10155_ VGND VGND VPWR VPWR _10156_ sky130_fd_sc_hd__xnor2_1
X_12729_ _04972_ _05001_ VGND VGND VPWR VPWR _05002_ sky130_fd_sc_hd__xor2_1
X_19285_ net3886 VGND VGND VPWR VPWR _11122_ sky130_fd_sc_hd__buf_1
XFILLER_0_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8561 net8564 VGND VGND VPWR VPWR net8561 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_73_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16497_ net2631 net2641 VGND VGND VPWR VPWR _08557_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18236_ net7142 net2554 _10037_ VGND VGND VPWR VPWR _10087_ sky130_fd_sc_hd__o21ai_1
X_15448_ _07513_ _07521_ VGND VGND VPWR VPWR _07522_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18167_ _10006_ _10008_ _10001_ VGND VGND VPWR VPWR _10018_ sky130_fd_sc_hd__a21o_1
X_15379_ net1878 net1275 VGND VGND VPWR VPWR _07453_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17118_ net1476 _09073_ net1221 VGND VGND VPWR VPWR _09074_ sky130_fd_sc_hd__o21ai_2
Xwire390 net391 VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__clkbuf_1
X_18098_ _09897_ _09948_ VGND VGND VPWR VPWR _09949_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17049_ net6486 net6464 VGND VGND VPWR VPWR _09008_ sky130_fd_sc_hd__or2_1
XFILLER_0_187_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_115_Right_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20060_ net3152 net3125 _11888_ VGND VGND VPWR VPWR _11889_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23750_ net4729 net4812 VGND VGND VPWR VPWR _03616_ sky130_fd_sc_hd__nand2_1
Xmax_length7407 matmul0.matmul_stage_inst.c\[10\] VGND VGND VPWR VPWR net7407 sky130_fd_sc_hd__clkbuf_1
X_20962_ net5924 VGND VGND VPWR VPWR _00978_ sky130_fd_sc_hd__inv_4
XFILLER_0_36_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22701_ _02642_ VGND VGND VPWR VPWR _00593_ sky130_fd_sc_hd__clkbuf_1
Xmax_length6717 svm0.counter\[7\] VGND VGND VPWR VPWR net6717 sky130_fd_sc_hd__clkbuf_2
X_23681_ net4768 net3746 VGND VGND VPWR VPWR _03548_ sky130_fd_sc_hd__or2_1
X_20893_ _00907_ _00908_ VGND VGND VPWR VPWR _00909_ sky130_fd_sc_hd__xnor2_1
X_25420_ clknet_leaf_98_clk _00303_ net8382 VGND VGND VPWR VPWR matmul0.cos\[7\] sky130_fd_sc_hd__dfrtp_1
X_22632_ _02560_ VGND VGND VPWR VPWR _02600_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_48_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25351_ clknet_leaf_83_clk _00234_ net8502 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22563_ net3768 net3093 VGND VGND VPWR VPWR _02547_ sky130_fd_sc_hd__and2_1
XFILLER_0_152_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24302_ _04123_ _04161_ VGND VGND VPWR VPWR _04162_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_161_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21514_ _01418_ _01525_ _01526_ VGND VGND VPWR VPWR _01527_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25282_ clknet_leaf_92_clk _00165_ net8429 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.c\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_22494_ _02429_ _02436_ _02431_ VGND VGND VPWR VPWR _02495_ sky130_fd_sc_hd__a21o_1
Xmax_length905 _06543_ VGND VGND VPWR VPWR net905 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6016 net6017 VGND VGND VPWR VPWR net6016 sky130_fd_sc_hd__clkbuf_1
X_24233_ net2022 net1656 VGND VGND VPWR VPWR _04094_ sky130_fd_sc_hd__xnor2_1
X_21445_ _01456_ _01457_ VGND VGND VPWR VPWR _01458_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6038 net6039 VGND VGND VPWR VPWR net6038 sky130_fd_sc_hd__buf_1
XFILLER_0_181_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6049 net6050 VGND VGND VPWR VPWR net6049 sky130_fd_sc_hd__buf_2
XFILLER_0_90_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5315 net5316 VGND VGND VPWR VPWR net5315 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5326 pid_d.out\[14\] VGND VGND VPWR VPWR net5326 sky130_fd_sc_hd__clkbuf_1
X_24164_ _04022_ net590 VGND VGND VPWR VPWR _04026_ sky130_fd_sc_hd__xnor2_1
Xwire5337 net5338 VGND VGND VPWR VPWR net5337 sky130_fd_sc_hd__clkbuf_1
X_21376_ _01263_ _01268_ _01389_ VGND VGND VPWR VPWR _01390_ sky130_fd_sc_hd__a21o_1
Xwire4603 net4604 VGND VGND VPWR VPWR net4603 sky130_fd_sc_hd__buf_1
Xwire5348 net5349 VGND VGND VPWR VPWR net5348 sky130_fd_sc_hd__clkbuf_1
Xwire4614 net4615 VGND VGND VPWR VPWR net4614 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5359 pid_d.out\[7\] VGND VGND VPWR VPWR net5359 sky130_fd_sc_hd__clkbuf_1
X_23115_ _02908_ _02919_ VGND VGND VPWR VPWR _02985_ sky130_fd_sc_hd__xor2_1
Xwire4625 net4626 VGND VGND VPWR VPWR net4625 sky130_fd_sc_hd__buf_1
X_20327_ _12129_ _12130_ _08885_ VGND VGND VPWR VPWR _12131_ sky130_fd_sc_hd__mux2_1
Xwire4636 net4637 VGND VGND VPWR VPWR net4636 sky130_fd_sc_hd__buf_1
Xwire4647 net4654 VGND VGND VPWR VPWR net4647 sky130_fd_sc_hd__buf_1
X_24095_ _03954_ net743 _03956_ VGND VGND VPWR VPWR _03957_ sky130_fd_sc_hd__a21o_1
Xwire3902 _10813_ VGND VGND VPWR VPWR net3902 sky130_fd_sc_hd__buf_1
Xwire4658 net4659 VGND VGND VPWR VPWR net4658 sky130_fd_sc_hd__clkbuf_1
Xwire3913 _10790_ VGND VGND VPWR VPWR net3913 sky130_fd_sc_hd__buf_1
Xwire3924 _10218_ VGND VGND VPWR VPWR net3924 sky130_fd_sc_hd__clkbuf_1
Xwire4669 net4670 VGND VGND VPWR VPWR net4669 sky130_fd_sc_hd__buf_1
X_23046_ _02897_ _02896_ VGND VGND VPWR VPWR _02916_ sky130_fd_sc_hd__xor2_1
X_20258_ _12070_ cordic0.slte0.opB\[12\] net2531 VGND VGND VPWR VPWR _12071_ sky130_fd_sc_hd__mux2_1
Xwire3935 _10064_ VGND VGND VPWR VPWR net3935 sky130_fd_sc_hd__clkbuf_1
Xwire3957 net3958 VGND VGND VPWR VPWR net3957 sky130_fd_sc_hd__clkbuf_1
Xwire3968 _09735_ VGND VGND VPWR VPWR net3968 sky130_fd_sc_hd__clkbuf_1
Xwire3979 net3980 VGND VGND VPWR VPWR net3979 sky130_fd_sc_hd__clkbuf_1
X_20189_ net244 _11967_ net3126 VGND VGND VPWR VPWR _12015_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24997_ net7498 net543 _04754_ net7472 VGND VGND VPWR VPWR _04755_ sky130_fd_sc_hd__a22o_1
X_14750_ net7454 _06835_ net7155 VGND VGND VPWR VPWR _06882_ sky130_fd_sc_hd__or3b_1
X_23948_ _03694_ _03696_ _03695_ VGND VGND VPWR VPWR _03812_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13701_ _05968_ _05969_ VGND VGND VPWR VPWR _05970_ sky130_fd_sc_hd__nor2_1
XFILLER_0_168_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14681_ net7156 _06830_ VGND VGND VPWR VPWR _06831_ sky130_fd_sc_hd__xor2_1
X_23879_ net4748 _03739_ net3049 VGND VGND VPWR VPWR _03744_ sky130_fd_sc_hd__or3b_1
X_16420_ net490 net571 VGND VGND VPWR VPWR _08482_ sky130_fd_sc_hd__or2_1
X_13632_ _05810_ _05811_ _05901_ VGND VGND VPWR VPWR _05902_ sky130_fd_sc_hd__a21o_1
X_25618_ clknet_leaf_110_clk _00491_ net8347 VGND VGND VPWR VPWR cordic0.slte0.opA\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_6_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16351_ net978 _08337_ _08333_ VGND VGND VPWR VPWR _08414_ sky130_fd_sc_hd__a21o_1
XFILLER_0_183_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13563_ net681 _05833_ VGND VGND VPWR VPWR _05834_ sky130_fd_sc_hd__xnor2_1
X_25549_ clknet_leaf_28_clk _00429_ net8649 VGND VGND VPWR VPWR pid_q.prev_int\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout7134 net7143 VGND VGND VPWR VPWR net7134 sky130_fd_sc_hd__buf_1
XFILLER_0_54_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15302_ _07372_ _07375_ VGND VGND VPWR VPWR _07376_ sky130_fd_sc_hd__xnor2_1
X_19070_ _10869_ _10889_ _10906_ VGND VGND VPWR VPWR _10907_ sky130_fd_sc_hd__a21o_1
X_16282_ _08185_ net1081 VGND VGND VPWR VPWR _08346_ sky130_fd_sc_hd__xor2_1
X_13494_ _05636_ _05650_ VGND VGND VPWR VPWR _05767_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7240 net7241 VGND VGND VPWR VPWR net7240 sky130_fd_sc_hd__clkbuf_1
X_18021_ net7052 _09641_ _09858_ _09870_ _09871_ VGND VGND VPWR VPWR _09872_ sky130_fd_sc_hd__a221o_1
Xwire7251 net7252 VGND VGND VPWR VPWR net7251 sky130_fd_sc_hd__clkbuf_1
Xfanout6444 state\[2\] VGND VGND VPWR VPWR net6444 sky130_fd_sc_hd__buf_1
X_15233_ net2711 net2797 net3443 _07306_ VGND VGND VPWR VPWR _07307_ sky130_fd_sc_hd__a31o_1
XFILLER_0_151_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6455 state\[0\] VGND VGND VPWR VPWR net6455 sky130_fd_sc_hd__buf_1
Xwire7262 net7263 VGND VGND VPWR VPWR net7262 sky130_fd_sc_hd__buf_1
Xwire7284 net7285 VGND VGND VPWR VPWR net7284 sky130_fd_sc_hd__buf_1
Xfanout6488 net6492 VGND VGND VPWR VPWR net6488 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7295 net7296 VGND VGND VPWR VPWR net7295 sky130_fd_sc_hd__clkbuf_1
Xwire6550 net6551 VGND VGND VPWR VPWR net6550 sky130_fd_sc_hd__buf_1
X_15164_ _07199_ net1892 VGND VGND VPWR VPWR _07238_ sky130_fd_sc_hd__xnor2_1
Xwire6561 net6562 VGND VGND VPWR VPWR net6561 sky130_fd_sc_hd__clkbuf_1
Xfanout5765 net5767 VGND VGND VPWR VPWR net5765 sky130_fd_sc_hd__buf_1
Xwire6583 net6580 VGND VGND VPWR VPWR net6583 sky130_fd_sc_hd__buf_1
X_14115_ _06349_ _06376_ VGND VGND VPWR VPWR _06377_ sky130_fd_sc_hd__xnor2_1
Xfanout5798 net5805 VGND VGND VPWR VPWR net5798 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5871 net5872 VGND VGND VPWR VPWR net5871 sky130_fd_sc_hd__clkbuf_1
X_19972_ net3153 net3199 net6027 net3880 VGND VGND VPWR VPWR _11803_ sky130_fd_sc_hd__o22a_1
X_15095_ _07125_ _07042_ VGND VGND VPWR VPWR _07169_ sky130_fd_sc_hd__nor2_1
Xmax_length1580 net1581 VGND VGND VPWR VPWR net1580 sky130_fd_sc_hd__buf_1
XFILLER_0_120_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14046_ _06246_ _06309_ VGND VGND VPWR VPWR _06310_ sky130_fd_sc_hd__xnor2_1
X_18923_ net3223 _10436_ net1427 _10762_ VGND VGND VPWR VPWR _10763_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_157_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18854_ net352 _10695_ VGND VGND VPWR VPWR _10697_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17805_ _09654_ _09655_ net7091 VGND VGND VPWR VPWR _09656_ sky130_fd_sc_hd__o21ai_1
X_15997_ net884 _07983_ VGND VGND VPWR VPWR _08065_ sky130_fd_sc_hd__and2_1
X_18785_ net1065 net1429 _10628_ VGND VGND VPWR VPWR _10629_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_167_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17736_ net8052 _09590_ _09591_ net6457 VGND VGND VPWR VPWR _00434_ sky130_fd_sc_hd__o2bb2a_1
X_14948_ net6620 net6640 matmul0.matmul_stage_inst.f\[8\] VGND VGND VPWR VPWR _07022_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17667_ net4021 svm0.tA\[5\] svm0.tA\[4\] net4011 VGND VGND VPWR VPWR _09547_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_187_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14879_ _06957_ VGND VGND VPWR VPWR _00210_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19406_ net812 net869 _11242_ VGND VGND VPWR VPWR _11243_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16618_ matmul0.matmul_stage_inst.mult2\[0\] matmul0.matmul_stage_inst.mult1\[0\]
+ VGND VGND VPWR VPWR _08659_ sky130_fd_sc_hd__xor2_1
X_17598_ _09477_ _09478_ VGND VGND VPWR VPWR _09479_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19337_ net3204 _10989_ _11133_ net3167 VGND VGND VPWR VPWR _11174_ sky130_fd_sc_hd__o211ai_1
X_16549_ _08606_ _08607_ VGND VGND VPWR VPWR _08608_ sky130_fd_sc_hd__or2b_1
XFILLER_0_156_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8380 net8386 VGND VGND VPWR VPWR net8380 sky130_fd_sc_hd__buf_1
X_19268_ _11103_ _11104_ _11096_ VGND VGND VPWR VPWR _11105_ sky130_fd_sc_hd__o21ai_1
X_18219_ net2546 _10069_ VGND VGND VPWR VPWR _10070_ sky130_fd_sc_hd__nand2_1
X_19199_ net6179 net6227 VGND VGND VPWR VPWR _11036_ sky130_fd_sc_hd__nand2_1
X_21230_ net4320 net480 _01243_ net4384 _01245_ VGND VGND VPWR VPWR _01246_ sky130_fd_sc_hd__a221o_1
Xhold201 pid_d.mult0.b\[8\] VGND VGND VPWR VPWR net9154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 svm0.tB\[10\] VGND VGND VPWR VPWR net9165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 svm0.tB\[11\] VGND VGND VPWR VPWR net9176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21161_ net5611 net5916 VGND VGND VPWR VPWR _01177_ sky130_fd_sc_hd__or2_1
Xhold234 cordic0.slte0.opA\[2\] VGND VGND VPWR VPWR net9187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 svm0.tC\[10\] VGND VGND VPWR VPWR net9198 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold256 pid_d.prev_int\[4\] VGND VGND VPWR VPWR net9209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 svm0.tA\[7\] VGND VGND VPWR VPWR net9220 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3209 _10829_ VGND VGND VPWR VPWR net3209 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20112_ _11939_ _11447_ _11890_ VGND VGND VPWR VPWR _11940_ sky130_fd_sc_hd__mux2_1
Xhold278 matmul0.a\[4\] VGND VGND VPWR VPWR net9231 sky130_fd_sc_hd__dlygate4sd3_1
X_21092_ _01106_ _01107_ _00871_ VGND VGND VPWR VPWR _01108_ sky130_fd_sc_hd__a21oi_1
Xhold289 matmul0.b\[11\] VGND VGND VPWR VPWR net9242 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2508 _11189_ VGND VGND VPWR VPWR net2508 sky130_fd_sc_hd__clkbuf_1
Xwire2519 _11053_ VGND VGND VPWR VPWR net2519 sky130_fd_sc_hd__buf_1
X_24920_ _04707_ VGND VGND VPWR VPWR _00747_ sky130_fd_sc_hd__clkbuf_1
X_20043_ _11848_ _11872_ VGND VGND VPWR VPWR _11873_ sky130_fd_sc_hd__xnor2_4
Xwire1807 net1809 VGND VGND VPWR VPWR net1807 sky130_fd_sc_hd__buf_1
Xwire1829 net1831 VGND VGND VPWR VPWR net1829 sky130_fd_sc_hd__buf_1
X_24851_ net4806 net2007 _04540_ net231 _04658_ VGND VGND VPWR VPWR _00727_ sky130_fd_sc_hd__a221o_1
X_23802_ net7503 _03666_ _03667_ VGND VGND VPWR VPWR _03668_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_0_Left_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24782_ net5214 net2390 VGND VGND VPWR VPWR _04609_ sky130_fd_sc_hd__nand2_1
X_21994_ _02000_ _02001_ _01894_ VGND VGND VPWR VPWR _02002_ sky130_fd_sc_hd__a21o_1
X_23733_ _03593_ _03598_ VGND VGND VPWR VPWR _03599_ sky130_fd_sc_hd__xnor2_1
X_20945_ _12556_ _00959_ net3825 VGND VGND VPWR VPWR _00961_ sky130_fd_sc_hd__and3_1
Xmax_length7259 net7249 VGND VGND VPWR VPWR net7259 sky130_fd_sc_hd__buf_1
Xmax_length6514 net6512 VGND VGND VPWR VPWR net6514 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6536 net6537 VGND VGND VPWR VPWR net6536 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_178_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23664_ _03411_ _03412_ _03413_ VGND VGND VPWR VPWR _03531_ sky130_fd_sc_hd__o21a_1
XFILLER_0_138_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20876_ _00891_ _00878_ _00887_ VGND VGND VPWR VPWR _00892_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25403_ clknet_leaf_72_clk _00286_ net8469 VGND VGND VPWR VPWR matmul0.a\[6\] sky130_fd_sc_hd__dfrtp_1
X_22615_ _02585_ net3770 _02586_ VGND VGND VPWR VPWR _02587_ sky130_fd_sc_hd__and3b_1
X_23595_ _03449_ _03462_ VGND VGND VPWR VPWR _03463_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25334_ clknet_leaf_82_clk _00217_ net8502 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_22546_ net9121 net2050 _02535_ VGND VGND VPWR VPWR _00545_ sky130_fd_sc_hd__a21o_1
XFILLER_0_161_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25265_ clknet_leaf_88_clk _00148_ net8435 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.b\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_22477_ net3829 _02433_ VGND VGND VPWR VPWR _02478_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5101 net5102 VGND VGND VPWR VPWR net5101 sky130_fd_sc_hd__clkbuf_1
Xwire5112 net5116 VGND VGND VPWR VPWR net5112 sky130_fd_sc_hd__buf_1
X_24216_ net2410 _04075_ net2021 VGND VGND VPWR VPWR _04077_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21428_ _01396_ _01409_ _01398_ VGND VGND VPWR VPWR _01441_ sky130_fd_sc_hd__o21ba_1
Xwire5123 net5117 VGND VGND VPWR VPWR net5123 sky130_fd_sc_hd__clkbuf_1
X_25196_ clknet_leaf_63_clk _00085_ net8665 VGND VGND VPWR VPWR matmul0.b_in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire5134 net5135 VGND VGND VPWR VPWR net5134 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5145 net5139 VGND VGND VPWR VPWR net5145 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4411 net4412 VGND VGND VPWR VPWR net4411 sky130_fd_sc_hd__clkbuf_1
X_24147_ net4788 net3052 VGND VGND VPWR VPWR _04009_ sky130_fd_sc_hd__nand2_1
Xwire4422 net4423 VGND VGND VPWR VPWR net4422 sky130_fd_sc_hd__clkbuf_1
Xwire5167 pid_q.curr_error\[12\] VGND VGND VPWR VPWR net5167 sky130_fd_sc_hd__buf_1
XFILLER_0_32_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21359_ net5844 net5476 VGND VGND VPWR VPWR _01373_ sky130_fd_sc_hd__nand2_1
Xwire5178 pid_q.curr_int\[7\] VGND VGND VPWR VPWR net5178 sky130_fd_sc_hd__clkbuf_2
Xwire4433 net4434 VGND VGND VPWR VPWR net4433 sky130_fd_sc_hd__clkbuf_1
Xwire4444 net4445 VGND VGND VPWR VPWR net4444 sky130_fd_sc_hd__clkbuf_1
Xwire3710 net3711 VGND VGND VPWR VPWR net3710 sky130_fd_sc_hd__buf_1
Xwire4455 net4456 VGND VGND VPWR VPWR net4455 sky130_fd_sc_hd__clkbuf_1
Xwire3721 net3722 VGND VGND VPWR VPWR net3721 sky130_fd_sc_hd__clkbuf_1
X_24078_ net595 net592 VGND VGND VPWR VPWR _03941_ sky130_fd_sc_hd__nand2_1
Xwire3732 net3733 VGND VGND VPWR VPWR net3732 sky130_fd_sc_hd__buf_1
Xwire3743 _03608_ VGND VGND VPWR VPWR net3743 sky130_fd_sc_hd__clkbuf_2
Xwire4488 net4489 VGND VGND VPWR VPWR net4488 sky130_fd_sc_hd__buf_1
Xwire4499 net4500 VGND VGND VPWR VPWR net4499 sky130_fd_sc_hd__buf_1
Xwire3754 net3755 VGND VGND VPWR VPWR net3754 sky130_fd_sc_hd__clkbuf_1
X_23029_ _02895_ _02896_ _02898_ VGND VGND VPWR VPWR _02899_ sky130_fd_sc_hd__a21oi_1
Xwire3765 net3766 VGND VGND VPWR VPWR net3765 sky130_fd_sc_hd__clkbuf_1
X_15920_ _07865_ _07867_ _07863_ VGND VGND VPWR VPWR _07989_ sky130_fd_sc_hd__o21a_1
Xwire3776 _01873_ VGND VGND VPWR VPWR net3776 sky130_fd_sc_hd__buf_1
XFILLER_0_127_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3798 net3799 VGND VGND VPWR VPWR net3798 sky130_fd_sc_hd__clkbuf_1
X_15851_ _07919_ _07920_ VGND VGND VPWR VPWR _07921_ sky130_fd_sc_hd__or2b_1
X_14802_ net3626 net7178 net3622 VGND VGND VPWR VPWR _06918_ sky130_fd_sc_hd__or3_1
X_15782_ _07762_ _07764_ _07851_ VGND VGND VPWR VPWR _07852_ sky130_fd_sc_hd__a21o_1
X_18570_ _10372_ _10417_ _10350_ VGND VGND VPWR VPWR _10418_ sky130_fd_sc_hd__a21o_1
XFILLER_0_157_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12994_ net7822 _04957_ _04959_ VGND VGND VPWR VPWR _05267_ sky130_fd_sc_hd__and3_1
X_17521_ net6742 _09405_ VGND VGND VPWR VPWR _09406_ sky130_fd_sc_hd__xor2_1
X_14733_ net3619 VGND VGND VPWR VPWR _06869_ sky130_fd_sc_hd__buf_1
Xmax_length8461 net8459 VGND VGND VPWR VPWR net8461 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_86_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17452_ net6743 _09341_ _09342_ net6736 VGND VGND VPWR VPWR _09347_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14664_ net7441 VGND VGND VPWR VPWR _06817_ sky130_fd_sc_hd__inv_2
Xmax_length7782 net7783 VGND VGND VPWR VPWR net7782 sky130_fd_sc_hd__clkbuf_1
X_16403_ _08447_ _08464_ VGND VGND VPWR VPWR _08465_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13615_ _05883_ _05884_ VGND VGND VPWR VPWR _05885_ sky130_fd_sc_hd__xor2_1
X_17383_ svm0.delta\[4\] _09288_ VGND VGND VPWR VPWR _09292_ sky130_fd_sc_hd__or2_1
X_14595_ net7209 net5195 VGND VGND VPWR VPWR _06769_ sky130_fd_sc_hd__xnor2_1
X_19122_ net2112 net2111 _10957_ VGND VGND VPWR VPWR _10959_ sky130_fd_sc_hd__a21o_1
X_16334_ net2654 net2218 VGND VGND VPWR VPWR _08397_ sky130_fd_sc_hd__nor2_1
X_13546_ _05745_ _05746_ VGND VGND VPWR VPWR _05817_ sky130_fd_sc_hd__nor2_1
XFILLER_0_165_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19053_ net2117 net2113 VGND VGND VPWR VPWR _10890_ sky130_fd_sc_hd__and2b_1
XFILLER_0_36_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16265_ net2651 net2659 _08328_ VGND VGND VPWR VPWR _08329_ sky130_fd_sc_hd__or3_1
X_13477_ net1574 net1572 VGND VGND VPWR VPWR _05750_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18004_ net3237 _09846_ _09854_ _09844_ net3337 VGND VGND VPWR VPWR _09855_ sky130_fd_sc_hd__o311a_1
X_15216_ _07288_ _07289_ VGND VGND VPWR VPWR _07290_ sky130_fd_sc_hd__xnor2_1
Xwire7081 net7083 VGND VGND VPWR VPWR net7081 sky130_fd_sc_hd__buf_1
XFILLER_0_51_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16196_ _08259_ _08260_ VGND VGND VPWR VPWR _08261_ sky130_fd_sc_hd__and2b_1
XFILLER_0_112_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6380 net6381 VGND VGND VPWR VPWR net6380 sky130_fd_sc_hd__clkbuf_1
Xwire6391 net6392 VGND VGND VPWR VPWR net6391 sky130_fd_sc_hd__clkbuf_1
X_15147_ net3464 _07129_ VGND VGND VPWR VPWR _07221_ sky130_fd_sc_hd__nand2_1
XFILLER_0_168_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5595 net5604 VGND VGND VPWR VPWR net5595 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout4894 net4898 VGND VGND VPWR VPWR net4894 sky130_fd_sc_hd__buf_1
Xwire5690 net5691 VGND VGND VPWR VPWR net5690 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19955_ net8997 net1202 _11786_ net1770 VGND VGND VPWR VPWR _00458_ sky130_fd_sc_hd__a22o_1
X_15078_ _07136_ VGND VGND VPWR VPWR _07152_ sky130_fd_sc_hd__clkbuf_2
X_14029_ _06291_ net1560 VGND VGND VPWR VPWR _06293_ sky130_fd_sc_hd__xor2_2
X_18906_ net302 _10729_ VGND VGND VPWR VPWR _10747_ sky130_fd_sc_hd__or2_1
X_19886_ _11717_ _11718_ net604 VGND VGND VPWR VPWR _11719_ sky130_fd_sc_hd__mux2_1
X_18837_ net3282 net3922 net6779 VGND VGND VPWR VPWR _10680_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_184_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18768_ _10561_ net764 net526 VGND VGND VPWR VPWR _10613_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17719_ pid_q.prev_int\[10\] net1455 net1788 net9202 VGND VGND VPWR VPWR _00424_
+ sky130_fd_sc_hd__a22o_1
X_18699_ net1066 _10544_ VGND VGND VPWR VPWR _10545_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20730_ _12499_ VGND VGND VPWR VPWR _12501_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20661_ net3152 net1816 _12437_ VGND VGND VPWR VPWR _12439_ sky130_fd_sc_hd__or3b_1
XFILLER_0_133_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22400_ pid_d.prev_error\[13\] net5965 _02401_ VGND VGND VPWR VPWR _02402_ sky130_fd_sc_hd__a21bo_1
X_23380_ _03248_ _03249_ VGND VGND VPWR VPWR _03250_ sky130_fd_sc_hd__xor2_1
X_20592_ net8057 net3164 _12373_ _12374_ VGND VGND VPWR VPWR _00507_ sky130_fd_sc_hd__a31o_1
XFILLER_0_34_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22331_ pid_d.curr_int\[12\] net4391 VGND VGND VPWR VPWR _02334_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25050_ _03955_ _04795_ pid_q.out\[7\] VGND VGND VPWR VPWR _04800_ sky130_fd_sc_hd__a21bo_1
X_22262_ pid_d.prev_error\[11\] net5966 VGND VGND VPWR VPWR _02266_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24001_ net5178 pid_q.prev_int\[7\] VGND VGND VPWR VPWR _03864_ sky130_fd_sc_hd__xor2_1
XFILLER_0_42_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21213_ net1732 _01010_ net1183 VGND VGND VPWR VPWR _01229_ sky130_fd_sc_hd__a21o_1
X_22193_ _02159_ _02188_ _02195_ net2062 _02197_ VGND VGND VPWR VPWR _02198_ sky130_fd_sc_hd__o221a_1
XFILLER_0_111_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21144_ net5617 net5881 VGND VGND VPWR VPWR _01160_ sky130_fd_sc_hd__nand2_1
Xwire3028 net3029 VGND VGND VPWR VPWR net3028 sky130_fd_sc_hd__buf_1
Xwire2 _08877_ VGND VGND VPWR VPWR net9247 sky130_fd_sc_hd__clkbuf_1
Xwire3039 _04348_ VGND VGND VPWR VPWR net3039 sky130_fd_sc_hd__clkbuf_1
Xwire2305 net2306 VGND VGND VPWR VPWR net2305 sky130_fd_sc_hd__buf_1
XFILLER_0_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2327 net2328 VGND VGND VPWR VPWR net2327 sky130_fd_sc_hd__buf_1
X_21075_ _01080_ _01081_ _01079_ VGND VGND VPWR VPWR _01091_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2338 net2339 VGND VGND VPWR VPWR net2338 sky130_fd_sc_hd__buf_1
Xwire2349 _04918_ VGND VGND VPWR VPWR net2349 sky130_fd_sc_hd__clkbuf_1
Xwire1604 _05037_ VGND VGND VPWR VPWR net1604 sky130_fd_sc_hd__buf_1
X_24903_ _04693_ VGND VGND VPWR VPWR _00744_ sky130_fd_sc_hd__clkbuf_1
Xwire1615 _04920_ VGND VGND VPWR VPWR net1615 sky130_fd_sc_hd__buf_1
X_20026_ net6081 _11800_ _11854_ _11855_ VGND VGND VPWR VPWR _11856_ sky130_fd_sc_hd__a31o_1
Xwire1637 _04701_ VGND VGND VPWR VPWR net1637 sky130_fd_sc_hd__buf_1
X_25883_ clknet_leaf_16_clk _00756_ net8625 VGND VGND VPWR VPWR pid_q.ki\[11\] sky130_fd_sc_hd__dfrtp_1
Xwire1648 _04507_ VGND VGND VPWR VPWR net1648 sky130_fd_sc_hd__buf_1
X_24834_ net7481 net738 net854 VGND VGND VPWR VPWR _04650_ sky130_fd_sc_hd__a21o_1
X_24765_ net7985 net4256 VGND VGND VPWR VPWR _04594_ sky130_fd_sc_hd__xnor2_1
X_21977_ _01980_ _01984_ VGND VGND VPWR VPWR _01985_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23716_ _03580_ _03581_ VGND VGND VPWR VPWR _03582_ sky130_fd_sc_hd__xnor2_1
Xmax_length6322 net6323 VGND VGND VPWR VPWR net6322 sky130_fd_sc_hd__buf_1
Xmax_length7067 net7066 VGND VGND VPWR VPWR net7067 sky130_fd_sc_hd__buf_1
XFILLER_0_68_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20928_ net5527 net5884 _00943_ VGND VGND VPWR VPWR _00944_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24696_ net4310 net3269 VGND VGND VPWR VPWR _04534_ sky130_fd_sc_hd__or2_1
Xmax_length5610 pid_d.mult0.a\[3\] VGND VGND VPWR VPWR net5610 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23647_ net4548 net5052 VGND VGND VPWR VPWR _03514_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20859_ _00862_ _00874_ VGND VGND VPWR VPWR _00875_ sky130_fd_sc_hd__xnor2_2
X_13400_ _05661_ _05667_ _05671_ _05672_ VGND VGND VPWR VPWR _05673_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14380_ net8285 net3637 VGND VGND VPWR VPWR _06588_ sky130_fd_sc_hd__and2_1
X_23578_ _03425_ _03445_ VGND VGND VPWR VPWR _03446_ sky130_fd_sc_hd__nor2_1
Xwire901 _06572_ VGND VGND VPWR VPWR net901 sky130_fd_sc_hd__buf_1
XFILLER_0_187_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire912 _05737_ VGND VGND VPWR VPWR net912 sky130_fd_sc_hd__buf_1
XFILLER_0_91_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire923 _04649_ VGND VGND VPWR VPWR net923 sky130_fd_sc_hd__clkbuf_1
X_13331_ _05590_ net844 VGND VGND VPWR VPWR _05604_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25317_ clknet_leaf_78_clk _00200_ net8439 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.f\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire934 net935 VGND VGND VPWR VPWR net934 sky130_fd_sc_hd__dlymetal6s2s_1
X_22529_ net5971 net2379 net2046 VGND VGND VPWR VPWR _02527_ sky130_fd_sc_hd__and3_1
Xwire945 _02078_ VGND VGND VPWR VPWR net945 sky130_fd_sc_hd__buf_1
Xwire956 net957 VGND VGND VPWR VPWR net956 sky130_fd_sc_hd__buf_1
XFILLER_0_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire967 net968 VGND VGND VPWR VPWR net967 sky130_fd_sc_hd__buf_1
XFILLER_0_17_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16050_ _08115_ _08116_ VGND VGND VPWR VPWR _08117_ sky130_fd_sc_hd__xnor2_1
X_13262_ _05533_ _05534_ VGND VGND VPWR VPWR _05535_ sky130_fd_sc_hd__xnor2_1
X_25248_ clknet_leaf_87_clk _00131_ net8436 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.a\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire978 _08335_ VGND VGND VPWR VPWR net978 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire989 _07727_ VGND VGND VPWR VPWR net989 sky130_fd_sc_hd__clkbuf_1
X_15001_ net1898 _07074_ VGND VGND VPWR VPWR _07075_ sky130_fd_sc_hd__xnor2_2
X_13193_ _05464_ _05465_ VGND VGND VPWR VPWR _05466_ sky130_fd_sc_hd__nand2_1
X_25179_ clknet_leaf_95_clk _00068_ net8448 VGND VGND VPWR VPWR matmul0.a_in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire4230 net4231 VGND VGND VPWR VPWR net4230 sky130_fd_sc_hd__clkbuf_1
Xwire4241 net4242 VGND VGND VPWR VPWR net4241 sky130_fd_sc_hd__buf_1
Xwire4252 net4253 VGND VGND VPWR VPWR net4252 sky130_fd_sc_hd__clkbuf_1
Xwire4263 net4264 VGND VGND VPWR VPWR net4263 sky130_fd_sc_hd__clkbuf_1
Xwire4274 net4276 VGND VGND VPWR VPWR net4274 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3540 _07049_ VGND VGND VPWR VPWR net3540 sky130_fd_sc_hd__clkbuf_1
Xwire4285 net4286 VGND VGND VPWR VPWR net4285 sky130_fd_sc_hd__buf_1
X_19740_ net3157 _11522_ _11164_ VGND VGND VPWR VPWR _11575_ sky130_fd_sc_hd__a21o_1
Xwire3551 net3552 VGND VGND VPWR VPWR net3551 sky130_fd_sc_hd__buf_1
Xwire4296 _04875_ VGND VGND VPWR VPWR net4296 sky130_fd_sc_hd__clkbuf_1
X_16952_ net4246 net2197 VGND VGND VPWR VPWR _08915_ sky130_fd_sc_hd__nor2_1
Xwire3562 net3563 VGND VGND VPWR VPWR net3562 sky130_fd_sc_hd__buf_1
XFILLER_0_47_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3573 net3574 VGND VGND VPWR VPWR net3573 sky130_fd_sc_hd__buf_1
X_15903_ net2734 net3425 net3427 net3460 VGND VGND VPWR VPWR _07972_ sky130_fd_sc_hd__a211o_1
Xwire2850 _06988_ VGND VGND VPWR VPWR net2850 sky130_fd_sc_hd__buf_1
Xwire3595 _06984_ VGND VGND VPWR VPWR net3595 sky130_fd_sc_hd__buf_1
X_19671_ net6198 net6238 net3154 net6156 VGND VGND VPWR VPWR _11507_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2861 _06838_ VGND VGND VPWR VPWR net2861 sky130_fd_sc_hd__dlymetal6s2s_1
X_16883_ _08827_ _08846_ net6525 VGND VGND VPWR VPWR _08847_ sky130_fd_sc_hd__mux2_1
Xwire2872 _06814_ VGND VGND VPWR VPWR net2872 sky130_fd_sc_hd__buf_1
XFILLER_0_194_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2883 net2884 VGND VGND VPWR VPWR net2883 sky130_fd_sc_hd__buf_1
X_18622_ net6919 _10223_ _10431_ VGND VGND VPWR VPWR _10469_ sky130_fd_sc_hd__nor3_1
XFILLER_0_189_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15834_ _07895_ net1263 VGND VGND VPWR VPWR _07904_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18553_ _10397_ _10401_ VGND VGND VPWR VPWR _10402_ sky130_fd_sc_hd__xor2_1
XFILLER_0_188_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12977_ net7759 net1986 net2364 VGND VGND VPWR VPWR _05250_ sky130_fd_sc_hd__and3_1
X_15765_ net3449 net3438 VGND VGND VPWR VPWR _07835_ sky130_fd_sc_hd__nor2_1
X_17504_ _09258_ net2571 _09389_ _09391_ VGND VGND VPWR VPWR _00401_ sky130_fd_sc_hd__a31o_1
X_14716_ matmul0.sin\[12\] _06856_ VGND VGND VPWR VPWR _06857_ sky130_fd_sc_hd__xnor2_1
X_15696_ net2676 _07672_ _07671_ VGND VGND VPWR VPWR _07767_ sky130_fd_sc_hd__a21o_1
X_18484_ _10332_ _10333_ VGND VGND VPWR VPWR _10334_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17435_ net7376 net3274 net6656 VGND VGND VPWR VPWR _09333_ sky130_fd_sc_hd__o21a_1
X_14647_ net7440 net7178 net2874 VGND VGND VPWR VPWR _06808_ sky130_fd_sc_hd__and3_1
XFILLER_0_184_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_72_Left_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17366_ net3276 VGND VGND VPWR VPWR _09278_ sky130_fd_sc_hd__buf_1
X_14578_ net7234 net5207 VGND VGND VPWR VPWR _06754_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_166_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19105_ net6243 _10941_ net3889 VGND VGND VPWR VPWR _10942_ sky130_fd_sc_hd__a21o_1
X_13529_ _05704_ net1128 net1129 VGND VGND VPWR VPWR _05800_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16317_ _08318_ _08351_ _08379_ VGND VGND VPWR VPWR _08380_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17297_ net7765 net7742 net7719 net1795 VGND VGND VPWR VPWR _09211_ sky130_fd_sc_hd__or4_1
XFILLER_0_166_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19036_ net6204 net6154 _10870_ VGND VGND VPWR VPWR _10873_ sky130_fd_sc_hd__and3_1
X_16248_ net3587 net2215 VGND VGND VPWR VPWR _08312_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5381 net5387 VGND VGND VPWR VPWR net5381 sky130_fd_sc_hd__buf_1
X_16179_ net672 _08222_ _08212_ VGND VGND VPWR VPWR _08244_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout4680 pid_q.mult0.a\[5\] VGND VGND VPWR VPWR net4680 sky130_fd_sc_hd__buf_1
XFILLER_0_103_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_81_Left_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19938_ net6013 _11448_ _11769_ VGND VGND VPWR VPWR _11770_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19869_ net6009 net6033 net2500 _11648_ VGND VGND VPWR VPWR _11702_ sky130_fd_sc_hd__or4_1
X_21900_ _01908_ _01812_ pid_d.prev_error\[6\] VGND VGND VPWR VPWR _01909_ sky130_fd_sc_hd__o21ba_1
X_22880_ net8898 _02775_ VGND VGND VPWR VPWR _02776_ sky130_fd_sc_hd__and2_1
XFILLER_0_179_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21831_ _01838_ _01839_ VGND VGND VPWR VPWR _01840_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_144_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24550_ _04357_ _04361_ _04362_ VGND VGND VPWR VPWR _04406_ sky130_fd_sc_hd__o21a_1
X_21762_ _01673_ _01675_ VGND VGND VPWR VPWR _01772_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_90_Left_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23501_ net1028 _03369_ VGND VGND VPWR VPWR _03370_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20713_ net2186 _12485_ _09023_ VGND VGND VPWR VPWR _12486_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24481_ net1650 _04306_ VGND VGND VPWR VPWR _04338_ sky130_fd_sc_hd__xor2_1
XFILLER_0_59_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21693_ net1720 _01702_ VGND VGND VPWR VPWR _01704_ sky130_fd_sc_hd__nand2_1
Xwire8507 net8508 VGND VGND VPWR VPWR net8507 sky130_fd_sc_hd__clkbuf_2
Xmax_length4205 net4206 VGND VGND VPWR VPWR net4205 sky130_fd_sc_hd__buf_1
X_23432_ _03200_ _03229_ _03183_ VGND VGND VPWR VPWR _03302_ sky130_fd_sc_hd__a21bo_1
Xwire7806 net7807 VGND VGND VPWR VPWR net7806 sky130_fd_sc_hd__buf_1
Xmax_length4238 _06503_ VGND VGND VPWR VPWR net4238 sky130_fd_sc_hd__clkbuf_1
X_20644_ _12421_ _12422_ VGND VGND VPWR VPWR _12423_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7817 net7818 VGND VGND VPWR VPWR net7817 sky130_fd_sc_hd__clkbuf_1
Xwire208 _08496_ VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__buf_1
Xwire219 _06321_ VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__buf_1
Xwire7828 net7829 VGND VGND VPWR VPWR net7828 sky130_fd_sc_hd__buf_1
X_23363_ _02932_ _02963_ net1032 VGND VGND VPWR VPWR _03233_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20575_ _12357_ _12358_ VGND VGND VPWR VPWR _12359_ sky130_fd_sc_hd__and2b_1
XFILLER_0_117_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25102_ _04836_ _04839_ _04844_ VGND VGND VPWR VPWR _04845_ sky130_fd_sc_hd__o21a_1
X_22314_ _02281_ _02317_ VGND VGND VPWR VPWR _02318_ sky130_fd_sc_hd__xnor2_2
X_23294_ net1031 _03162_ VGND VGND VPWR VPWR _03164_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25033_ _04783_ net1628 net2147 VGND VGND VPWR VPWR _04786_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22245_ _02249_ VGND VGND VPWR VPWR _02250_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22176_ pid_d.curr_int\[10\] net3843 net2487 _02181_ VGND VGND VPWR VPWR _00529_
+ sky130_fd_sc_hd__a22o_1
Xwire2102 _11468_ VGND VGND VPWR VPWR net2102 sky130_fd_sc_hd__clkbuf_1
X_21127_ _01139_ _01133_ VGND VGND VPWR VPWR _01143_ sky130_fd_sc_hd__and2b_1
Xwire2113 net2114 VGND VGND VPWR VPWR net2113 sky130_fd_sc_hd__clkbuf_1
Xwire2124 _10771_ VGND VGND VPWR VPWR net2124 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2135 net2136 VGND VGND VPWR VPWR net2135 sky130_fd_sc_hd__buf_1
Xwire1401 net1402 VGND VGND VPWR VPWR net1401 sky130_fd_sc_hd__clkbuf_1
Xwire1412 net1413 VGND VGND VPWR VPWR net1412 sky130_fd_sc_hd__buf_1
X_25935_ clknet_leaf_24_clk _00808_ net8589 VGND VGND VPWR VPWR pid_d.prev_int\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21058_ net3121 _01072_ _01073_ VGND VGND VPWR VPWR _01074_ sky130_fd_sc_hd__o21ba_1
Xwire1423 net1424 VGND VGND VPWR VPWR net1423 sky130_fd_sc_hd__clkbuf_1
Xwire2168 _09096_ VGND VGND VPWR VPWR net2168 sky130_fd_sc_hd__buf_1
Xwire2179 net2180 VGND VGND VPWR VPWR net2179 sky130_fd_sc_hd__buf_1
Xwire1434 _10471_ VGND VGND VPWR VPWR net1434 sky130_fd_sc_hd__clkbuf_1
X_12900_ _05171_ _05172_ VGND VGND VPWR VPWR _05173_ sky130_fd_sc_hd__xor2_1
Xwire1445 net1446 VGND VGND VPWR VPWR net1445 sky130_fd_sc_hd__buf_1
Xwire1456 net1457 VGND VGND VPWR VPWR net1456 sky130_fd_sc_hd__buf_1
X_20009_ _11838_ VGND VGND VPWR VPWR _11839_ sky130_fd_sc_hd__inv_2
X_13880_ net532 _06080_ VGND VGND VPWR VPWR _06147_ sky130_fd_sc_hd__or2_1
X_25866_ clknet_leaf_16_clk _00739_ net8625 VGND VGND VPWR VPWR pid_q.mult0.a\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1467 net1468 VGND VGND VPWR VPWR net1467 sky130_fd_sc_hd__clkbuf_1
Xwire1478 _09036_ VGND VGND VPWR VPWR net1478 sky130_fd_sc_hd__buf_1
Xwire1489 net1498 VGND VGND VPWR VPWR net1489 sky130_fd_sc_hd__clkbuf_1
X_24817_ net7949 _04639_ VGND VGND VPWR VPWR _04640_ sky130_fd_sc_hd__xnor2_1
X_12831_ net7875 _04956_ net2975 VGND VGND VPWR VPWR _05104_ sky130_fd_sc_hd__and3_1
X_25797_ clknet_leaf_32_clk _00670_ net8682 VGND VGND VPWR VPWR pid_q.curr_int\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_185_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15550_ _07617_ _07622_ VGND VGND VPWR VPWR _07623_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_55_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24748_ _04577_ net8002 _04571_ _04570_ VGND VGND VPWR VPWR _04579_ sky130_fd_sc_hd__a211o_1
X_12762_ net7337 _04892_ net3695 VGND VGND VPWR VPWR _05035_ sky130_fd_sc_hd__nand3_1
XFILLER_0_97_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14501_ net9058 net832 net1292 _06683_ VGND VGND VPWR VPWR _00106_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15481_ _07475_ _07554_ VGND VGND VPWR VPWR _07555_ sky130_fd_sc_hd__xor2_1
XFILLER_0_84_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12693_ net7905 net1963 VGND VGND VPWR VPWR _04966_ sky130_fd_sc_hd__nand2_1
X_24679_ pid_q.curr_error\[11\] net3021 net1646 VGND VGND VPWR VPWR _04522_ sky130_fd_sc_hd__and3_1
X_14432_ net8194 net3632 VGND VGND VPWR VPWR _06628_ sky130_fd_sc_hd__and2_1
X_17220_ net6788 net1821 _09167_ VGND VGND VPWR VPWR _09169_ sky130_fd_sc_hd__or3_1
XFILLER_0_166_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17151_ net6932 _09075_ _09103_ VGND VGND VPWR VPWR _09105_ sky130_fd_sc_hd__or3_1
X_14363_ net4233 VGND VGND VPWR VPWR _06575_ sky130_fd_sc_hd__buf_1
Xwire720 net721 VGND VGND VPWR VPWR net720 sky130_fd_sc_hd__buf_1
XFILLER_0_25_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire731 _05605_ VGND VGND VPWR VPWR net731 sky130_fd_sc_hd__buf_1
Xinput16 angle_in[9] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_1
Xinput27 currA_in[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire742 _03952_ VGND VGND VPWR VPWR net742 sky130_fd_sc_hd__clkbuf_1
Xmax_length4794 net4787 VGND VGND VPWR VPWR net4794 sky130_fd_sc_hd__buf_1
X_16102_ _08105_ _08165_ _08167_ VGND VGND VPWR VPWR _08168_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_181_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire753 net754 VGND VGND VPWR VPWR net753 sky130_fd_sc_hd__clkbuf_1
X_13314_ _05585_ _05586_ VGND VGND VPWR VPWR _05587_ sky130_fd_sc_hd__xnor2_1
Xinput38 currB_in[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_1
Xinput49 currT_in[0] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
X_17082_ _08977_ _09018_ _09014_ VGND VGND VPWR VPWR _09040_ sky130_fd_sc_hd__o21bai_1
Xwire764 _10563_ VGND VGND VPWR VPWR net764 sky130_fd_sc_hd__buf_2
X_14294_ net68 net2901 net2264 net7670 VGND VGND VPWR VPWR _00063_ sky130_fd_sc_hd__a22o_1
Xwire775 _08169_ VGND VGND VPWR VPWR net775 sky130_fd_sc_hd__clkbuf_1
Xwire786 net787 VGND VGND VPWR VPWR net786 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire797 net798 VGND VGND VPWR VPWR net797 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16033_ net2239 _08056_ VGND VGND VPWR VPWR _08100_ sky130_fd_sc_hd__nand2_1
X_13245_ net7845 net1947 VGND VGND VPWR VPWR _05518_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13176_ _05432_ _05433_ net1000 net999 VGND VGND VPWR VPWR _05449_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_23_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4060 _08832_ VGND VGND VPWR VPWR net4060 sky130_fd_sc_hd__buf_1
XFILLER_0_196_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4071 net4072 VGND VGND VPWR VPWR net4071 sky130_fd_sc_hd__buf_1
XFILLER_0_20_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4082 _07515_ VGND VGND VPWR VPWR net4082 sky130_fd_sc_hd__clkbuf_1
X_17984_ _09825_ net1779 VGND VGND VPWR VPWR _09835_ sky130_fd_sc_hd__or2_1
Xwire4093 _07369_ VGND VGND VPWR VPWR net4093 sky130_fd_sc_hd__clkbuf_1
Xwire3370 net3371 VGND VGND VPWR VPWR net3370 sky130_fd_sc_hd__clkbuf_2
X_19723_ _11557_ _11543_ net3857 VGND VGND VPWR VPWR _11558_ sky130_fd_sc_hd__mux2_1
Xwire3381 net3382 VGND VGND VPWR VPWR net3381 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_165_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16935_ _08889_ _08894_ _08895_ _08898_ net3360 VGND VGND VPWR VPWR _08899_ sky130_fd_sc_hd__o2111a_1
Xwire3392 net3393 VGND VGND VPWR VPWR net3392 sky130_fd_sc_hd__buf_1
Xwire2680 _07560_ VGND VGND VPWR VPWR net2680 sky130_fd_sc_hd__buf_1
X_19654_ net6002 net6022 VGND VGND VPWR VPWR _11490_ sky130_fd_sc_hd__nand2_2
Xwire2691 net2692 VGND VGND VPWR VPWR net2691 sky130_fd_sc_hd__buf_1
X_16866_ _08829_ net4061 _08825_ VGND VGND VPWR VPWR _08831_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18605_ net1196 _10452_ VGND VGND VPWR VPWR _10453_ sky130_fd_sc_hd__and2_1
Xwire1990 _04859_ VGND VGND VPWR VPWR net1990 sky130_fd_sc_hd__buf_1
X_15817_ _07885_ _07886_ VGND VGND VPWR VPWR _07887_ sky130_fd_sc_hd__or2_1
X_19585_ _11358_ _11420_ _11421_ VGND VGND VPWR VPWR _11422_ sky130_fd_sc_hd__a21o_1
XFILLER_0_177_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16797_ _08788_ VGND VGND VPWR VPWR _00297_ sky130_fd_sc_hd__clkbuf_1
X_18536_ _10322_ net1205 _10308_ VGND VGND VPWR VPWR _10385_ sky130_fd_sc_hd__o21ba_1
X_15748_ _07800_ _07818_ VGND VGND VPWR VPWR _07819_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_90_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18467_ _10309_ _10312_ _10316_ VGND VGND VPWR VPWR _10317_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15679_ net2671 net2668 net3395 net2235 VGND VGND VPWR VPWR _07750_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17418_ svm0.delta\[11\] _09316_ VGND VGND VPWR VPWR _09320_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18398_ _10217_ _10248_ VGND VGND VPWR VPWR _10249_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_99_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17349_ net3278 _09261_ _09262_ VGND VGND VPWR VPWR _09263_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_114_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20360_ _12156_ _12160_ VGND VGND VPWR VPWR _12161_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_141_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19019_ net6265 net6298 net6317 VGND VGND VPWR VPWR _10856_ sky130_fd_sc_hd__and3b_1
X_20291_ net1482 _12096_ net2604 VGND VGND VPWR VPWR _12097_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22030_ _01932_ _01937_ _01927_ VGND VGND VPWR VPWR _02037_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_12_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23981_ _03843_ _03844_ VGND VGND VPWR VPWR _03845_ sky130_fd_sc_hd__nor2_1
X_25720_ clknet_leaf_11_clk _00593_ net8603 VGND VGND VPWR VPWR pid_d.mult0.a\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_22932_ _02813_ _02820_ _02821_ VGND VGND VPWR VPWR _02822_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_119_Left_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25651_ clknet_leaf_1_clk _00524_ net8404 VGND VGND VPWR VPWR pid_d.curr_int\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_22863_ net5981 _02747_ _02759_ net5980 VGND VGND VPWR VPWR _02760_ sky130_fd_sc_hd__a211o_1
XFILLER_0_35_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24602_ net5170 pid_q.prev_int\[14\] VGND VGND VPWR VPWR _04457_ sky130_fd_sc_hd__or2_1
X_21814_ _01821_ _01822_ VGND VGND VPWR VPWR _01823_ sky130_fd_sc_hd__xnor2_1
X_25582_ clknet_leaf_86_clk _00455_ net8532 VGND VGND VPWR VPWR cordic0.cos\[2\] sky130_fd_sc_hd__dfrtp_1
X_22794_ pid_d.kp\[9\] net3070 net1687 VGND VGND VPWR VPWR _02705_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24533_ _04329_ _04389_ net9066 _02867_ VGND VGND VPWR VPWR _00678_ sky130_fd_sc_hd__a2bb2o_1
X_21745_ _01661_ _01663_ _01754_ VGND VGND VPWR VPWR _01755_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_176_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8304 net19 VGND VGND VPWR VPWR net8304 sky130_fd_sc_hd__clkbuf_1
Xwire8315 net8316 VGND VGND VPWR VPWR net8315 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_171_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8326 net8327 VGND VGND VPWR VPWR net8326 sky130_fd_sc_hd__clkbuf_1
X_24464_ pid_q.prev_error\[12\] net5167 VGND VGND VPWR VPWR _04322_ sky130_fd_sc_hd__or2_1
X_21676_ _01658_ _01686_ VGND VGND VPWR VPWR _01687_ sky130_fd_sc_hd__xnor2_1
Xwire8337 net8334 VGND VGND VPWR VPWR net8337 sky130_fd_sc_hd__buf_1
Xmax_length4035 _09196_ VGND VGND VPWR VPWR net4035 sky130_fd_sc_hd__buf_1
XFILLER_0_175_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7603 net7604 VGND VGND VPWR VPWR net7603 sky130_fd_sc_hd__buf_1
Xfanout6807 net6821 VGND VGND VPWR VPWR net6807 sky130_fd_sc_hd__dlymetal6s2s_1
X_23415_ net4637 net4989 VGND VGND VPWR VPWR _03285_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7636 net7637 VGND VGND VPWR VPWR net7636 sky130_fd_sc_hd__clkbuf_1
X_20627_ net3848 net3847 net2593 VGND VGND VPWR VPWR _12407_ sky130_fd_sc_hd__mux2_1
Xmax_length4068 net4069 VGND VGND VPWR VPWR net4068 sky130_fd_sc_hd__buf_1
X_24395_ pid_q.prev_error\[11\] pid_q.curr_error\[11\] VGND VGND VPWR VPWR _04254_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7647 net7646 VGND VGND VPWR VPWR net7647 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire6902 net6903 VGND VGND VPWR VPWR net6902 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7658 net7659 VGND VGND VPWR VPWR net7658 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_129_Right_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length3345 _08924_ VGND VGND VPWR VPWR net3345 sky130_fd_sc_hd__clkbuf_2
Xwire6913 net6905 VGND VGND VPWR VPWR net6913 sky130_fd_sc_hd__clkbuf_1
Xwire7669 net7665 VGND VGND VPWR VPWR net7669 sky130_fd_sc_hd__buf_1
XFILLER_0_116_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6924 net6926 VGND VGND VPWR VPWR net6924 sky130_fd_sc_hd__buf_1
X_23346_ _02939_ _02944_ _03215_ VGND VGND VPWR VPWR _03216_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_128_Left_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20558_ net1480 _12342_ VGND VGND VPWR VPWR _12343_ sky130_fd_sc_hd__nand2_1
Xwire6946 net6951 VGND VGND VPWR VPWR net6946 sky130_fd_sc_hd__buf_1
XFILLER_0_105_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length2644 _07838_ VGND VGND VPWR VPWR net2644 sky130_fd_sc_hd__buf_1
Xwire6968 net6961 VGND VGND VPWR VPWR net6968 sky130_fd_sc_hd__buf_1
XFILLER_0_46_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire6979 net6980 VGND VGND VPWR VPWR net6979 sky130_fd_sc_hd__dlymetal6s2s_1
X_23277_ _03114_ _03128_ _03146_ VGND VGND VPWR VPWR _03147_ sky130_fd_sc_hd__o21a_1
XFILLER_0_21_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20489_ net7129 net7113 net7088 net7056 net6507 net6489 VGND VGND VPWR VPWR _12277_
+ sky130_fd_sc_hd__mux4_1
X_25016_ _04768_ _04769_ VGND VGND VPWR VPWR _04771_ sky130_fd_sc_hd__or2_1
X_13030_ net920 _05302_ VGND VGND VPWR VPWR _05303_ sky130_fd_sc_hd__xnor2_2
X_22228_ _02221_ _02232_ VGND VGND VPWR VPWR _02233_ sky130_fd_sc_hd__xnor2_2
X_22159_ _02159_ _02164_ VGND VGND VPWR VPWR _02165_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14981_ net4198 net4197 VGND VGND VPWR VPWR _07055_ sky130_fd_sc_hd__nor2_1
XFILLER_0_195_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1220 _09250_ VGND VGND VPWR VPWR net1220 sky130_fd_sc_hd__clkbuf_1
Xwire1231 net1232 VGND VGND VPWR VPWR net1231 sky130_fd_sc_hd__buf_1
Xwire1242 _08615_ VGND VGND VPWR VPWR net1242 sky130_fd_sc_hd__buf_1
X_16720_ matmul0.matmul_stage_inst.mult2\[15\] matmul0.matmul_stage_inst.mult1\[15\]
+ VGND VGND VPWR VPWR _08746_ sky130_fd_sc_hd__xor2_1
XFILLER_0_191_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13932_ _06189_ _06197_ VGND VGND VPWR VPWR _06198_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_137_Left_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25918_ clknet_leaf_28_clk _00791_ net8651 VGND VGND VPWR VPWR pid_q.out\[14\] sky130_fd_sc_hd__dfrtp_1
Xwire1253 _08184_ VGND VGND VPWR VPWR net1253 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_135_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1264 _07845_ VGND VGND VPWR VPWR net1264 sky130_fd_sc_hd__buf_1
Xwire1275 _07324_ VGND VGND VPWR VPWR net1275 sky130_fd_sc_hd__clkbuf_2
Xwire1286 _07070_ VGND VGND VPWR VPWR net1286 sky130_fd_sc_hd__dlymetal6s2s_1
X_13863_ net3676 _06028_ VGND VGND VPWR VPWR _06130_ sky130_fd_sc_hd__nor2_1
X_16651_ _08686_ _08682_ matmul0.matmul_stage_inst.mult2\[4\] VGND VGND VPWR VPWR
+ _08687_ sky130_fd_sc_hd__o21ba_1
X_25849_ clknet_leaf_20_clk _00722_ net8616 VGND VGND VPWR VPWR pid_q.mult0.b\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12814_ _04955_ net1343 _05085_ _05086_ VGND VGND VPWR VPWR _05087_ sky130_fd_sc_hd__o211ai_1
X_15602_ net2676 _07673_ VGND VGND VPWR VPWR _07674_ sky130_fd_sc_hd__xnor2_1
X_19370_ _11206_ VGND VGND VPWR VPWR _11207_ sky130_fd_sc_hd__dlymetal6s2s_1
X_13794_ _06060_ _06061_ VGND VGND VPWR VPWR _06062_ sky130_fd_sc_hd__xor2_1
XFILLER_0_9_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16582_ _08638_ VGND VGND VPWR VPWR _00232_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_186_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18321_ _10169_ _10171_ VGND VGND VPWR VPWR _10172_ sky130_fd_sc_hd__xor2_2
X_12745_ _05008_ _05010_ _05017_ VGND VGND VPWR VPWR _05018_ sky130_fd_sc_hd__a21boi_1
X_15533_ net4207 net4201 net4083 net4081 VGND VGND VPWR VPWR _07606_ sky130_fd_sc_hd__o22a_1
XFILLER_0_155_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8743 net8747 VGND VGND VPWR VPWR net8743 sky130_fd_sc_hd__buf_1
X_15464_ net1861 net1860 VGND VGND VPWR VPWR _07538_ sky130_fd_sc_hd__xor2_1
X_18252_ net6920 net6893 VGND VGND VPWR VPWR _10103_ sky130_fd_sc_hd__nor2b_1
X_12676_ net7844 net2356 net1978 VGND VGND VPWR VPWR _04949_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14415_ _06615_ VGND VGND VPWR VPWR _00088_ sky130_fd_sc_hd__clkbuf_1
X_17203_ _09146_ _09152_ VGND VGND VPWR VPWR _09153_ sky130_fd_sc_hd__xor2_1
Xwire8860 net8861 VGND VGND VPWR VPWR net8860 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_146_Left_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15395_ _07339_ net725 _07467_ _07468_ VGND VGND VPWR VPWR _07469_ sky130_fd_sc_hd__and4_1
XFILLER_0_37_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18183_ net7063 net3254 VGND VGND VPWR VPWR _10034_ sky130_fd_sc_hd__nand2_1
XFILLER_0_182_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8882 net8883 VGND VGND VPWR VPWR net8882 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8893 net8894 VGND VGND VPWR VPWR net8893 sky130_fd_sc_hd__buf_1
XFILLER_0_181_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire550 _02385_ VGND VGND VPWR VPWR net550 sky130_fd_sc_hd__clkbuf_1
X_17134_ _09086_ _09088_ VGND VGND VPWR VPWR _09089_ sky130_fd_sc_hd__xnor2_1
X_14346_ _06561_ matmul0.a_in\[6\] net904 VGND VGND VPWR VPWR _06562_ sky130_fd_sc_hd__mux2_1
Xwire561 net562 VGND VGND VPWR VPWR net561 sky130_fd_sc_hd__buf_1
XFILLER_0_40_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire572 net573 VGND VGND VPWR VPWR net572 sky130_fd_sc_hd__buf_1
Xwire583 net584 VGND VGND VPWR VPWR net583 sky130_fd_sc_hd__buf_1
XFILLER_0_100_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire594 _03940_ VGND VGND VPWR VPWR net594 sky130_fd_sc_hd__clkbuf_1
X_17065_ net2179 _09022_ net3320 VGND VGND VPWR VPWR _09024_ sky130_fd_sc_hd__a21o_1
X_14277_ net53 net2914 _06517_ net9042 VGND VGND VPWR VPWR _00048_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16016_ _08007_ VGND VGND VPWR VPWR _08084_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13228_ _05491_ _05500_ VGND VGND VPWR VPWR _05501_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_176_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13159_ _05372_ net1138 VGND VGND VPWR VPWR _05432_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_155_Left_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17967_ net6924 net6884 _09157_ VGND VGND VPWR VPWR _09818_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19706_ _11532_ _11541_ VGND VGND VPWR VPWR _11542_ sky130_fd_sc_hd__xnor2_2
X_16918_ _08880_ _08881_ cordic0.slte0.opA\[17\] _08855_ VGND VGND VPWR VPWR _08882_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_192_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17898_ net7132 net3263 _09748_ net7091 _09650_ VGND VGND VPWR VPWR _09749_ sky130_fd_sc_hd__o221a_1
XFILLER_0_189_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19637_ net6012 _11348_ _11411_ VGND VGND VPWR VPWR _11474_ sky130_fd_sc_hd__and3_1
X_16849_ _08815_ VGND VGND VPWR VPWR _00322_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19568_ net1418 _11404_ VGND VGND VPWR VPWR _11405_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_75_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18519_ net6872 net3932 _10367_ _10174_ VGND VGND VPWR VPWR _10368_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_186_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19499_ net6116 net6128 VGND VGND VPWR VPWR _11336_ sky130_fd_sc_hd__or2_1
XFILLER_0_186_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21530_ pid_d.prev_int\[3\] _01438_ _01541_ VGND VGND VPWR VPWR _01542_ sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_164_Left_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21461_ _01360_ _01362_ _01473_ VGND VGND VPWR VPWR _01474_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_141_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6209 net6210 VGND VGND VPWR VPWR net6209 sky130_fd_sc_hd__buf_2
X_23200_ _03062_ VGND VGND VPWR VPWR _03070_ sky130_fd_sc_hd__inv_2
X_20412_ cordic0.slte0.opA\[9\] _12198_ net811 VGND VGND VPWR VPWR _12209_ sky130_fd_sc_hd__a21o_1
X_24180_ pid_q.curr_int\[9\] pid_q.prev_int\[9\] VGND VGND VPWR VPWR _04041_ sky130_fd_sc_hd__xor2_1
XFILLER_0_43_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21392_ net5444 net3812 net3789 _00821_ VGND VGND VPWR VPWR _01406_ sky130_fd_sc_hd__or4_1
Xwire5508 net5509 VGND VGND VPWR VPWR net5508 sky130_fd_sc_hd__clkbuf_1
Xwire5519 net5520 VGND VGND VPWR VPWR net5519 sky130_fd_sc_hd__clkbuf_1
X_23131_ _02993_ net2431 _03000_ VGND VGND VPWR VPWR _03001_ sky130_fd_sc_hd__o21ba_1
Xmax_length1217 net1218 VGND VGND VPWR VPWR net1217 sky130_fd_sc_hd__buf_1
X_20343_ net3668 _12133_ VGND VGND VPWR VPWR _12145_ sky130_fd_sc_hd__nor2_2
XFILLER_0_4_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4807 net4808 VGND VGND VPWR VPWR net4807 sky130_fd_sc_hd__buf_1
XFILLER_0_113_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4818 net4814 VGND VGND VPWR VPWR net4818 sky130_fd_sc_hd__clkbuf_1
X_23062_ net2026 net1678 VGND VGND VPWR VPWR _02932_ sky130_fd_sc_hd__xnor2_2
X_20274_ _12082_ VGND VGND VPWR VPWR _00481_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22013_ net5976 pid_d.prev_int\[9\] VGND VGND VPWR VPWR _02020_ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_173_Left_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23964_ _03803_ _03827_ VGND VGND VPWR VPWR _03828_ sky130_fd_sc_hd__xnor2_1
Xmax_length8813 net8808 VGND VGND VPWR VPWR net8813 sky130_fd_sc_hd__clkbuf_1
X_22915_ net5340 _02806_ net3064 VGND VGND VPWR VPWR _02807_ sky130_fd_sc_hd__mux2_1
X_25703_ clknet_leaf_2_clk _00576_ net8572 VGND VGND VPWR VPWR pid_d.mult0.b\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23895_ _03758_ _03759_ VGND VGND VPWR VPWR _03760_ sky130_fd_sc_hd__nor2_1
XFILLER_0_190_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25634_ clknet_leaf_104_clk _00507_ net8361 VGND VGND VPWR VPWR cordic0.vec\[0\]\[6\]
+ sky130_fd_sc_hd__dfstp_1
X_22846_ pid_d.out\[3\] VGND VGND VPWR VPWR _02745_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25565_ clknet_leaf_100_clk _00438_ net8390 VGND VGND VPWR VPWR cordic0.out_valid
+ sky130_fd_sc_hd__dfrtp_1
X_22777_ _02696_ VGND VGND VPWR VPWR _00615_ sky130_fd_sc_hd__clkbuf_1
Xwire8101 net89 VGND VGND VPWR VPWR net8101 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24516_ _04372_ VGND VGND VPWR VPWR _04373_ sky130_fd_sc_hd__inv_2
Xwire8112 net8113 VGND VGND VPWR VPWR net8112 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21728_ _01736_ _01646_ _01737_ VGND VGND VPWR VPWR _01738_ sky130_fd_sc_hd__a21o_1
X_25496_ clknet_leaf_42_clk _00376_ net8771 VGND VGND VPWR VPWR svm0.delta\[1\] sky130_fd_sc_hd__dfrtp_1
Xwire8123 net8124 VGND VGND VPWR VPWR net8123 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8134 net8135 VGND VGND VPWR VPWR net8134 sky130_fd_sc_hd__clkbuf_1
Xwire8145 net44 VGND VGND VPWR VPWR net8145 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24447_ _04298_ _04304_ VGND VGND VPWR VPWR _04305_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7411 net7412 VGND VGND VPWR VPWR net7411 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8156 net42 VGND VGND VPWR VPWR net8156 sky130_fd_sc_hd__clkbuf_1
X_21659_ _01666_ _01669_ VGND VGND VPWR VPWR _01670_ sky130_fd_sc_hd__xnor2_2
Xwire8167 net40 VGND VGND VPWR VPWR net8167 sky130_fd_sc_hd__clkbuf_1
Xfanout6626 net6633 VGND VGND VPWR VPWR net6626 sky130_fd_sc_hd__clkbuf_1
Xwire8178 net8179 VGND VGND VPWR VPWR net8178 sky130_fd_sc_hd__clkbuf_1
Xwire7433 matmul0.matmul_stage_inst.b\[2\] VGND VGND VPWR VPWR net7433 sky130_fd_sc_hd__buf_1
X_14200_ _06456_ _06458_ VGND VGND VPWR VPWR _06460_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5903 net5916 VGND VGND VPWR VPWR net5903 sky130_fd_sc_hd__clkbuf_1
Xwire7444 net7447 VGND VGND VPWR VPWR net7444 sky130_fd_sc_hd__clkbuf_1
Xwire8189 net36 VGND VGND VPWR VPWR net8189 sky130_fd_sc_hd__clkbuf_1
Xwire6710 svm0.counter\[9\] VGND VGND VPWR VPWR net6710 sky130_fd_sc_hd__buf_1
Xwire6721 net6722 VGND VGND VPWR VPWR net6721 sky130_fd_sc_hd__buf_1
XFILLER_0_163_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15180_ _07237_ _07239_ _07253_ VGND VGND VPWR VPWR _07254_ sky130_fd_sc_hd__a21o_1
X_24378_ _04227_ net1012 VGND VGND VPWR VPWR _04237_ sky130_fd_sc_hd__xnor2_1
Xwire6732 svm0.counter\[4\] VGND VGND VPWR VPWR net6732 sky130_fd_sc_hd__buf_1
Xwire7477 pid_q.state\[4\] VGND VGND VPWR VPWR net7477 sky130_fd_sc_hd__buf_1
Xfanout5936 net5942 VGND VGND VPWR VPWR net5936 sky130_fd_sc_hd__buf_1
Xwire6743 svm0.delta\[2\] VGND VGND VPWR VPWR net6743 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire7488 net7489 VGND VGND VPWR VPWR net7488 sky130_fd_sc_hd__buf_1
X_14131_ _06377_ _06392_ VGND VGND VPWR VPWR _06393_ sky130_fd_sc_hd__xor2_1
Xwire7499 net7500 VGND VGND VPWR VPWR net7499 sky130_fd_sc_hd__buf_1
Xwire6754 matmul0.state\[1\] VGND VGND VPWR VPWR net6754 sky130_fd_sc_hd__buf_1
Xfanout5958 pid_d.mult0.b\[0\] VGND VGND VPWR VPWR net5958 sky130_fd_sc_hd__buf_1
X_23329_ _03196_ net3059 VGND VGND VPWR VPWR _03199_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_162_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2463 net2465 VGND VGND VPWR VPWR net2463 sky130_fd_sc_hd__buf_1
XFILLER_0_104_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6787 cordic0.vec\[1\]\[17\] VGND VGND VPWR VPWR net6787 sky130_fd_sc_hd__clkbuf_1
X_14062_ _06307_ _06305_ _06324_ VGND VGND VPWR VPWR _06325_ sky130_fd_sc_hd__o21a_1
XFILLER_0_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13013_ net7246 _04892_ _04894_ net2991 net7546 VGND VGND VPWR VPWR _05286_ sky130_fd_sc_hd__a32o_1
X_18870_ net2589 _10677_ _10711_ VGND VGND VPWR VPWR _10712_ sky130_fd_sc_hd__nor3b_1
X_17821_ _09629_ _09659_ _09670_ _09671_ VGND VGND VPWR VPWR _09672_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold5 matmul0.matmul_stage_inst.a\[7\] VGND VGND VPWR VPWR net8958 sky130_fd_sc_hd__dlygate4sd3_1
X_17752_ _09601_ _09602_ VGND VGND VPWR VPWR _09603_ sky130_fd_sc_hd__xnor2_2
X_14964_ net4126 net4124 VGND VGND VPWR VPWR _07038_ sky130_fd_sc_hd__nor2_1
Xwire1050 _01302_ VGND VGND VPWR VPWR net1050 sky130_fd_sc_hd__buf_1
Xwire1061 net1062 VGND VGND VPWR VPWR net1061 sky130_fd_sc_hd__buf_1
X_16703_ net383 _08731_ VGND VGND VPWR VPWR _08732_ sky130_fd_sc_hd__xnor2_1
X_13915_ net1965 net1583 net7611 VGND VGND VPWR VPWR _06181_ sky130_fd_sc_hd__o21a_1
Xwire1072 _10356_ VGND VGND VPWR VPWR net1072 sky130_fd_sc_hd__clkbuf_1
X_17683_ svm0.tA\[15\] _09520_ _09562_ VGND VGND VPWR VPWR _09563_ sky130_fd_sc_hd__o21ai_1
Xwire1083 _08316_ VGND VGND VPWR VPWR net1083 sky130_fd_sc_hd__buf_1
Xwire1094 net1095 VGND VGND VPWR VPWR net1094 sky130_fd_sc_hd__buf_1
X_14895_ net6615 net6638 matmul0.matmul_stage_inst.f\[2\] VGND VGND VPWR VPWR _06969_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_187_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19422_ net6355 _10916_ VGND VGND VPWR VPWR _11259_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16634_ _08665_ _08666_ _08671_ VGND VGND VPWR VPWR _08672_ sky130_fd_sc_hd__a21o_1
X_13846_ _06106_ VGND VGND VPWR VPWR _06113_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19353_ net6288 net6203 VGND VGND VPWR VPWR _11190_ sky130_fd_sc_hd__or2b_1
XFILLER_0_174_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13777_ _05977_ _06043_ _06044_ VGND VGND VPWR VPWR _06045_ sky130_fd_sc_hd__a21o_1
X_16565_ _08581_ _08585_ VGND VGND VPWR VPWR _08624_ sky130_fd_sc_hd__nand2_1
XFILLER_0_168_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18304_ net6857 net6811 VGND VGND VPWR VPWR _10155_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15516_ net1272 _07588_ VGND VGND VPWR VPWR _07589_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_167_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8551 net8554 VGND VGND VPWR VPWR net8551 sky130_fd_sc_hd__buf_1
X_12728_ _04998_ _04999_ _05000_ VGND VGND VPWR VPWR _05001_ sky130_fd_sc_hd__and3_1
X_19284_ net6290 _11120_ _11049_ VGND VGND VPWR VPWR _11121_ sky130_fd_sc_hd__a21o_1
X_16496_ net2621 net2217 VGND VGND VPWR VPWR _08556_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout8573 net8578 VGND VGND VPWR VPWR net8573 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18235_ net7144 _10076_ _10079_ _10082_ _10085_ VGND VGND VPWR VPWR _10086_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_183_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12659_ net2335 VGND VGND VPWR VPWR _04932_ sky130_fd_sc_hd__buf_1
X_15447_ _07517_ _07520_ VGND VGND VPWR VPWR _07521_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_128_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18166_ net819 net818 _10013_ _10016_ VGND VGND VPWR VPWR _10017_ sky130_fd_sc_hd__a211o_1
X_15378_ _07437_ _07448_ _07451_ VGND VGND VPWR VPWR _07452_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17117_ _09058_ VGND VGND VPWR VPWR _09073_ sky130_fd_sc_hd__inv_2
Xwire380 _02513_ VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__clkbuf_1
X_14329_ net7346 net1299 net2896 pid_d.out\[2\] _06548_ VGND VGND VPWR VPWR _06549_
+ sky130_fd_sc_hd__a221o_1
X_18097_ _09856_ _09883_ VGND VGND VPWR VPWR _09948_ sky130_fd_sc_hd__xor2_1
Xwire391 net392 VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17048_ net2601 net5993 _08931_ net3326 VGND VGND VPWR VPWR _09007_ sky130_fd_sc_hd__o22a_1
XFILLER_0_110_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18999_ _10800_ VGND VGND VPWR VPWR _10836_ sky130_fd_sc_hd__buf_1
X_20961_ net5553 VGND VGND VPWR VPWR _00977_ sky130_fd_sc_hd__inv_2
XFILLER_0_174_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22700_ _02641_ net5478 net3095 VGND VGND VPWR VPWR _02642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23680_ _03455_ _03457_ _03546_ VGND VGND VPWR VPWR _03547_ sky130_fd_sc_hd__o21ai_1
X_20892_ _12521_ _12522_ VGND VGND VPWR VPWR _00908_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_177_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6729 svm0.counter\[5\] VGND VGND VPWR VPWR net6729 sky130_fd_sc_hd__buf_1
X_22631_ net3774 VGND VGND VPWR VPWR _02599_ sky130_fd_sc_hd__buf_1
XFILLER_0_49_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25350_ clknet_leaf_83_clk _00233_ net8502 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_22562_ net8887 net4301 net3774 VGND VGND VPWR VPWR _02546_ sky130_fd_sc_hd__and3_1
X_24301_ _04152_ _04160_ VGND VGND VPWR VPWR _04161_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21513_ net860 net806 net757 VGND VGND VPWR VPWR _01526_ sky130_fd_sc_hd__and3_1
X_25281_ clknet_leaf_92_clk _00164_ net8428 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.c\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22493_ _02481_ _02493_ VGND VGND VPWR VPWR _02494_ sky130_fd_sc_hd__xnor2_1
X_24232_ _04091_ _04092_ net4624 VGND VGND VPWR VPWR _04093_ sky130_fd_sc_hd__mux2_1
Xwire6006 net6003 VGND VGND VPWR VPWR net6006 sky130_fd_sc_hd__buf_1
X_21444_ net5724 net5565 VGND VGND VPWR VPWR _01457_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6017 net6014 VGND VGND VPWR VPWR net6017 sky130_fd_sc_hd__buf_1
XFILLER_0_90_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6039 net6040 VGND VGND VPWR VPWR net6039 sky130_fd_sc_hd__clkbuf_1
Xwire5305 net5306 VGND VGND VPWR VPWR net5305 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_82_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24163_ _03935_ _04023_ _04024_ VGND VGND VPWR VPWR _04025_ sky130_fd_sc_hd__o21ai_1
Xwire5316 net5317 VGND VGND VPWR VPWR net5316 sky130_fd_sc_hd__clkbuf_1
Xwire5327 pid_d.out\[13\] VGND VGND VPWR VPWR net5327 sky130_fd_sc_hd__dlymetal6s2s_1
X_21375_ _01263_ _01268_ _01261_ VGND VGND VPWR VPWR _01389_ sky130_fd_sc_hd__o21a_1
XFILLER_0_102_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5338 pid_d.out\[12\] VGND VGND VPWR VPWR net5338 sky130_fd_sc_hd__clkbuf_1
Xwire4604 net4605 VGND VGND VPWR VPWR net4604 sky130_fd_sc_hd__buf_1
Xwire5349 net5350 VGND VGND VPWR VPWR net5349 sky130_fd_sc_hd__clkbuf_1
Xwire4615 net4616 VGND VGND VPWR VPWR net4615 sky130_fd_sc_hd__buf_1
X_23114_ _02968_ net1677 VGND VGND VPWR VPWR _02984_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4626 net4627 VGND VGND VPWR VPWR net4626 sky130_fd_sc_hd__buf_1
X_20326_ net1911 _12128_ VGND VGND VPWR VPWR _12130_ sky130_fd_sc_hd__nor2_1
X_24094_ _03954_ net743 _03955_ VGND VGND VPWR VPWR _03956_ sky130_fd_sc_hd__o21a_1
Xwire4637 net4638 VGND VGND VPWR VPWR net4637 sky130_fd_sc_hd__buf_1
XFILLER_0_101_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4648 net4649 VGND VGND VPWR VPWR net4648 sky130_fd_sc_hd__clkbuf_1
Xwire3903 _10812_ VGND VGND VPWR VPWR net3903 sky130_fd_sc_hd__clkbuf_1
Xwire4659 net4660 VGND VGND VPWR VPWR net4659 sky130_fd_sc_hd__clkbuf_1
Xwire3914 net3917 VGND VGND VPWR VPWR net3914 sky130_fd_sc_hd__clkbuf_1
X_23045_ _02881_ _02914_ VGND VGND VPWR VPWR _02915_ sky130_fd_sc_hd__xnor2_2
Xwire3925 _10211_ VGND VGND VPWR VPWR net3925 sky130_fd_sc_hd__buf_1
X_20257_ net2 _12069_ VGND VGND VPWR VPWR _12070_ sky130_fd_sc_hd__xor2_1
Xwire3936 net3937 VGND VGND VPWR VPWR net3936 sky130_fd_sc_hd__buf_1
Xwire3947 net3948 VGND VGND VPWR VPWR net3947 sky130_fd_sc_hd__buf_1
Xwire3958 net3959 VGND VGND VPWR VPWR net3958 sky130_fd_sc_hd__clkbuf_1
Xwire3969 _09703_ VGND VGND VPWR VPWR net3969 sky130_fd_sc_hd__buf_1
X_20188_ _11995_ _12013_ VGND VGND VPWR VPWR _12014_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_192_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24996_ pid_q.out\[0\] net5183 VGND VGND VPWR VPWR _04754_ sky130_fd_sc_hd__xor2_1
XFILLER_0_188_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23947_ _03807_ _03810_ VGND VGND VPWR VPWR _03811_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_25_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length8654 net8655 VGND VGND VPWR VPWR net8654 sky130_fd_sc_hd__buf_1
X_13700_ net7615 net1338 net1563 VGND VGND VPWR VPWR _05969_ sky130_fd_sc_hd__a21oi_1
Xmax_length8665 net8667 VGND VGND VPWR VPWR net8665 sky130_fd_sc_hd__buf_1
Xmax_length8676 net8673 VGND VGND VPWR VPWR net8676 sky130_fd_sc_hd__buf_1
X_14680_ net7160 net7164 net7158 net7453 VGND VGND VPWR VPWR _06830_ sky130_fd_sc_hd__o31a_1
X_23878_ _03738_ _03741_ _03742_ VGND VGND VPWR VPWR _03743_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_6_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13631_ _05810_ _05811_ net7722 net1598 VGND VGND VPWR VPWR _05901_ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25617_ clknet_leaf_110_clk _00490_ net8343 VGND VGND VPWR VPWR cordic0.slte0.opA\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_22829_ net5365 net5983 VGND VGND VPWR VPWR _02730_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13562_ _05821_ _05832_ VGND VGND VPWR VPWR _05833_ sky130_fd_sc_hd__xnor2_2
X_16350_ _08408_ _08412_ VGND VGND VPWR VPWR _08413_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_149_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25548_ clknet_leaf_30_clk _00428_ net8673 VGND VGND VPWR VPWR pid_q.prev_int\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_181_Right_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15301_ _07373_ _07374_ VGND VGND VPWR VPWR _07375_ sky130_fd_sc_hd__xnor2_1
X_16281_ net1250 _08344_ VGND VGND VPWR VPWR _08345_ sky130_fd_sc_hd__xnor2_1
X_25479_ clknet_leaf_45_clk _00359_ net8787 VGND VGND VPWR VPWR svm0.tA\[1\] sky130_fd_sc_hd__dfrtp_1
X_13493_ _05645_ _05647_ _05763_ _05765_ VGND VGND VPWR VPWR _05766_ sky130_fd_sc_hd__a31o_1
XFILLER_0_81_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7230 net7231 VGND VGND VPWR VPWR net7230 sky130_fd_sc_hd__clkbuf_1
X_18020_ net7052 net7081 VGND VGND VPWR VPWR _09871_ sky130_fd_sc_hd__nor2_1
Xwire7241 net7242 VGND VGND VPWR VPWR net7241 sky130_fd_sc_hd__clkbuf_1
X_15232_ net3509 net3504 net4121 net4116 VGND VGND VPWR VPWR _07306_ sky130_fd_sc_hd__o22a_1
Xwire7252 net7253 VGND VGND VPWR VPWR net7252 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7263 matmul0.alpha_pass\[10\] VGND VGND VPWR VPWR net7263 sky130_fd_sc_hd__clkbuf_1
Xfanout6467 net6469 VGND VGND VPWR VPWR net6467 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_140_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout5744 net5754 VGND VGND VPWR VPWR net5744 sky130_fd_sc_hd__buf_1
Xwire7285 net7286 VGND VGND VPWR VPWR net7285 sky130_fd_sc_hd__clkbuf_1
X_15163_ _07232_ _07236_ VGND VGND VPWR VPWR _07237_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6551 net6552 VGND VGND VPWR VPWR net6551 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire7296 net7297 VGND VGND VPWR VPWR net7296 sky130_fd_sc_hd__clkbuf_1
Xwire6562 net6553 VGND VGND VPWR VPWR net6562 sky130_fd_sc_hd__buf_1
Xfanout5766 net5770 VGND VGND VPWR VPWR net5766 sky130_fd_sc_hd__buf_1
Xwire6573 net6574 VGND VGND VPWR VPWR net6573 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout5777 net5788 VGND VGND VPWR VPWR net5777 sky130_fd_sc_hd__buf_1
X_14114_ net834 _06375_ VGND VGND VPWR VPWR _06376_ sky130_fd_sc_hd__xnor2_1
Xwire5850 net5851 VGND VGND VPWR VPWR net5850 sky130_fd_sc_hd__clkbuf_1
X_19971_ _11797_ _11801_ VGND VGND VPWR VPWR _11802_ sky130_fd_sc_hd__xnor2_1
X_15094_ _07075_ _07167_ VGND VGND VPWR VPWR _07168_ sky130_fd_sc_hd__xnor2_1
Xwire6595 net6596 VGND VGND VPWR VPWR net6595 sky130_fd_sc_hd__buf_1
Xwire5861 net5865 VGND VGND VPWR VPWR net5861 sky130_fd_sc_hd__buf_1
Xwire5872 net5874 VGND VGND VPWR VPWR net5872 sky130_fd_sc_hd__buf_1
X_14045_ _06305_ _06308_ VGND VGND VPWR VPWR _06309_ sky130_fd_sc_hd__xnor2_2
X_18922_ _10717_ _10760_ _10761_ _10713_ VGND VGND VPWR VPWR _10762_ sky130_fd_sc_hd__a2bb2o_1
Xwire5894 net5888 VGND VGND VPWR VPWR net5894 sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_length1592 _05293_ VGND VGND VPWR VPWR net1592 sky130_fd_sc_hd__buf_1
XFILLER_0_66_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18853_ net352 _10695_ VGND VGND VPWR VPWR _10696_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17804_ net7061 _09613_ VGND VGND VPWR VPWR _09655_ sky130_fd_sc_hd__nor2_1
X_18784_ net1065 net1429 _10591_ VGND VGND VPWR VPWR _10628_ sky130_fd_sc_hd__a21bo_1
X_15996_ _08018_ _08063_ VGND VGND VPWR VPWR _08064_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_173_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17735_ net8052 net6509 _08943_ VGND VGND VPWR VPWR _09591_ sky130_fd_sc_hd__and3_1
X_14947_ net4146 VGND VGND VPWR VPWR _07021_ sky130_fd_sc_hd__clkbuf_1
X_17666_ net4013 svm0.tA\[1\] _09545_ net6740 VGND VGND VPWR VPWR _09546_ sky130_fd_sc_hd__a2bb2o_1
X_14878_ net9225 matmul0.matmul_stage_inst.f\[11\] net3604 VGND VGND VPWR VPWR _06957_
+ sky130_fd_sc_hd__mux2_1
X_19405_ _11092_ _11241_ VGND VGND VPWR VPWR _11242_ sky130_fd_sc_hd__xnor2_1
X_16617_ _08658_ VGND VGND VPWR VPWR _00247_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_187_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13829_ _06092_ _06095_ VGND VGND VPWR VPWR _06096_ sky130_fd_sc_hd__xnor2_2
X_17597_ svm0.tB\[6\] net6721 VGND VGND VPWR VPWR _09478_ sky130_fd_sc_hd__and2b_1
XFILLER_0_159_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19336_ net6259 net6230 _11159_ net1752 VGND VGND VPWR VPWR _11173_ sky130_fd_sc_hd__a31o_1
X_16548_ net2621 net2208 net2628 _08605_ VGND VGND VPWR VPWR _08607_ sky130_fd_sc_hd__a211o_1
XFILLER_0_45_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19267_ _11099_ _11102_ _11045_ VGND VGND VPWR VPWR _11104_ sky130_fd_sc_hd__a21oi_1
X_16479_ _08537_ _08539_ VGND VGND VPWR VPWR _08540_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18218_ net2545 VGND VGND VPWR VPWR _10069_ sky130_fd_sc_hd__inv_2
Xfanout7691 svm0.periodTop\[11\] VGND VGND VPWR VPWR net7691 sky130_fd_sc_hd__clkbuf_1
X_19198_ net6115 VGND VGND VPWR VPWR _11035_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18149_ _09954_ _09957_ VGND VGND VPWR VPWR _10000_ sky130_fd_sc_hd__nor2_1
Xhold202 svm0.tB\[0\] VGND VGND VPWR VPWR net9155 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold213 pid_q.out\[5\] VGND VGND VPWR VPWR net9166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 pid_q.prev_error\[0\] VGND VGND VPWR VPWR net9177 sky130_fd_sc_hd__dlygate4sd3_1
X_21160_ _01173_ _01175_ VGND VGND VPWR VPWR _01176_ sky130_fd_sc_hd__nand2_1
Xhold235 cordic0.slte0.opA\[8\] VGND VGND VPWR VPWR net9188 sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 svm0.calc_ready VGND VGND VPWR VPWR net9199 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold257 cordic0.cos\[11\] VGND VGND VPWR VPWR net9210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 pid_q.prev_int\[7\] VGND VGND VPWR VPWR net9221 sky130_fd_sc_hd__dlygate4sd3_1
X_20111_ net6052 _11938_ VGND VGND VPWR VPWR _11939_ sky130_fd_sc_hd__and2_1
Xhold279 svm0.tA\[11\] VGND VGND VPWR VPWR net9232 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21091_ net5564 _01079_ _01080_ VGND VGND VPWR VPWR _01107_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2509 net2510 VGND VGND VPWR VPWR net2509 sky130_fd_sc_hd__clkbuf_2
X_20042_ _11870_ _11871_ VGND VGND VPWR VPWR _11872_ sky130_fd_sc_hd__xor2_2
Xwire1808 net1809 VGND VGND VPWR VPWR net1808 sky130_fd_sc_hd__buf_1
Xwire1819 net1820 VGND VGND VPWR VPWR net1819 sky130_fd_sc_hd__buf_1
X_24850_ net7488 _04540_ net227 VGND VGND VPWR VPWR _04658_ sky130_fd_sc_hd__and3_1
X_23801_ _03664_ _03665_ VGND VGND VPWR VPWR _03667_ sky130_fd_sc_hd__or2_1
X_24781_ net7974 VGND VGND VPWR VPWR _04608_ sky130_fd_sc_hd__inv_2
X_21993_ _01892_ _01896_ VGND VGND VPWR VPWR _02001_ sky130_fd_sc_hd__or2_1
X_23732_ _03595_ _03597_ VGND VGND VPWR VPWR _03598_ sky130_fd_sc_hd__xnor2_1
X_20944_ net5779 net5804 VGND VGND VPWR VPWR _00960_ sky130_fd_sc_hd__and2_1
X_23663_ _03526_ _03529_ VGND VGND VPWR VPWR _03530_ sky130_fd_sc_hd__xnor2_1
X_20875_ _00880_ net2482 VGND VGND VPWR VPWR _00891_ sky130_fd_sc_hd__or2_1
X_22614_ net7250 net7237 net7227 _02576_ VGND VGND VPWR VPWR _02586_ sky130_fd_sc_hd__or4_1
X_25402_ clknet_leaf_69_clk _00285_ net8450 VGND VGND VPWR VPWR matmul0.a\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length5836 net5837 VGND VGND VPWR VPWR net5836 sky130_fd_sc_hd__buf_1
X_23594_ _03451_ _03461_ VGND VGND VPWR VPWR _03462_ sky130_fd_sc_hd__xor2_1
XFILLER_0_76_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25333_ clknet_leaf_82_clk _00216_ net8503 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult1\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_22545_ pid_d.curr_error\[10\] net3016 net2461 VGND VGND VPWR VPWR _02535_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25264_ clknet_leaf_88_clk _00147_ net8435 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.b\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_22476_ net2055 _02476_ VGND VGND VPWR VPWR _02477_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_161_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24215_ net3743 _03887_ VGND VGND VPWR VPWR _04076_ sky130_fd_sc_hd__nand2_1
X_21427_ _01438_ _01439_ VGND VGND VPWR VPWR _01440_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_101_Left_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5113 net5114 VGND VGND VPWR VPWR net5113 sky130_fd_sc_hd__clkbuf_1
X_25195_ clknet_leaf_62_clk _00084_ net8708 VGND VGND VPWR VPWR matmul0.b_in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire5124 net5125 VGND VGND VPWR VPWR net5124 sky130_fd_sc_hd__buf_1
XFILLER_0_133_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5135 net5136 VGND VGND VPWR VPWR net5135 sky130_fd_sc_hd__buf_1
X_24146_ net4605 net4625 net3052 net4788 _04007_ VGND VGND VPWR VPWR _04008_ sky130_fd_sc_hd__a32o_1
Xwire4401 pid_q.out\[13\] VGND VGND VPWR VPWR net4401 sky130_fd_sc_hd__clkbuf_2
Xwire5157 net5158 VGND VGND VPWR VPWR net5157 sky130_fd_sc_hd__buf_1
Xwire4412 pid_q.out\[12\] VGND VGND VPWR VPWR net4412 sky130_fd_sc_hd__clkbuf_1
X_21358_ net1729 _01371_ VGND VGND VPWR VPWR _01372_ sky130_fd_sc_hd__xnor2_1
Xwire5168 pid_q.curr_error\[1\] VGND VGND VPWR VPWR net5168 sky130_fd_sc_hd__clkbuf_2
Xwire4423 pid_q.out\[10\] VGND VGND VPWR VPWR net4423 sky130_fd_sc_hd__clkbuf_1
Xwire5179 net5180 VGND VGND VPWR VPWR net5179 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4434 net4435 VGND VGND VPWR VPWR net4434 sky130_fd_sc_hd__clkbuf_1
Xwire3700 net3701 VGND VGND VPWR VPWR net3700 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4445 net4446 VGND VGND VPWR VPWR net4445 sky130_fd_sc_hd__clkbuf_1
Xwire3711 net3712 VGND VGND VPWR VPWR net3711 sky130_fd_sc_hd__clkbuf_2
X_20309_ _12102_ _12113_ VGND VGND VPWR VPWR _12114_ sky130_fd_sc_hd__nand2_1
X_24077_ _03837_ _03844_ _03842_ VGND VGND VPWR VPWR _03940_ sky130_fd_sc_hd__o21ai_1
Xwire4456 pid_q.out\[4\] VGND VGND VPWR VPWR net4456 sky130_fd_sc_hd__clkbuf_1
Xwire3722 net3723 VGND VGND VPWR VPWR net3722 sky130_fd_sc_hd__clkbuf_1
Xwire4467 net4468 VGND VGND VPWR VPWR net4467 sky130_fd_sc_hd__clkbuf_1
X_21289_ net1737 net1736 _01303_ VGND VGND VPWR VPWR _01304_ sky130_fd_sc_hd__o21a_2
Xwire4478 pid_q.kp\[5\] VGND VGND VPWR VPWR net4478 sky130_fd_sc_hd__clkbuf_1
Xwire3733 _04172_ VGND VGND VPWR VPWR net3733 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4489 net4490 VGND VGND VPWR VPWR net4489 sky130_fd_sc_hd__buf_1
Xwire3744 net3745 VGND VGND VPWR VPWR net3744 sky130_fd_sc_hd__buf_1
X_23028_ _02895_ _02896_ _02897_ VGND VGND VPWR VPWR _02898_ sky130_fd_sc_hd__o21a_1
Xwire3755 net3756 VGND VGND VPWR VPWR net3755 sky130_fd_sc_hd__clkbuf_1
Xwire3766 _02659_ VGND VGND VPWR VPWR net3766 sky130_fd_sc_hd__clkbuf_1
Xwire3777 net3779 VGND VGND VPWR VPWR net3777 sky130_fd_sc_hd__clkbuf_1
Xwire3788 _01709_ VGND VGND VPWR VPWR net3788 sky130_fd_sc_hd__buf_1
Xwire3799 net3800 VGND VGND VPWR VPWR net3799 sky130_fd_sc_hd__clkbuf_1
X_15850_ _07914_ _07918_ VGND VGND VPWR VPWR _07920_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14801_ net9019 net3006 _06917_ VGND VGND VPWR VPWR _00172_ sky130_fd_sc_hd__o21a_1
X_15781_ _07762_ _07764_ _07760_ VGND VGND VPWR VPWR _07851_ sky130_fd_sc_hd__o21a_1
X_24979_ _04744_ VGND VGND VPWR VPWR _00769_ sky130_fd_sc_hd__clkbuf_1
X_12993_ net7802 net2324 net2320 VGND VGND VPWR VPWR _05266_ sky130_fd_sc_hd__and3_1
X_17520_ _09319_ _09400_ _09404_ VGND VGND VPWR VPWR _09405_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_19_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14732_ net7444 net7160 VGND VGND VPWR VPWR _06868_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length8484 net8485 VGND VGND VPWR VPWR net8484 sky130_fd_sc_hd__buf_1
XFILLER_0_169_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17451_ net6736 _09345_ _09346_ _09344_ VGND VGND VPWR VPWR _00393_ sky130_fd_sc_hd__a22o_1
X_14663_ net8982 _06814_ _06816_ VGND VGND VPWR VPWR _00135_ sky130_fd_sc_hd__a21o_1
X_16402_ _08453_ net1246 VGND VGND VPWR VPWR _08464_ sky130_fd_sc_hd__xnor2_2
X_13614_ net7790 net2950 net3669 VGND VGND VPWR VPWR _05884_ sky130_fd_sc_hd__and3_1
X_17382_ svm0.delta\[5\] VGND VGND VPWR VPWR _09291_ sky130_fd_sc_hd__inv_2
X_14594_ _06761_ _06766_ _06767_ net281 VGND VGND VPWR VPWR _06768_ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19121_ net2112 net2111 _10957_ VGND VGND VPWR VPWR _10958_ sky130_fd_sc_hd__nand3_1
XFILLER_0_27_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16333_ _08394_ _08395_ VGND VGND VPWR VPWR _08396_ sky130_fd_sc_hd__nor2_1
X_13545_ net7698 net1352 _05745_ _05746_ VGND VGND VPWR VPWR _05816_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_54_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6220 net6223 VGND VGND VPWR VPWR net6220 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_109_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19052_ net2117 _10888_ VGND VGND VPWR VPWR _10889_ sky130_fd_sc_hd__nor2_1
X_13476_ net1574 net1572 net1945 VGND VGND VPWR VPWR _05749_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16264_ _08326_ _08327_ VGND VGND VPWR VPWR _08328_ sky130_fd_sc_hd__nor2_1
Xfanout6253 cordic0.vec\[0\]\[5\] VGND VGND VPWR VPWR net6253 sky130_fd_sc_hd__buf_1
X_18003_ _09026_ net2555 VGND VGND VPWR VPWR _09854_ sky130_fd_sc_hd__xnor2_1
Xfanout6264 net6273 VGND VGND VPWR VPWR net6264 sky130_fd_sc_hd__clkbuf_1
Xwire7060 net7061 VGND VGND VPWR VPWR net7060 sky130_fd_sc_hd__buf_1
Xfanout6275 net6285 VGND VGND VPWR VPWR net6275 sky130_fd_sc_hd__buf_1
X_15215_ _07272_ _07273_ VGND VGND VPWR VPWR _07289_ sky130_fd_sc_hd__xnor2_1
Xfanout5541 net5554 VGND VGND VPWR VPWR net5541 sky130_fd_sc_hd__buf_1
Xwire7082 net7083 VGND VGND VPWR VPWR net7082 sky130_fd_sc_hd__buf_1
XFILLER_0_180_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6286 net6301 VGND VGND VPWR VPWR net6286 sky130_fd_sc_hd__clkbuf_1
X_16195_ net2682 net2670 _07932_ _08257_ VGND VGND VPWR VPWR _08260_ sky130_fd_sc_hd__a211o_1
XFILLER_0_22_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout6297 net6302 VGND VGND VPWR VPWR net6297 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5563 net5568 VGND VGND VPWR VPWR net5563 sky130_fd_sc_hd__clkbuf_1
Xwire6370 cordic0.slte0.opA\[12\] VGND VGND VPWR VPWR net6370 sky130_fd_sc_hd__buf_1
XFILLER_0_164_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15146_ net2251 net2790 VGND VGND VPWR VPWR _07220_ sky130_fd_sc_hd__nand2_1
Xwire6381 net6382 VGND VGND VPWR VPWR net6381 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire6392 cordic0.slte0.opB\[15\] VGND VGND VPWR VPWR net6392 sky130_fd_sc_hd__clkbuf_1
Xfanout4862 net4883 VGND VGND VPWR VPWR net4862 sky130_fd_sc_hd__buf_1
XFILLER_0_11_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5680 net5673 VGND VGND VPWR VPWR net5680 sky130_fd_sc_hd__buf_1
X_19954_ _11736_ _11785_ VGND VGND VPWR VPWR _11786_ sky130_fd_sc_hd__xnor2_1
X_15077_ _07135_ VGND VGND VPWR VPWR _07151_ sky130_fd_sc_hd__clkbuf_2
Xwire5691 net5692 VGND VGND VPWR VPWR net5691 sky130_fd_sc_hd__buf_1
X_14028_ net7625 _05608_ _05609_ VGND VGND VPWR VPWR _06292_ sky130_fd_sc_hd__and3_1
X_18905_ _10743_ _10745_ VGND VGND VPWR VPWR _10746_ sky130_fd_sc_hd__xnor2_1
Xwire4990 net4991 VGND VGND VPWR VPWR net4990 sky130_fd_sc_hd__buf_1
X_19885_ _11544_ _11545_ _11609_ VGND VGND VPWR VPWR _11718_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18836_ _10676_ _10678_ VGND VGND VPWR VPWR _10679_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18767_ _10610_ _10611_ VGND VGND VPWR VPWR _10612_ sky130_fd_sc_hd__or2_1
X_15979_ _07935_ _07938_ _08046_ VGND VGND VPWR VPWR _08047_ sky130_fd_sc_hd__o21a_1
X_17718_ net9223 net1216 net1453 pid_q.curr_int\[9\] VGND VGND VPWR VPWR _00423_ sky130_fd_sc_hd__a22o_1
X_18698_ net1430 _10543_ VGND VGND VPWR VPWR _10544_ sky130_fd_sc_hd__xor2_1
XFILLER_0_188_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17649_ net6707 net6746 VGND VGND VPWR VPWR _09529_ sky130_fd_sc_hd__or2_1
XFILLER_0_175_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20660_ net1837 _12437_ net8061 VGND VGND VPWR VPWR _12438_ sky130_fd_sc_hd__o21a_1
XFILLER_0_85_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19319_ net6186 _10930_ VGND VGND VPWR VPWR _11156_ sky130_fd_sc_hd__xor2_2
XFILLER_0_46_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20591_ net1237 _12372_ net3164 VGND VGND VPWR VPWR _12374_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22330_ pid_d.curr_int\[12\] net4391 net381 VGND VGND VPWR VPWR _02333_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_144_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22261_ pid_d.prev_error\[11\] net5966 VGND VGND VPWR VPWR _02265_ sky130_fd_sc_hd__nor2_1
XFILLER_0_170_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24000_ _03860_ _03773_ _03862_ VGND VGND VPWR VPWR _03863_ sky130_fd_sc_hd__a21o_1
X_21212_ _01009_ _01227_ _01022_ VGND VGND VPWR VPWR _01228_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_13_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22192_ _02059_ _02196_ net859 VGND VGND VPWR VPWR _02197_ sky130_fd_sc_hd__or3b_1
Xwire3007 net3008 VGND VGND VPWR VPWR net3007 sky130_fd_sc_hd__buf_1
X_21143_ net3816 _01151_ VGND VGND VPWR VPWR _01159_ sky130_fd_sc_hd__nor2_1
Xwire3018 _04874_ VGND VGND VPWR VPWR net3018 sky130_fd_sc_hd__buf_1
Xwire3029 _04857_ VGND VGND VPWR VPWR net3029 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_6_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2306 _05130_ VGND VGND VPWR VPWR net2306 sky130_fd_sc_hd__clkbuf_1
Xwire2317 net2318 VGND VGND VPWR VPWR net2317 sky130_fd_sc_hd__buf_1
X_21074_ _01045_ _01089_ VGND VGND VPWR VPWR _01090_ sky130_fd_sc_hd__xnor2_2
Xwire2328 net2329 VGND VGND VPWR VPWR net2328 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2339 _04930_ VGND VGND VPWR VPWR net2339 sky130_fd_sc_hd__buf_1
Xwire1605 net1606 VGND VGND VPWR VPWR net1605 sky130_fd_sc_hd__buf_1
X_24902_ _04692_ net4492 net2399 VGND VGND VPWR VPWR _04693_ sky130_fd_sc_hd__mux2_1
Xwire1616 net1617 VGND VGND VPWR VPWR net1616 sky130_fd_sc_hd__buf_1
X_20025_ net6081 _11797_ _11800_ VGND VGND VPWR VPWR _11855_ sky130_fd_sc_hd__nor3_1
X_25882_ clknet_leaf_16_clk _00755_ net8625 VGND VGND VPWR VPWR pid_q.ki\[10\] sky130_fd_sc_hd__dfrtp_1
Xwire1627 _04785_ VGND VGND VPWR VPWR net1627 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1638 net1639 VGND VGND VPWR VPWR net1638 sky130_fd_sc_hd__buf_1
Xwire1649 net1650 VGND VGND VPWR VPWR net1649 sky130_fd_sc_hd__clkbuf_2
X_24833_ net5021 _04642_ net2000 net922 VGND VGND VPWR VPWR _00718_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24764_ net7990 _04588_ _04592_ VGND VGND VPWR VPWR _04593_ sky130_fd_sc_hd__o21ai_2
X_21976_ _01799_ net1044 VGND VGND VPWR VPWR _01984_ sky130_fd_sc_hd__xor2_1
XFILLER_0_96_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23715_ pid_q.curr_int\[4\] pid_q.prev_int\[4\] VGND VGND VPWR VPWR _03581_ sky130_fd_sc_hd__xor2_1
Xmax_length7057 net7053 VGND VGND VPWR VPWR net7057 sky130_fd_sc_hd__clkbuf_2
X_20927_ _00939_ _00940_ _00942_ VGND VGND VPWR VPWR _00943_ sky130_fd_sc_hd__a21boi_2
X_24695_ net3727 net3034 VGND VGND VPWR VPWR _04533_ sky130_fd_sc_hd__nor2_1
Xmax_length6334 net6335 VGND VGND VPWR VPWR net6334 sky130_fd_sc_hd__buf_1
XFILLER_0_49_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6356 net6357 VGND VGND VPWR VPWR net6356 sky130_fd_sc_hd__buf_1
X_23646_ net4530 net5078 VGND VGND VPWR VPWR _03513_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length6367 cordic0.vec\[0\]\[0\] VGND VGND VPWR VPWR net6367 sky130_fd_sc_hd__clkbuf_1
X_20858_ _00864_ _00873_ VGND VGND VPWR VPWR _00874_ sky130_fd_sc_hd__xor2_1
XFILLER_0_187_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length5644 net5639 VGND VGND VPWR VPWR net5644 sky130_fd_sc_hd__buf_1
XFILLER_0_64_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23577_ _03439_ _03444_ VGND VGND VPWR VPWR _03445_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_147_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_115_clk clknet_4_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_115_clk
+ sky130_fd_sc_hd__clkbuf_16
Xmax_length4943 net4944 VGND VGND VPWR VPWR net4943 sky130_fd_sc_hd__clkbuf_1
X_20789_ net5615 net5741 VGND VGND VPWR VPWR _12560_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length5688 net5685 VGND VGND VPWR VPWR net5688 sky130_fd_sc_hd__buf_1
Xwire902 net903 VGND VGND VPWR VPWR net902 sky130_fd_sc_hd__clkbuf_2
Xwire913 net914 VGND VGND VPWR VPWR net913 sky130_fd_sc_hd__buf_1
X_13330_ _05595_ _05602_ VGND VGND VPWR VPWR _05603_ sky130_fd_sc_hd__xor2_1
XFILLER_0_18_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire924 net925 VGND VGND VPWR VPWR net924 sky130_fd_sc_hd__clkbuf_1
X_25316_ clknet_leaf_75_clk _00199_ net8463 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.f\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_22528_ net9182 net1699 _02526_ VGND VGND VPWR VPWR _00536_ sky130_fd_sc_hd__a21o_1
Xwire935 net936 VGND VGND VPWR VPWR net935 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire946 _01734_ VGND VGND VPWR VPWR net946 sky130_fd_sc_hd__buf_1
Xwire957 _11598_ VGND VGND VPWR VPWR net957 sky130_fd_sc_hd__clkbuf_1
X_13261_ net7879 net3684 net4254 VGND VGND VPWR VPWR _05534_ sky130_fd_sc_hd__and3_1
Xwire968 net969 VGND VGND VPWR VPWR net968 sky130_fd_sc_hd__clkbuf_1
X_22459_ pid_d.curr_int\[14\] _12499_ net2488 _02408_ _02460_ VGND VGND VPWR VPWR
+ _00533_ sky130_fd_sc_hd__a221o_1
X_25247_ clknet_leaf_87_clk _00130_ net8436 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.a\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire979 net980 VGND VGND VPWR VPWR net979 sky130_fd_sc_hd__buf_1
XFILLER_0_150_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15000_ net1896 _07060_ VGND VGND VPWR VPWR _07074_ sky130_fd_sc_hd__xor2_1
XFILLER_0_33_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13192_ _05463_ _05448_ _05449_ VGND VGND VPWR VPWR _05465_ sky130_fd_sc_hd__nand3_1
X_25178_ clknet_leaf_72_clk _00067_ net8469 VGND VGND VPWR VPWR matmul0.a_in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire4220 _06963_ VGND VGND VPWR VPWR net4220 sky130_fd_sc_hd__buf_1
X_24129_ net2408 _03990_ VGND VGND VPWR VPWR _03991_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4242 net4243 VGND VGND VPWR VPWR net4242 sky130_fd_sc_hd__clkbuf_1
Xwire4253 _05776_ VGND VGND VPWR VPWR net4253 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_138_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3530 net3531 VGND VGND VPWR VPWR net3530 sky130_fd_sc_hd__clkbuf_1
Xwire4275 _04898_ VGND VGND VPWR VPWR net4275 sky130_fd_sc_hd__clkbuf_1
X_16951_ _08913_ VGND VGND VPWR VPWR _08914_ sky130_fd_sc_hd__buf_1
Xwire3541 net3542 VGND VGND VPWR VPWR net3541 sky130_fd_sc_hd__buf_1
Xwire4286 _04883_ VGND VGND VPWR VPWR net4286 sky130_fd_sc_hd__buf_1
Xwire4297 _04872_ VGND VGND VPWR VPWR net4297 sky130_fd_sc_hd__buf_1
Xwire3552 net3553 VGND VGND VPWR VPWR net3552 sky130_fd_sc_hd__buf_1
Xwire3563 net3564 VGND VGND VPWR VPWR net3563 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3574 net3576 VGND VGND VPWR VPWR net3574 sky130_fd_sc_hd__buf_1
X_15902_ net2846 net2695 net3439 net2803 VGND VGND VPWR VPWR _07971_ sky130_fd_sc_hd__a211o_1
Xwire3585 net3586 VGND VGND VPWR VPWR net3585 sky130_fd_sc_hd__buf_1
Xwire2840 net2841 VGND VGND VPWR VPWR net2840 sky130_fd_sc_hd__buf_1
X_19670_ net6113 net6136 VGND VGND VPWR VPWR _11506_ sky130_fd_sc_hd__nand2_1
Xwire2851 net2852 VGND VGND VPWR VPWR net2851 sky130_fd_sc_hd__buf_1
XFILLER_0_194_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16882_ net6133 net6092 net6504 VGND VGND VPWR VPWR _08846_ sky130_fd_sc_hd__mux2_1
Xwire2862 _06838_ VGND VGND VPWR VPWR net2862 sky130_fd_sc_hd__buf_1
Xwire2873 net2875 VGND VGND VPWR VPWR net2873 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2884 net2885 VGND VGND VPWR VPWR net2884 sky130_fd_sc_hd__clkbuf_1
X_18621_ net3959 _10429_ _10223_ VGND VGND VPWR VPWR _10468_ sky130_fd_sc_hd__mux2_1
Xwire2895 _06569_ VGND VGND VPWR VPWR net2895 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15833_ _07897_ _07899_ _07902_ VGND VGND VPWR VPWR _07903_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18552_ net607 _10333_ net765 _10400_ VGND VGND VPWR VPWR _10401_ sky130_fd_sc_hd__a31o_1
X_15764_ net3499 net3399 VGND VGND VPWR VPWR _07834_ sky130_fd_sc_hd__nor2_1
X_12976_ net7785 net1355 VGND VGND VPWR VPWR _05249_ sky130_fd_sc_hd__nand2_1
X_17503_ _09258_ _09390_ VGND VGND VPWR VPWR _09391_ sky130_fd_sc_hd__nor2_1
X_14715_ net7456 _06855_ VGND VGND VPWR VPWR _06856_ sky130_fd_sc_hd__nand2_1
X_18483_ _10331_ net663 net659 VGND VGND VPWR VPWR _10333_ sky130_fd_sc_hd__and3_1
X_15695_ _07760_ _07765_ VGND VGND VPWR VPWR _07766_ sky130_fd_sc_hd__xnor2_1
X_17434_ net4067 VGND VGND VPWR VPWR _09332_ sky130_fd_sc_hd__buf_1
X_14646_ net8969 net2879 _06807_ VGND VGND VPWR VPWR _00127_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17365_ net7377 svm0.delta\[1\] _09276_ VGND VGND VPWR VPWR _09277_ sky130_fd_sc_hd__o21a_1
XFILLER_0_172_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_106_clk clknet_4_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_106_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_7_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14577_ net7244 net5213 VGND VGND VPWR VPWR _06753_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19104_ net6340 net6353 VGND VGND VPWR VPWR _10941_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16316_ _08318_ _08351_ _08310_ VGND VGND VPWR VPWR _08379_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_166_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13528_ _05704_ net1128 VGND VGND VPWR VPWR _05799_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17296_ net7787 _09209_ VGND VGND VPWR VPWR _09210_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19035_ net6204 net6154 _10871_ VGND VGND VPWR VPWR _10872_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16247_ net979 _08287_ _08286_ VGND VGND VPWR VPWR _08311_ sky130_fd_sc_hd__a21oi_2
X_13459_ net7710 net2321 net2317 VGND VGND VPWR VPWR _05732_ sky130_fd_sc_hd__and3_1
XFILLER_0_153_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16178_ _08226_ _08229_ _08242_ VGND VGND VPWR VPWR _08243_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15129_ _07183_ net1278 VGND VGND VPWR VPWR _07203_ sky130_fd_sc_hd__nor2_1
Xfanout4692 net4714 VGND VGND VPWR VPWR net4692 sky130_fd_sc_hd__buf_1
X_19937_ net3137 net2096 VGND VGND VPWR VPWR _11769_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19868_ _11700_ VGND VGND VPWR VPWR _11701_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18819_ _10627_ _10649_ _10650_ VGND VGND VPWR VPWR _10662_ sky130_fd_sc_hd__a21o_1
X_19799_ net2104 _11582_ net6151 VGND VGND VPWR VPWR _11633_ sky130_fd_sc_hd__a21o_1
X_21830_ net5719 net5499 VGND VGND VPWR VPWR _01839_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21761_ _01673_ _01675_ VGND VGND VPWR VPWR _01771_ sky130_fd_sc_hd__nand2_1
XFILLER_0_194_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23500_ _03349_ _03368_ VGND VGND VPWR VPWR _03369_ sky130_fd_sc_hd__xor2_1
X_20712_ _12481_ _12484_ VGND VGND VPWR VPWR _12485_ sky130_fd_sc_hd__xor2_1
X_24480_ _04333_ _04336_ VGND VGND VPWR VPWR _04337_ sky130_fd_sc_hd__xnor2_1
X_21692_ net1720 _01702_ VGND VGND VPWR VPWR _01703_ sky130_fd_sc_hd__nor2_1
Xwire8508 net8509 VGND VGND VPWR VPWR net8508 sky130_fd_sc_hd__buf_1
Xwire8519 net8520 VGND VGND VPWR VPWR net8519 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23431_ net1675 net3059 _03300_ VGND VGND VPWR VPWR _03301_ sky130_fd_sc_hd__a21o_1
XFILLER_0_190_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20643_ net6164 _12412_ _12411_ VGND VGND VPWR VPWR _12422_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire7807 net7811 VGND VGND VPWR VPWR net7807 sky130_fd_sc_hd__buf_1
Xwire7818 net7812 VGND VGND VPWR VPWR net7818 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire209 net210 VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__buf_1
Xwire7829 net7830 VGND VGND VPWR VPWR net7829 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23362_ net2026 net1678 VGND VGND VPWR VPWR _03232_ sky130_fd_sc_hd__nand2_1
X_20574_ _12356_ _12348_ _12349_ VGND VGND VPWR VPWR _12358_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_61_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22313_ _02313_ _02316_ VGND VGND VPWR VPWR _02317_ sky130_fd_sc_hd__xnor2_1
X_25101_ _04836_ _04839_ net4400 VGND VGND VPWR VPWR _04844_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_2_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2826 _07087_ VGND VGND VPWR VPWR net2826 sky130_fd_sc_hd__buf_1
X_23293_ net1031 _03162_ VGND VGND VPWR VPWR _03163_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25032_ _04784_ VGND VGND VPWR VPWR _04785_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22244_ _02245_ _02247_ VGND VGND VPWR VPWR _02249_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22175_ net4381 _02113_ _02173_ net4314 net410 VGND VGND VPWR VPWR _02181_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21126_ _01141_ _01100_ VGND VGND VPWR VPWR _01142_ sky130_fd_sc_hd__xnor2_1
Xwire2103 _11402_ VGND VGND VPWR VPWR net2103 sky130_fd_sc_hd__buf_1
Xwire2114 net2115 VGND VGND VPWR VPWR net2114 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2125 _10588_ VGND VGND VPWR VPWR net2125 sky130_fd_sc_hd__buf_1
Xwire2136 net2137 VGND VGND VPWR VPWR net2136 sky130_fd_sc_hd__clkbuf_1
X_25934_ clknet_leaf_25_clk _00807_ net8583 VGND VGND VPWR VPWR pid_d.prev_int\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire2147 net2148 VGND VGND VPWR VPWR net2147 sky130_fd_sc_hd__clkbuf_2
Xwire1402 net1403 VGND VGND VPWR VPWR net1402 sky130_fd_sc_hd__clkbuf_1
X_21057_ net3823 net3121 _01060_ _01001_ VGND VGND VPWR VPWR _01073_ sky130_fd_sc_hd__o211a_1
Xwire2158 _09193_ VGND VGND VPWR VPWR net2158 sky130_fd_sc_hd__buf_1
Xwire1413 net1414 VGND VGND VPWR VPWR net1413 sky130_fd_sc_hd__clkbuf_1
Xwire1424 net1425 VGND VGND VPWR VPWR net1424 sky130_fd_sc_hd__clkbuf_1
Xwire2169 _09081_ VGND VGND VPWR VPWR net2169 sky130_fd_sc_hd__clkbuf_1
Xwire1435 _10418_ VGND VGND VPWR VPWR net1435 sky130_fd_sc_hd__clkbuf_1
X_20008_ _11835_ _11837_ net487 VGND VGND VPWR VPWR _11838_ sky130_fd_sc_hd__mux2_1
X_25865_ clknet_leaf_16_clk _00738_ net8619 VGND VGND VPWR VPWR pid_q.mult0.a\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1457 _09579_ VGND VGND VPWR VPWR net1457 sky130_fd_sc_hd__buf_1
Xwire1468 net1469 VGND VGND VPWR VPWR net1468 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24816_ net1626 _04634_ _04637_ _04638_ VGND VGND VPWR VPWR _04639_ sky130_fd_sc_hd__a31oi_1
X_12830_ net7906 net1603 VGND VGND VPWR VPWR _05103_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25796_ clknet_leaf_33_clk _00669_ net8679 VGND VGND VPWR VPWR pid_q.curr_int\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_68_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24747_ net8002 _04572_ _04577_ VGND VGND VPWR VPWR _04578_ sky130_fd_sc_hd__a21o_1
X_12761_ net7823 _04904_ net2989 VGND VGND VPWR VPWR _05034_ sky130_fd_sc_hd__and3_2
XFILLER_0_33_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21959_ net5817 _01963_ _01966_ VGND VGND VPWR VPWR _01967_ sky130_fd_sc_hd__a21o_1
Xmax_length6131 net6127 VGND VGND VPWR VPWR net6131 sky130_fd_sc_hd__buf_1
XFILLER_0_57_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14500_ _06679_ _06682_ VGND VGND VPWR VPWR _06683_ sky130_fd_sc_hd__xnor2_1
X_12692_ _04964_ VGND VGND VPWR VPWR _04965_ sky130_fd_sc_hd__clkbuf_1
X_15480_ _07543_ _07553_ VGND VGND VPWR VPWR _07554_ sky130_fd_sc_hd__xor2_1
XFILLER_0_16_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24678_ net9127 net1648 _04521_ VGND VGND VPWR VPWR _00691_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14431_ _06627_ VGND VGND VPWR VPWR _00092_ sky130_fd_sc_hd__clkbuf_1
X_23629_ net4641 net4940 _03494_ _03495_ VGND VGND VPWR VPWR _03496_ sky130_fd_sc_hd__a31o_1
Xmax_length6197 net6198 VGND VGND VPWR VPWR net6197 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length4740 net4734 VGND VGND VPWR VPWR net4740 sky130_fd_sc_hd__buf_1
XFILLER_0_126_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17150_ net6932 _09075_ _09076_ _09103_ _09064_ VGND VGND VPWR VPWR _09104_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_135_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14362_ net1548 VGND VGND VPWR VPWR _06574_ sky130_fd_sc_hd__buf_1
Xwire710 net711 VGND VGND VPWR VPWR net710 sky130_fd_sc_hd__clkbuf_1
Xwire721 net722 VGND VGND VPWR VPWR net721 sky130_fd_sc_hd__clkbuf_1
Xwire732 _05517_ VGND VGND VPWR VPWR net732 sky130_fd_sc_hd__clkbuf_2
Xinput17 currA_in[0] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
Xwire743 _03863_ VGND VGND VPWR VPWR net743 sky130_fd_sc_hd__buf_1
Xinput28 currA_in[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
X_16101_ _08105_ _08165_ net1515 net1526 VGND VGND VPWR VPWR _08167_ sky130_fd_sc_hd__a211o_1
Xwire754 _03240_ VGND VGND VPWR VPWR net754 sky130_fd_sc_hd__clkbuf_1
X_13313_ net7698 net1982 net2360 VGND VGND VPWR VPWR _05586_ sky130_fd_sc_hd__and3_1
Xinput39 currB_in[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
X_14293_ net67 net2901 net2264 net7684 VGND VGND VPWR VPWR _00062_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17081_ net1478 _09038_ VGND VGND VPWR VPWR _09039_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_24_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire765 net766 VGND VGND VPWR VPWR net765 sky130_fd_sc_hd__clkbuf_2
Xwire776 net777 VGND VGND VPWR VPWR net776 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire787 net788 VGND VGND VPWR VPWR net787 sky130_fd_sc_hd__clkbuf_1
Xwire798 net799 VGND VGND VPWR VPWR net798 sky130_fd_sc_hd__clkbuf_1
X_13244_ _05501_ _05516_ VGND VGND VPWR VPWR _05517_ sky130_fd_sc_hd__xnor2_1
X_16032_ net2239 _08056_ net2812 VGND VGND VPWR VPWR _08099_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13175_ _05432_ _05433_ net1000 net999 VGND VGND VPWR VPWR _05448_ sky130_fd_sc_hd__or4_1
XFILLER_0_131_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4050 net4051 VGND VGND VPWR VPWR net4050 sky130_fd_sc_hd__clkbuf_1
Xwire4061 _08830_ VGND VGND VPWR VPWR net4061 sky130_fd_sc_hd__clkbuf_1
Xwire4072 net4073 VGND VGND VPWR VPWR net4072 sky130_fd_sc_hd__buf_1
XFILLER_0_102_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17983_ _09825_ net1779 VGND VGND VPWR VPWR _09834_ sky130_fd_sc_hd__nand2_1
Xwire4083 net4084 VGND VGND VPWR VPWR net4083 sky130_fd_sc_hd__buf_1
Xwire4094 _07352_ VGND VGND VPWR VPWR net4094 sky130_fd_sc_hd__buf_1
X_19722_ _11553_ net604 _11556_ net569 VGND VGND VPWR VPWR _11557_ sky130_fd_sc_hd__o22a_1
X_16934_ net6416 _08890_ _08871_ _08897_ VGND VGND VPWR VPWR _08898_ sky130_fd_sc_hd__o211a_1
Xwire3371 net3377 VGND VGND VPWR VPWR net3371 sky130_fd_sc_hd__clkbuf_1
Xwire3382 _08759_ VGND VGND VPWR VPWR net3382 sky130_fd_sc_hd__buf_1
Xwire3393 _07723_ VGND VGND VPWR VPWR net3393 sky130_fd_sc_hd__buf_1
Xwire2670 _07694_ VGND VGND VPWR VPWR net2670 sky130_fd_sc_hd__buf_1
XFILLER_0_74_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19653_ net3880 VGND VGND VPWR VPWR _11489_ sky130_fd_sc_hd__buf_1
X_16865_ net6363 net6344 net6325 net6309 net6518 net6498 VGND VGND VPWR VPWR _08830_
+ sky130_fd_sc_hd__mux4_1
Xwire2681 _07560_ VGND VGND VPWR VPWR net2681 sky130_fd_sc_hd__buf_1
X_18604_ net1070 _10451_ VGND VGND VPWR VPWR _10452_ sky130_fd_sc_hd__xnor2_1
X_15816_ _07883_ _07879_ _07880_ VGND VGND VPWR VPWR _07886_ sky130_fd_sc_hd__and3_1
X_19584_ _11353_ _11361_ VGND VGND VPWR VPWR _11421_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16796_ net9240 net7182 net3369 VGND VGND VPWR VPWR _08788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18535_ net1071 _10383_ VGND VGND VPWR VPWR _10384_ sky130_fd_sc_hd__xnor2_2
X_15747_ _07802_ _07817_ VGND VGND VPWR VPWR _07818_ sky130_fd_sc_hd__xor2_1
XFILLER_0_176_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12959_ net1003 _05231_ _05221_ VGND VGND VPWR VPWR _05232_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18466_ _10313_ _10314_ _10315_ VGND VGND VPWR VPWR _10316_ sky130_fd_sc_hd__mux2_1
X_15678_ net3395 _07746_ _07747_ net3397 _07748_ VGND VGND VPWR VPWR _07749_ sky130_fd_sc_hd__a221o_1
XFILLER_0_114_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17417_ svm0.delta\[12\] VGND VGND VPWR VPWR _09319_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14629_ net2881 _06785_ VGND VGND VPWR VPWR _06797_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18397_ _10245_ net1210 VGND VGND VPWR VPWR _10248_ sky130_fd_sc_hd__xor2_1
XFILLER_0_117_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17348_ net3278 _09212_ _09259_ _09260_ VGND VGND VPWR VPWR _09262_ sky130_fd_sc_hd__and4_1
XFILLER_0_172_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17279_ net7606 net2983 net153 net2158 net9190 VGND VGND VPWR VPWR _00373_ sky130_fd_sc_hd__a32o_1
XFILLER_0_114_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19018_ net6208 _10796_ _10798_ _10853_ _10854_ VGND VGND VPWR VPWR _10855_ sky130_fd_sc_hd__a221o_1
XFILLER_0_140_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20290_ _12095_ VGND VGND VPWR VPWR _12096_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23980_ _03839_ _03841_ VGND VGND VPWR VPWR _03844_ sky130_fd_sc_hd__nor2_1
XFILLER_0_177_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22931_ net5327 pid_d.curr_int\[13\] VGND VGND VPWR VPWR _02821_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25650_ clknet_leaf_1_clk _00523_ net8403 VGND VGND VPWR VPWR pid_d.curr_int\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_22862_ net5981 _02747_ pid_d.out\[4\] VGND VGND VPWR VPWR _02759_ sky130_fd_sc_hd__o21a_1
X_24601_ net5170 pid_q.prev_int\[14\] VGND VGND VPWR VPWR _04456_ sky130_fd_sc_hd__and2_1
XFILLER_0_196_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21813_ net5978 pid_d.prev_int\[7\] VGND VGND VPWR VPWR _01822_ sky130_fd_sc_hd__xor2_1
X_22793_ _02704_ VGND VGND VPWR VPWR _00623_ sky130_fd_sc_hd__clkbuf_1
X_25581_ clknet_leaf_86_clk _00454_ net8531 VGND VGND VPWR VPWR cordic0.cos\[1\] sky130_fd_sc_hd__dfrtp_1
X_24532_ _04330_ _04337_ net200 _04383_ net265 VGND VGND VPWR VPWR _04389_ sky130_fd_sc_hd__o221a_1
X_21744_ _01661_ _01663_ _01662_ VGND VGND VPWR VPWR _01754_ sky130_fd_sc_hd__o21a_1
XFILLER_0_182_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8305 net8306 VGND VGND VPWR VPWR net8305 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4003 _09451_ VGND VGND VPWR VPWR net4003 sky130_fd_sc_hd__buf_1
XFILLER_0_175_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8316 net8317 VGND VGND VPWR VPWR net8316 sky130_fd_sc_hd__clkbuf_1
Xwire8327 net148 VGND VGND VPWR VPWR net8327 sky130_fd_sc_hd__clkbuf_1
X_24463_ pid_q.prev_error\[12\] net5167 VGND VGND VPWR VPWR _04321_ sky130_fd_sc_hd__nand2_1
X_21675_ _01672_ _01685_ VGND VGND VPWR VPWR _01686_ sky130_fd_sc_hd__xnor2_1
Xwire7604 net7601 VGND VGND VPWR VPWR net7604 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire8349 net8352 VGND VGND VPWR VPWR net8349 sky130_fd_sc_hd__buf_1
X_23414_ net4963 net4666 VGND VGND VPWR VPWR _03284_ sky130_fd_sc_hd__nand2_1
Xwire7615 net7616 VGND VGND VPWR VPWR net7615 sky130_fd_sc_hd__clkbuf_2
X_20626_ net6173 _12400_ _12401_ VGND VGND VPWR VPWR _12406_ sky130_fd_sc_hd__o21ai_1
Xmax_length4047 net4048 VGND VGND VPWR VPWR net4047 sky130_fd_sc_hd__clkbuf_1
Xfanout6819 cordic0.vec\[1\]\[15\] VGND VGND VPWR VPWR net6819 sky130_fd_sc_hd__buf_1
XFILLER_0_191_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24394_ _04251_ _04180_ _04252_ VGND VGND VPWR VPWR _04253_ sky130_fd_sc_hd__a21o_1
Xwire7626 net7627 VGND VGND VPWR VPWR net7626 sky130_fd_sc_hd__buf_1
Xmax_length4058 _08834_ VGND VGND VPWR VPWR net4058 sky130_fd_sc_hd__buf_1
Xwire7648 net7646 VGND VGND VPWR VPWR net7648 sky130_fd_sc_hd__buf_1
XFILLER_0_11_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6903 net6901 VGND VGND VPWR VPWR net6903 sky130_fd_sc_hd__buf_1
Xmax_length2601 net2602 VGND VGND VPWR VPWR net2601 sky130_fd_sc_hd__buf_1
X_23345_ _02939_ _02944_ net2432 VGND VGND VPWR VPWR _03215_ sky130_fd_sc_hd__o21a_1
Xwire7659 svm0.periodTop\[13\] VGND VGND VPWR VPWR net7659 sky130_fd_sc_hd__clkbuf_1
X_20557_ net2082 net2084 _12329_ VGND VGND VPWR VPWR _12342_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6925 net6927 VGND VGND VPWR VPWR net6925 sky130_fd_sc_hd__buf_1
XFILLER_0_6_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2634 net2635 VGND VGND VPWR VPWR net2634 sky130_fd_sc_hd__buf_1
Xwire6958 net6959 VGND VGND VPWR VPWR net6958 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23276_ _03114_ _03128_ _03120_ VGND VGND VPWR VPWR _03146_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20488_ net6935 net6917 net6904 net6890 net6513 net6491 VGND VGND VPWR VPWR _12276_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_30_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22227_ net1704 net1703 VGND VGND VPWR VPWR _02232_ sky130_fd_sc_hd__xor2_1
X_25015_ _04768_ _04769_ VGND VGND VPWR VPWR _04770_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22158_ net2476 _02163_ VGND VGND VPWR VPWR _02164_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21109_ _01117_ _01118_ VGND VGND VPWR VPWR _01125_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_195_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22089_ _02095_ VGND VGND VPWR VPWR _02096_ sky130_fd_sc_hd__inv_2
X_14980_ net1901 _07053_ VGND VGND VPWR VPWR _07054_ sky130_fd_sc_hd__xnor2_1
Xwire1210 _10247_ VGND VGND VPWR VPWR net1210 sky130_fd_sc_hd__buf_1
Xwire1221 net1222 VGND VGND VPWR VPWR net1221 sky130_fd_sc_hd__buf_1
X_13931_ _06191_ _06196_ VGND VGND VPWR VPWR _06197_ sky130_fd_sc_hd__xnor2_1
X_25917_ clknet_leaf_28_clk _00790_ net8657 VGND VGND VPWR VPWR pid_q.out\[13\] sky130_fd_sc_hd__dfrtp_1
Xwire1232 net1233 VGND VGND VPWR VPWR net1232 sky130_fd_sc_hd__buf_1
Xwire1243 _08578_ VGND VGND VPWR VPWR net1243 sky130_fd_sc_hd__buf_1
Xwire1254 net1255 VGND VGND VPWR VPWR net1254 sky130_fd_sc_hd__buf_1
XFILLER_0_156_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1265 _07807_ VGND VGND VPWR VPWR net1265 sky130_fd_sc_hd__buf_1
Xwire1276 _07294_ VGND VGND VPWR VPWR net1276 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_88_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16650_ matmul0.matmul_stage_inst.mult1\[4\] VGND VGND VPWR VPWR _08686_ sky130_fd_sc_hd__inv_2
X_13862_ net7767 net1579 VGND VGND VPWR VPWR _06129_ sky130_fd_sc_hd__and2_1
X_25848_ clknet_leaf_20_clk _00721_ net8615 VGND VGND VPWR VPWR pid_q.mult0.b\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1287 _07054_ VGND VGND VPWR VPWR net1287 sky130_fd_sc_hd__buf_1
XFILLER_0_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15601_ _07671_ _07672_ VGND VGND VPWR VPWR _07673_ sky130_fd_sc_hd__xnor2_1
X_12813_ _04955_ _04941_ net1343 _04969_ VGND VGND VPWR VPWR _05086_ sky130_fd_sc_hd__a31o_1
XFILLER_0_158_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16581_ matmul0.matmul_stage_inst.mult2\[1\] net440 net2620 VGND VGND VPWR VPWR _08638_
+ sky130_fd_sc_hd__mux2_1
X_13793_ net1563 net1148 net7615 VGND VGND VPWR VPWR _06061_ sky130_fd_sc_hd__nand3b_1
X_25779_ clknet_leaf_81_clk _00652_ net8500 VGND VGND VPWR VPWR matmul0.beta_pass\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_18320_ net6852 _10170_ VGND VGND VPWR VPWR _10171_ sky130_fd_sc_hd__xnor2_4
X_15532_ net3597 net3591 net4092 net4089 VGND VGND VPWR VPWR _07605_ sky130_fd_sc_hd__o22a_1
XFILLER_0_84_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12744_ _05013_ _05016_ VGND VGND VPWR VPWR _05017_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout8722 net8732 VGND VGND VPWR VPWR net8722 sky130_fd_sc_hd__buf_1
XFILLER_0_195_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18251_ net6857 net6811 VGND VGND VPWR VPWR _10102_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_167_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15463_ _07390_ _07535_ _07536_ VGND VGND VPWR VPWR _07537_ sky130_fd_sc_hd__a21o_1
X_12675_ _04946_ _04947_ VGND VGND VPWR VPWR _04948_ sky130_fd_sc_hd__xnor2_1
X_17202_ _09148_ _09151_ VGND VGND VPWR VPWR _09152_ sky130_fd_sc_hd__nand2_1
X_14414_ _06614_ matmul0.b_in\[5\] _06606_ VGND VGND VPWR VPWR _06615_ sky130_fd_sc_hd__mux2_1
Xwire8850 net8851 VGND VGND VPWR VPWR net8850 sky130_fd_sc_hd__clkbuf_1
X_18182_ _10031_ _10032_ _10030_ VGND VGND VPWR VPWR _10033_ sky130_fd_sc_hd__o21a_1
Xwire8861 net147 VGND VGND VPWR VPWR net8861 sky130_fd_sc_hd__clkbuf_1
X_15394_ net829 _07334_ VGND VGND VPWR VPWR _07468_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8872 net8869 VGND VGND VPWR VPWR net8872 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8883 net8884 VGND VGND VPWR VPWR net8883 sky130_fd_sc_hd__clkbuf_1
X_17133_ _09075_ _09077_ _09087_ VGND VGND VPWR VPWR _09088_ sky130_fd_sc_hd__o21a_1
Xwire540 net541 VGND VGND VPWR VPWR net540 sky130_fd_sc_hd__buf_1
Xwire8894 net8890 VGND VGND VPWR VPWR net8894 sky130_fd_sc_hd__buf_1
X_14345_ net7299 net1301 net2898 net5361 _06560_ VGND VGND VPWR VPWR _06561_ sky130_fd_sc_hd__a221o_1
Xwire551 _02339_ VGND VGND VPWR VPWR net551 sky130_fd_sc_hd__buf_1
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire562 net563 VGND VGND VPWR VPWR net562 sky130_fd_sc_hd__clkbuf_1
Xwire573 _08093_ VGND VGND VPWR VPWR net573 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire584 net585 VGND VGND VPWR VPWR net584 sky130_fd_sc_hd__clkbuf_1
X_17064_ net4246 VGND VGND VPWR VPWR _09023_ sky130_fd_sc_hd__buf_1
X_14276_ net52 net2903 net2266 net7973 VGND VGND VPWR VPWR _00047_ sky130_fd_sc_hd__a22o_1
Xwire595 net596 VGND VGND VPWR VPWR net595 sky130_fd_sc_hd__buf_1
XFILLER_0_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16015_ _08081_ _08082_ VGND VGND VPWR VPWR _08083_ sky130_fd_sc_hd__nand2_1
X_13227_ net1135 _05499_ VGND VGND VPWR VPWR _05500_ sky130_fd_sc_hd__xor2_1
XFILLER_0_21_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13158_ net918 _05430_ VGND VGND VPWR VPWR _05431_ sky130_fd_sc_hd__xnor2_1
X_13089_ _05262_ _05277_ VGND VGND VPWR VPWR _05362_ sky130_fd_sc_hd__or2_1
X_17966_ _09807_ _09816_ VGND VGND VPWR VPWR _09817_ sky130_fd_sc_hd__xnor2_1
Xwire3190 _10938_ VGND VGND VPWR VPWR net3190 sky130_fd_sc_hd__clkbuf_2
X_16917_ net6369 _08879_ VGND VGND VPWR VPWR _08881_ sky130_fd_sc_hd__nand2_1
X_19705_ _11534_ net1057 VGND VGND VPWR VPWR _11541_ sky130_fd_sc_hd__xor2_1
XFILLER_0_100_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17897_ net3348 net3969 net3995 VGND VGND VPWR VPWR _09748_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19636_ _11348_ _11411_ VGND VGND VPWR VPWR _11473_ sky130_fd_sc_hd__or2_1
X_16848_ cordic0.sin\[12\] matmul0.sin\[12\] net4287 VGND VGND VPWR VPWR _08815_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_195_Right_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19567_ net1417 _11403_ VGND VGND VPWR VPWR _11404_ sky130_fd_sc_hd__xnor2_1
X_16779_ net7598 matmul0.a\[9\] net3379 VGND VGND VPWR VPWR _08779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18518_ net3310 net3989 _10063_ net6872 VGND VGND VPWR VPWR _10367_ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19498_ net6182 net6205 _11333_ _11334_ VGND VGND VPWR VPWR _11335_ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18449_ net6998 _10294_ _10296_ _10297_ _10298_ VGND VGND VPWR VPWR _10299_ sky130_fd_sc_hd__o221a_1
XFILLER_0_75_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21460_ _01360_ _01362_ _01361_ VGND VGND VPWR VPWR _01473_ sky130_fd_sc_hd__o21a_1
X_20411_ _12206_ _12207_ _12182_ net603 VGND VGND VPWR VPWR _12208_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_43_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21391_ net5462 VGND VGND VPWR VPWR _01405_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5509 net5510 VGND VGND VPWR VPWR net5509 sky130_fd_sc_hd__buf_1
Xclkbuf_4_6__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_4_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_23130_ net5143 net4631 _02998_ _02999_ VGND VGND VPWR VPWR _03000_ sky130_fd_sc_hd__a31o_1
X_20342_ _12141_ _12143_ _12144_ net9218 VGND VGND VPWR VPWR _00487_ sky130_fd_sc_hd__a22o_1
Xwire4808 net4809 VGND VGND VPWR VPWR net4808 sky130_fd_sc_hd__buf_1
Xwire4819 net4820 VGND VGND VPWR VPWR net4819 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23061_ _02894_ _02905_ _02906_ VGND VGND VPWR VPWR _02931_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_141_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20273_ net8122 cordic0.domain\[0\] net2533 VGND VGND VPWR VPWR _12082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22012_ _02016_ _01919_ _02018_ VGND VGND VPWR VPWR _02019_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_179_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23963_ _03824_ _03826_ VGND VGND VPWR VPWR _03827_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_166_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_95_clk clknet_4_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_95_clk sky130_fd_sc_hd__clkbuf_16
X_25702_ clknet_leaf_2_clk _00575_ net8572 VGND VGND VPWR VPWR pid_d.mult0.b\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_22914_ net4333 _02804_ _02805_ net298 net4362 VGND VGND VPWR VPWR _02806_ sky130_fd_sc_hd__a32o_1
X_23894_ _03757_ _03679_ _03680_ VGND VGND VPWR VPWR _03759_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_162_Right_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25633_ clknet_leaf_105_clk _00506_ net8356 VGND VGND VPWR VPWR cordic0.vec\[0\]\[5\]
+ sky130_fd_sc_hd__dfstp_1
X_22845_ net5982 VGND VGND VPWR VPWR _02744_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25564_ clknet_leaf_66_clk _00437_ net8659 VGND VGND VPWR VPWR state\[2\] sky130_fd_sc_hd__dfrtp_1
X_22776_ pid_d.kp\[0\] _02653_ net1679 VGND VGND VPWR VPWR _02696_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8102 net88 VGND VGND VPWR VPWR net8102 sky130_fd_sc_hd__clkbuf_1
X_24515_ _04366_ _04371_ VGND VGND VPWR VPWR _04372_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_94_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21727_ _01736_ _01646_ pid_d.curr_int\[5\] VGND VGND VPWR VPWR _01737_ sky130_fd_sc_hd__o21ba_1
Xwire8113 net8114 VGND VGND VPWR VPWR net8113 sky130_fd_sc_hd__clkbuf_1
X_25495_ clknet_leaf_48_clk _00375_ net8759 VGND VGND VPWR VPWR svm0.rising sky130_fd_sc_hd__dfstp_1
XFILLER_0_54_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8124 net8125 VGND VGND VPWR VPWR net8124 sky130_fd_sc_hd__clkbuf_1
Xwire8135 net46 VGND VGND VPWR VPWR net8135 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7401 net7402 VGND VGND VPWR VPWR net7401 sky130_fd_sc_hd__clkbuf_1
Xwire8146 net8147 VGND VGND VPWR VPWR net8146 sky130_fd_sc_hd__clkbuf_1
X_24446_ _04302_ _04303_ VGND VGND VPWR VPWR _04304_ sky130_fd_sc_hd__or2_1
X_21658_ _01667_ _01668_ VGND VGND VPWR VPWR _01669_ sky130_fd_sc_hd__xor2_1
Xwire8157 net8158 VGND VGND VPWR VPWR net8157 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7412 matmul0.matmul_stage_inst.c\[6\] VGND VGND VPWR VPWR net7412 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7423 matmul0.matmul_stage_inst.b\[8\] VGND VGND VPWR VPWR net7423 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8168 net8169 VGND VGND VPWR VPWR net8168 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3121 _00872_ VGND VGND VPWR VPWR net3121 sky130_fd_sc_hd__buf_1
Xwire8179 net38 VGND VGND VPWR VPWR net8179 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7434 net7435 VGND VGND VPWR VPWR net7434 sky130_fd_sc_hd__clkbuf_1
Xfanout6638 net6641 VGND VGND VPWR VPWR net6638 sky130_fd_sc_hd__buf_1
XFILLER_0_136_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20609_ net1740 _12385_ _12387_ _12389_ net6216 VGND VGND VPWR VPWR _12390_ sky130_fd_sc_hd__o32a_1
Xmax_length3143 net3144 VGND VGND VPWR VPWR net3143 sky130_fd_sc_hd__buf_1
Xwire7456 net7457 VGND VGND VPWR VPWR net7456 sky130_fd_sc_hd__buf_1
Xwire6722 net6723 VGND VGND VPWR VPWR net6722 sky130_fd_sc_hd__buf_1
Xwire7467 net7466 VGND VGND VPWR VPWR net7467 sky130_fd_sc_hd__buf_1
X_24377_ _04229_ _04235_ VGND VGND VPWR VPWR _04236_ sky130_fd_sc_hd__xnor2_1
X_21589_ _01595_ _01600_ VGND VGND VPWR VPWR _01601_ sky130_fd_sc_hd__xnor2_2
Xwire6733 net6734 VGND VGND VPWR VPWR net6733 sky130_fd_sc_hd__buf_1
X_14130_ _06384_ _06391_ VGND VGND VPWR VPWR _06392_ sky130_fd_sc_hd__xor2_1
Xfanout5948 net5955 VGND VGND VPWR VPWR net5948 sky130_fd_sc_hd__clkbuf_1
X_23328_ _02925_ _03197_ _02922_ net3751 VGND VGND VPWR VPWR _03198_ sky130_fd_sc_hd__or4b_1
XFILLER_0_104_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length3198 _10911_ VGND VGND VPWR VPWR net3198 sky130_fd_sc_hd__buf_1
Xwire6766 net6767 VGND VGND VPWR VPWR net6766 sky130_fd_sc_hd__buf_1
XFILLER_0_34_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2464 net2465 VGND VGND VPWR VPWR net2464 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14061_ _06307_ _06305_ net1561 VGND VGND VPWR VPWR _06324_ sky130_fd_sc_hd__a21bo_1
Xwire6799 net6801 VGND VGND VPWR VPWR net6799 sky130_fd_sc_hd__buf_1
X_23259_ _03120_ _03128_ VGND VGND VPWR VPWR _03129_ sky130_fd_sc_hd__xnor2_1
X_13012_ net3693 VGND VGND VPWR VPWR _05285_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_20_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17820_ _09666_ _09669_ VGND VGND VPWR VPWR _09671_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17751_ net6908 net6948 VGND VGND VPWR VPWR _09602_ sky130_fd_sc_hd__xor2_4
Xhold6 matmul0.matmul_stage_inst.a\[2\] VGND VGND VPWR VPWR net8959 sky130_fd_sc_hd__dlygate4sd3_1
X_14963_ net6612 net7432 matmul0.matmul_stage_inst.a\[2\] net6583 VGND VGND VPWR VPWR
+ _07037_ sky130_fd_sc_hd__a22o_1
Xwire1040 _02053_ VGND VGND VPWR VPWR net1040 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_86_clk clknet_4_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_86_clk sky130_fd_sc_hd__clkbuf_16
Xwire1051 _01013_ VGND VGND VPWR VPWR net1051 sky130_fd_sc_hd__buf_1
X_16702_ matmul0.matmul_stage_inst.mult2\[12\] matmul0.matmul_stage_inst.mult1\[12\]
+ VGND VGND VPWR VPWR _08731_ sky130_fd_sc_hd__xor2_1
X_13914_ _06117_ net1311 _06179_ net4248 VGND VGND VPWR VPWR _06180_ sky130_fd_sc_hd__o22a_1
Xwire1062 net1063 VGND VGND VPWR VPWR net1062 sky130_fd_sc_hd__clkbuf_1
X_17682_ svm0.tA\[15\] _09520_ net4030 VGND VGND VPWR VPWR _09562_ sky130_fd_sc_hd__a21o_1
Xwire1073 _10184_ VGND VGND VPWR VPWR net1073 sky130_fd_sc_hd__dlymetal6s2s_1
X_14894_ net3602 net3601 VGND VGND VPWR VPWR _06968_ sky130_fd_sc_hd__nor2_1
Xwire1084 net1085 VGND VGND VPWR VPWR net1084 sky130_fd_sc_hd__buf_1
XFILLER_0_18_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19421_ _11255_ _11256_ _11257_ VGND VGND VPWR VPWR _11258_ sky130_fd_sc_hd__a21o_1
Xwire1095 net1096 VGND VGND VPWR VPWR net1095 sky130_fd_sc_hd__clkbuf_1
X_16633_ matmul0.matmul_stage_inst.mult1\[2\] VGND VGND VPWR VPWR _08671_ sky130_fd_sc_hd__inv_2
X_13845_ _06105_ _06111_ VGND VGND VPWR VPWR _06112_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_162_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19352_ net6295 _11147_ _10991_ VGND VGND VPWR VPWR _11189_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16564_ _08582_ _08585_ _08581_ VGND VGND VPWR VPWR _08623_ sky130_fd_sc_hd__a21oi_1
X_13776_ _05965_ _05966_ _05968_ _05969_ VGND VGND VPWR VPWR _06044_ sky130_fd_sc_hd__o22a_1
X_18303_ net6774 net3926 VGND VGND VPWR VPWR _10154_ sky130_fd_sc_hd__nand2_1
XFILLER_0_174_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15515_ _07478_ _07494_ _07492_ VGND VGND VPWR VPWR _07588_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_73_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12727_ _04994_ _04997_ net1611 _04979_ VGND VGND VPWR VPWR _05000_ sky130_fd_sc_hd__a211o_1
X_19283_ net6323 net6335 VGND VGND VPWR VPWR _11120_ sky130_fd_sc_hd__or2b_1
Xfanout8530 net8546 VGND VGND VPWR VPWR net8530 sky130_fd_sc_hd__buf_1
X_16495_ net2634 net2628 VGND VGND VPWR VPWR _08555_ sky130_fd_sc_hd__nor2_2
X_18234_ _10083_ _10084_ _09810_ VGND VGND VPWR VPWR _10085_ sky130_fd_sc_hd__a21boi_1
X_15446_ _07518_ _07519_ VGND VGND VPWR VPWR _07520_ sky130_fd_sc_hd__xnor2_1
Xfanout8585 net8593 VGND VGND VPWR VPWR net8585 sky130_fd_sc_hd__clkbuf_1
X_12658_ net7364 _04892_ net4278 net2990 svm0.vC\[0\] VGND VGND VPWR VPWR _04931_
+ sky130_fd_sc_hd__a32oi_1
Xfanout7851 net7856 VGND VGND VPWR VPWR net7851 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout7873 net7885 VGND VGND VPWR VPWR net7873 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18165_ _10006_ _10014_ _10015_ _10012_ VGND VGND VPWR VPWR _10016_ sky130_fd_sc_hd__o211a_1
XFILLER_0_170_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8691 net8687 VGND VGND VPWR VPWR net8691 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_111_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15377_ net2811 net2249 _07450_ VGND VGND VPWR VPWR _07451_ sky130_fd_sc_hd__and3_1
X_12589_ net4365 VGND VGND VPWR VPWR _04872_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_10_clk clknet_4_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_128_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17116_ net5990 net2170 _09071_ VGND VGND VPWR VPWR _09072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire370 net371 VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14328_ net8262 net3642 VGND VGND VPWR VPWR _06548_ sky130_fd_sc_hd__and2_1
Xwire7990 net7991 VGND VGND VPWR VPWR net7990 sky130_fd_sc_hd__clkbuf_2
Xwire381 _02272_ VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__buf_1
XFILLER_0_29_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18096_ _09901_ _09942_ _09946_ VGND VGND VPWR VPWR _09947_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_111_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire392 net393 VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17047_ _09005_ VGND VGND VPWR VPWR _09006_ sky130_fd_sc_hd__buf_1
X_14259_ net6455 net6445 VGND VGND VPWR VPWR _06513_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_14__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_4_14__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_18998_ _10817_ _10834_ VGND VGND VPWR VPWR _10835_ sky130_fd_sc_hd__nand2_1
XFILLER_0_174_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17949_ net7115 net7124 VGND VGND VPWR VPWR _09800_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_77_clk clknet_4_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_77_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_75_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20960_ _00954_ _00975_ VGND VGND VPWR VPWR _00976_ sky130_fd_sc_hd__xnor2_1
Xmax_length7409 matmul0.matmul_stage_inst.c\[9\] VGND VGND VPWR VPWR net7409 sky130_fd_sc_hd__clkbuf_1
X_19619_ _11382_ net3907 _11272_ _11455_ VGND VGND VPWR VPWR _11456_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_45_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20891_ net5579 net5822 VGND VGND VPWR VPWR _00907_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22630_ net9061 _02544_ net2042 _02598_ VGND VGND VPWR VPWR _00566_ sky130_fd_sc_hd__a22o_1
X_22561_ net6754 net6603 net4347 VGND VGND VPWR VPWR _02545_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24300_ _04153_ _04159_ VGND VGND VPWR VPWR _04160_ sky130_fd_sc_hd__xnor2_2
X_21512_ _01524_ VGND VGND VPWR VPWR _01525_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22492_ _02490_ _02492_ VGND VGND VPWR VPWR _02493_ sky130_fd_sc_hd__xnor2_1
X_25280_ clknet_leaf_92_clk _00163_ net8434 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.c\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24231_ net4802 _03981_ _04090_ VGND VGND VPWR VPWR _04092_ sky130_fd_sc_hd__a21oi_1
X_21443_ net5705 net5582 VGND VGND VPWR VPWR _01456_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24162_ _03869_ _03937_ VGND VGND VPWR VPWR _04024_ sky130_fd_sc_hd__nand2_1
Xwire5306 matmul0.beta_pass\[1\] VGND VGND VPWR VPWR net5306 sky130_fd_sc_hd__buf_1
Xwire5317 net5318 VGND VGND VPWR VPWR net5317 sky130_fd_sc_hd__clkbuf_1
X_21374_ _01284_ _01286_ _01387_ VGND VGND VPWR VPWR _01388_ sky130_fd_sc_hd__o21ai_1
Xwire5328 net5329 VGND VGND VPWR VPWR net5328 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23113_ _02973_ _02978_ _02982_ VGND VGND VPWR VPWR _02983_ sky130_fd_sc_hd__a21o_1
Xwire4605 net4606 VGND VGND VPWR VPWR net4605 sky130_fd_sc_hd__buf_1
XFILLER_0_160_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20325_ net2182 _12128_ net4241 VGND VGND VPWR VPWR _12129_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4616 net4617 VGND VGND VPWR VPWR net4616 sky130_fd_sc_hd__buf_1
X_24093_ net5178 VGND VGND VPWR VPWR _03955_ sky130_fd_sc_hd__inv_2
Xwire4627 net4628 VGND VGND VPWR VPWR net4627 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4638 net4630 VGND VGND VPWR VPWR net4638 sky130_fd_sc_hd__buf_1
Xwire4649 net4650 VGND VGND VPWR VPWR net4649 sky130_fd_sc_hd__clkbuf_1
Xwire3904 net3905 VGND VGND VPWR VPWR net3904 sky130_fd_sc_hd__clkbuf_1
X_23044_ _02882_ _02883_ VGND VGND VPWR VPWR _02914_ sky130_fd_sc_hd__xnor2_1
Xwire3915 net3916 VGND VGND VPWR VPWR net3915 sky130_fd_sc_hd__buf_1
X_20256_ net15 net16 _12061_ net8121 VGND VGND VPWR VPWR _12069_ sky130_fd_sc_hd__a31o_1
Xwire3926 _10123_ VGND VGND VPWR VPWR net3926 sky130_fd_sc_hd__buf_1
Xwire3937 net3939 VGND VGND VPWR VPWR net3937 sky130_fd_sc_hd__clkbuf_1
Xwire3948 net3951 VGND VGND VPWR VPWR net3948 sky130_fd_sc_hd__buf_1
Xwire3959 net3960 VGND VGND VPWR VPWR net3959 sky130_fd_sc_hd__buf_1
XFILLER_0_177_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20187_ net952 net867 VGND VGND VPWR VPWR _12013_ sky130_fd_sc_hd__xor2_1
X_24995_ net7483 net3270 net8874 VGND VGND VPWR VPWR _04753_ sky130_fd_sc_hd__nor3b_1
Xclkbuf_leaf_68_clk clknet_4_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_16
X_23946_ _03808_ _03809_ VGND VGND VPWR VPWR _03810_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_192_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length8644 net8633 VGND VGND VPWR VPWR net8644 sky130_fd_sc_hd__buf_1
XFILLER_0_193_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length8666 net8667 VGND VGND VPWR VPWR net8666 sky130_fd_sc_hd__buf_1
X_23877_ net4729 net3747 _03738_ VGND VGND VPWR VPWR _03742_ sky130_fd_sc_hd__or3_1
Xmax_length8699 net8700 VGND VGND VPWR VPWR net8699 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13630_ _05896_ _05899_ VGND VGND VPWR VPWR _05900_ sky130_fd_sc_hd__xnor2_2
X_25616_ clknet_leaf_109_clk _00489_ net8346 VGND VGND VPWR VPWR cordic0.slte0.opA\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_22828_ _02727_ _02728_ VGND VGND VPWR VPWR _02729_ sky130_fd_sc_hd__nand2_1
X_13561_ _05830_ _05831_ VGND VGND VPWR VPWR _05832_ sky130_fd_sc_hd__or2b_1
X_25547_ clknet_leaf_28_clk _00427_ net8649 VGND VGND VPWR VPWR pid_q.prev_int\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22759_ net4302 net8086 VGND VGND VPWR VPWR _02684_ sky130_fd_sc_hd__and2_1
Xfanout7103 net7109 VGND VGND VPWR VPWR net7103 sky130_fd_sc_hd__buf_1
Xfanout7114 cordic0.vec\[1\]\[2\] VGND VGND VPWR VPWR net7114 sky130_fd_sc_hd__buf_1
X_15300_ net4207 net4201 net4216 net4214 VGND VGND VPWR VPWR _07374_ sky130_fd_sc_hd__o22a_1
XFILLER_0_137_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout7125 cordic0.vec\[1\]\[1\] VGND VGND VPWR VPWR net7125 sky130_fd_sc_hd__buf_1
XFILLER_0_66_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16280_ net2682 _08342_ _08343_ VGND VGND VPWR VPWR _08344_ sky130_fd_sc_hd__a21o_1
X_25478_ clknet_leaf_46_clk _00358_ net8787 VGND VGND VPWR VPWR svm0.tA\[0\] sky130_fd_sc_hd__dfrtp_1
X_13492_ net7947 net1130 net1564 VGND VGND VPWR VPWR _05765_ sky130_fd_sc_hd__and3_1
XFILLER_0_164_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire7220 net7221 VGND VGND VPWR VPWR net7220 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7231 net7236 VGND VGND VPWR VPWR net7231 sky130_fd_sc_hd__clkbuf_1
X_15231_ _07304_ VGND VGND VPWR VPWR _07305_ sky130_fd_sc_hd__clkbuf_1
X_24429_ net4872 net4504 VGND VGND VPWR VPWR _04287_ sky130_fd_sc_hd__nand2_1
Xwire7242 net7243 VGND VGND VPWR VPWR net7242 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5701 net5716 VGND VGND VPWR VPWR net5701 sky130_fd_sc_hd__buf_1
Xfanout5712 pid_d.mult0.b\[12\] VGND VGND VPWR VPWR net5712 sky130_fd_sc_hd__buf_1
Xwire7253 net7254 VGND VGND VPWR VPWR net7253 sky130_fd_sc_hd__clkbuf_1
Xfanout6457 net6463 VGND VGND VPWR VPWR net6457 sky130_fd_sc_hd__buf_1
Xwire7264 net7270 VGND VGND VPWR VPWR net7264 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_151_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7275 net7276 VGND VGND VPWR VPWR net7275 sky130_fd_sc_hd__clkbuf_1
Xfanout6479 net6482 VGND VGND VPWR VPWR net6479 sky130_fd_sc_hd__buf_1
Xwire6530 cordic0.gm0.iter\[0\] VGND VGND VPWR VPWR net6530 sky130_fd_sc_hd__buf_1
XFILLER_0_34_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15162_ _07223_ net1884 VGND VGND VPWR VPWR _07236_ sky130_fd_sc_hd__xnor2_1
Xwire6541 net6539 VGND VGND VPWR VPWR net6541 sky130_fd_sc_hd__buf_1
Xwire7286 matmul0.alpha_pass\[7\] VGND VGND VPWR VPWR net7286 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6552 net6547 VGND VGND VPWR VPWR net6552 sky130_fd_sc_hd__buf_1
Xwire7297 net7298 VGND VGND VPWR VPWR net7297 sky130_fd_sc_hd__clkbuf_1
Xwire6563 net6564 VGND VGND VPWR VPWR net6563 sky130_fd_sc_hd__buf_1
X_14113_ net7680 _06374_ VGND VGND VPWR VPWR _06375_ sky130_fd_sc_hd__nand2_1
Xwire6585 net6584 VGND VGND VPWR VPWR net6585 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_120_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5851 net5852 VGND VGND VPWR VPWR net5851 sky130_fd_sc_hd__buf_1
X_19970_ _11799_ _11800_ VGND VGND VPWR VPWR _11801_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15093_ net1285 net1283 VGND VGND VPWR VPWR _07167_ sky130_fd_sc_hd__xnor2_1
Xmax_length2283 net2284 VGND VGND VPWR VPWR net2283 sky130_fd_sc_hd__clkbuf_1
Xwire6596 net6591 VGND VGND VPWR VPWR net6596 sky130_fd_sc_hd__clkbuf_1
Xwire5862 net5863 VGND VGND VPWR VPWR net5862 sky130_fd_sc_hd__buf_1
X_14044_ net1561 _06307_ VGND VGND VPWR VPWR _06308_ sky130_fd_sc_hd__xor2_1
X_18921_ _10716_ _10738_ net6777 VGND VGND VPWR VPWR _10761_ sky130_fd_sc_hd__a21o_1
Xwire5884 net5883 VGND VGND VPWR VPWR net5884 sky130_fd_sc_hd__buf_1
XFILLER_0_24_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18852_ net6376 _10694_ VGND VGND VPWR VPWR _10695_ sky130_fd_sc_hd__nand2_1
X_17803_ net7061 net3262 _09613_ VGND VGND VPWR VPWR _09654_ sky130_fd_sc_hd__and3_1
X_18783_ _10572_ _10593_ _10626_ VGND VGND VPWR VPWR _10627_ sky130_fd_sc_hd__o21a_1
X_15995_ _08061_ _08062_ VGND VGND VPWR VPWR _08063_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_59_clk clknet_4_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_16
X_17734_ net6509 net6457 _08943_ net3668 VGND VGND VPWR VPWR _09590_ sky130_fd_sc_hd__a31o_1
X_14946_ net6537 matmul0.matmul_stage_inst.c\[3\] matmul0.matmul_stage_inst.b\[3\]
+ net6617 VGND VGND VPWR VPWR _07020_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_192_Left_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17665_ svm0.tA\[0\] VGND VGND VPWR VPWR _09545_ sky130_fd_sc_hd__inv_2
X_14877_ _06956_ VGND VGND VPWR VPWR _00209_ sky130_fd_sc_hd__clkbuf_1
X_19404_ _11070_ _11093_ VGND VGND VPWR VPWR _11241_ sky130_fd_sc_hd__and2b_1
X_16616_ matmul0.matmul_stage_inst.mult2\[15\] net161 net3467 VGND VGND VPWR VPWR
+ _08658_ sky130_fd_sc_hd__mux2_1
X_13828_ _06093_ _06094_ VGND VGND VPWR VPWR _06095_ sky130_fd_sc_hd__xor2_1
X_17596_ net6721 svm0.tB\[6\] VGND VGND VPWR VPWR _09477_ sky130_fd_sc_hd__and2b_1
XFILLER_0_15_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19335_ _11169_ _10901_ _11170_ _10900_ _11171_ _11158_ VGND VGND VPWR VPWR _11172_
+ sky130_fd_sc_hd__mux4_1
X_16547_ net2628 _08605_ net2621 net2208 VGND VGND VPWR VPWR _08606_ sky130_fd_sc_hd__o211a_1
X_13759_ net2300 net2296 net7768 VGND VGND VPWR VPWR _06027_ sky130_fd_sc_hd__or3b_1
XFILLER_0_72_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19266_ _11099_ _11102_ VGND VGND VPWR VPWR _11103_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16478_ _08538_ VGND VGND VPWR VPWR _08539_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18217_ net3947 _10066_ _10064_ VGND VGND VPWR VPWR _10068_ sky130_fd_sc_hd__nor3_1
XFILLER_0_142_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15429_ _07398_ _07400_ _07387_ VGND VGND VPWR VPWR _07503_ sky130_fd_sc_hd__o21a_1
XFILLER_0_54_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout7670 svm0.periodTop\[12\] VGND VGND VPWR VPWR net7670 sky130_fd_sc_hd__buf_1
X_19197_ net3183 _11028_ VGND VGND VPWR VPWR _11034_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18148_ _09998_ _09957_ VGND VGND VPWR VPWR _09999_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold203 pid_d.mult0.b\[11\] VGND VGND VPWR VPWR net9156 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold214 svm0.tB\[3\] VGND VGND VPWR VPWR net9167 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold225 pid_q.prev_error\[2\] VGND VGND VPWR VPWR net9178 sky130_fd_sc_hd__dlygate4sd3_1
X_18079_ _09914_ _09923_ _09929_ VGND VGND VPWR VPWR _09930_ sky130_fd_sc_hd__nand3_1
Xhold236 pid_q.prev_int\[14\] VGND VGND VPWR VPWR net9189 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold247 pid_q.prev_int\[8\] VGND VGND VPWR VPWR net9200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 pid_q.prev_int\[6\] VGND VGND VPWR VPWR net9211 sky130_fd_sc_hd__dlygate4sd3_1
X_20110_ net6063 net6005 VGND VGND VPWR VPWR _11938_ sky130_fd_sc_hd__xor2_1
Xhold269 svm0.tC\[11\] VGND VGND VPWR VPWR net9222 sky130_fd_sc_hd__dlygate4sd3_1
X_21090_ net5581 _01054_ _01105_ net3805 VGND VGND VPWR VPWR _01106_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_13_Left_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20041_ net2581 net2498 VGND VGND VPWR VPWR _11871_ sky130_fd_sc_hd__nor2_1
Xwire1809 _08918_ VGND VGND VPWR VPWR net1809 sky130_fd_sc_hd__buf_1
XFILLER_0_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23800_ _03664_ _03665_ VGND VGND VPWR VPWR _03666_ sky130_fd_sc_hd__nand2_1
X_24780_ net7980 _04598_ _04606_ net2385 VGND VGND VPWR VPWR _04607_ sky130_fd_sc_hd__a2bb2o_1
X_21992_ _01893_ _01897_ _01744_ VGND VGND VPWR VPWR _02000_ sky130_fd_sc_hd__o21ai_1
X_23731_ _03526_ _03528_ _03596_ VGND VGND VPWR VPWR _03597_ sky130_fd_sc_hd__a21oi_2
X_20943_ net5613 net5759 VGND VGND VPWR VPWR _00959_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23662_ _03527_ _03528_ VGND VGND VPWR VPWR _03529_ sky130_fd_sc_hd__xnor2_1
Xmax_length6527 net6524 VGND VGND VPWR VPWR net6527 sky130_fd_sc_hd__clkbuf_1
X_20874_ _00878_ _00887_ _00889_ VGND VGND VPWR VPWR _00890_ sky130_fd_sc_hd__o21bai_1
X_25401_ clknet_leaf_68_clk _00284_ net8450 VGND VGND VPWR VPWR matmul0.a\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22613_ net7250 net7237 _02576_ net7227 VGND VGND VPWR VPWR _02585_ sky130_fd_sc_hd__o31a_1
X_23593_ _03453_ _03460_ VGND VGND VPWR VPWR _03461_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_165_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25332_ clknet_leaf_82_clk _00215_ net8503 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.mult1\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_22544_ net9105 net1701 _02534_ VGND VGND VPWR VPWR _00544_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25263_ clknet_leaf_77_clk _00146_ net8437 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.b\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22475_ net3778 _02474_ _02475_ VGND VGND VPWR VPWR _02476_ sky130_fd_sc_hd__or3_1
X_24214_ _03975_ VGND VGND VPWR VPWR _04075_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21426_ pid_d.curr_int\[3\] pid_d.prev_int\[3\] VGND VGND VPWR VPWR _01439_ sky130_fd_sc_hd__xnor2_1
X_25194_ clknet_leaf_63_clk _00083_ net8665 VGND VGND VPWR VPWR matmul0.b_in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire5114 net5115 VGND VGND VPWR VPWR net5114 sky130_fd_sc_hd__clkbuf_1
Xfanout4318 net4323 VGND VGND VPWR VPWR net4318 sky130_fd_sc_hd__buf_1
Xwire5125 net5126 VGND VGND VPWR VPWR net5125 sky130_fd_sc_hd__clkbuf_1
Xwire5136 net5137 VGND VGND VPWR VPWR net5136 sky130_fd_sc_hd__clkbuf_1
Xwire5147 net5148 VGND VGND VPWR VPWR net5147 sky130_fd_sc_hd__clkbuf_1
X_24145_ net4651 VGND VGND VPWR VPWR _04007_ sky130_fd_sc_hd__inv_2
Xwire4402 net4403 VGND VGND VPWR VPWR net4402 sky130_fd_sc_hd__clkbuf_1
X_21357_ _01359_ _01370_ VGND VGND VPWR VPWR _01371_ sky130_fd_sc_hd__xor2_1
Xwire4413 net4414 VGND VGND VPWR VPWR net4413 sky130_fd_sc_hd__clkbuf_1
Xwire5158 net5159 VGND VGND VPWR VPWR net5158 sky130_fd_sc_hd__buf_1
Xwire5169 pid_q.curr_int\[15\] VGND VGND VPWR VPWR net5169 sky130_fd_sc_hd__clkbuf_2
X_20308_ _12089_ _12100_ cordic0.slte0.opA\[1\] VGND VGND VPWR VPWR _12113_ sky130_fd_sc_hd__o21bai_1
Xwire3701 _04882_ VGND VGND VPWR VPWR net3701 sky130_fd_sc_hd__buf_1
Xwire4446 net4447 VGND VGND VPWR VPWR net4446 sky130_fd_sc_hd__clkbuf_1
Xwire3712 net3713 VGND VGND VPWR VPWR net3712 sky130_fd_sc_hd__clkbuf_1
X_24076_ _03869_ _03938_ VGND VGND VPWR VPWR _03939_ sky130_fd_sc_hd__xnor2_1
X_21288_ net1737 net1736 _00834_ VGND VGND VPWR VPWR _01303_ sky130_fd_sc_hd__a21bo_1
Xwire3723 net3724 VGND VGND VPWR VPWR net3723 sky130_fd_sc_hd__clkbuf_1
Xwire4468 net4469 VGND VGND VPWR VPWR net4468 sky130_fd_sc_hd__clkbuf_1
Xwire3734 net3735 VGND VGND VPWR VPWR net3734 sky130_fd_sc_hd__buf_1
Xwire4479 net4480 VGND VGND VPWR VPWR net4479 sky130_fd_sc_hd__clkbuf_1
X_23027_ net5062 net4647 VGND VGND VPWR VPWR _02897_ sky130_fd_sc_hd__nand2_1
Xwire3745 _03605_ VGND VGND VPWR VPWR net3745 sky130_fd_sc_hd__dlymetal6s2s_1
X_20239_ net13 _12055_ VGND VGND VPWR VPWR _12056_ sky130_fd_sc_hd__xnor2_1
Xwire3767 _02560_ VGND VGND VPWR VPWR net3767 sky130_fd_sc_hd__buf_1
Xwire3778 net3779 VGND VGND VPWR VPWR net3778 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3789 net3790 VGND VGND VPWR VPWR net3789 sky130_fd_sc_hd__buf_1
XFILLER_0_36_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14800_ net3624 net7180 net3618 VGND VGND VPWR VPWR _06917_ sky130_fd_sc_hd__or3_1
X_15780_ _07846_ _07849_ VGND VGND VPWR VPWR _07850_ sky130_fd_sc_hd__xnor2_1
X_24978_ pid_q.kp\[8\] _04718_ net1358 VGND VGND VPWR VPWR _04744_ sky130_fd_sc_hd__mux2_1
X_12992_ net7847 net1602 VGND VGND VPWR VPWR _05265_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14731_ _06827_ _06866_ net7444 VGND VGND VPWR VPWR _06867_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_169_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23929_ _03791_ _03792_ VGND VGND VPWR VPWR _03793_ sky130_fd_sc_hd__xor2_2
Xmax_length8452 net8450 VGND VGND VPWR VPWR net8452 sky130_fd_sc_hd__clkbuf_2
Xmax_length8474 net8471 VGND VGND VPWR VPWR net8474 sky130_fd_sc_hd__buf_1
X_17450_ net6736 net2577 VGND VGND VPWR VPWR _09346_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14662_ net7442 net7167 net2873 VGND VGND VPWR VPWR _06816_ sky130_fd_sc_hd__and3_1
Xmax_length8496 net8497 VGND VGND VPWR VPWR net8496 sky130_fd_sc_hd__clkbuf_2
Xmax_length7762 net7755 VGND VGND VPWR VPWR net7762 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16401_ net2628 _08459_ _08461_ net3402 _08462_ VGND VGND VPWR VPWR _08463_ sky130_fd_sc_hd__o221a_1
X_13613_ net7832 net2946 net1938 VGND VGND VPWR VPWR _05883_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17381_ _09287_ net614 _09288_ _09290_ VGND VGND VPWR VPWR _00379_ sky130_fd_sc_hd__a31o_1
XFILLER_0_157_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14593_ net3641 _06762_ VGND VGND VPWR VPWR _06767_ sky130_fd_sc_hd__nor2_1
X_19120_ net2110 net2109 VGND VGND VPWR VPWR _10957_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_184_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16332_ _08040_ net2636 net2697 net3431 VGND VGND VPWR VPWR _08395_ sky130_fd_sc_hd__o211a_1
X_13544_ _05732_ _05733_ VGND VGND VPWR VPWR _05815_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19051_ _10884_ _10886_ net2113 VGND VGND VPWR VPWR _10888_ sky130_fd_sc_hd__a21boi_1
X_16263_ net2626 net2636 net2697 net3587 VGND VGND VPWR VPWR _08327_ sky130_fd_sc_hd__o211a_1
X_13475_ _05744_ _05747_ VGND VGND VPWR VPWR _05748_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_36_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6243 net6251 VGND VGND VPWR VPWR net6243 sky130_fd_sc_hd__buf_1
X_18002_ _09026_ net6940 _09845_ _09852_ net7050 VGND VGND VPWR VPWR _09853_ sky130_fd_sc_hd__o311a_1
Xwire7061 net7058 VGND VGND VPWR VPWR net7061 sky130_fd_sc_hd__clkbuf_2
X_15214_ net2715 _07125_ VGND VGND VPWR VPWR _07288_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7072 net7066 VGND VGND VPWR VPWR net7072 sky130_fd_sc_hd__buf_1
X_16194_ _07932_ _08257_ net2682 _08258_ VGND VGND VPWR VPWR _08259_ sky130_fd_sc_hd__o211a_1
Xwire7083 net7084 VGND VGND VPWR VPWR net7083 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_140_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7094 net7095 VGND VGND VPWR VPWR net7094 sky130_fd_sc_hd__buf_1
Xwire6360 net6361 VGND VGND VPWR VPWR net6360 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire6371 cordic0.slte0.opA\[11\] VGND VGND VPWR VPWR net6371 sky130_fd_sc_hd__dlymetal6s2s_1
X_15145_ net830 _07218_ VGND VGND VPWR VPWR _07219_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_105_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6382 net6383 VGND VGND VPWR VPWR net6382 sky130_fd_sc_hd__buf_1
Xfanout5575 net5587 VGND VGND VPWR VPWR net5575 sky130_fd_sc_hd__buf_1
Xfanout4841 net4849 VGND VGND VPWR VPWR net4841 sky130_fd_sc_hd__clkbuf_1
Xfanout5586 pid_d.mult0.a\[4\] VGND VGND VPWR VPWR net5586 sky130_fd_sc_hd__buf_1
XFILLER_0_121_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6393 net6394 VGND VGND VPWR VPWR net6393 sky130_fd_sc_hd__buf_1
Xfanout4874 net4879 VGND VGND VPWR VPWR net4874 sky130_fd_sc_hd__buf_1
Xwire5670 net5671 VGND VGND VPWR VPWR net5670 sky130_fd_sc_hd__buf_1
Xfanout4885 net4908 VGND VGND VPWR VPWR net4885 sky130_fd_sc_hd__buf_1
Xwire5681 net5682 VGND VGND VPWR VPWR net5681 sky130_fd_sc_hd__clkbuf_1
X_15076_ net4099 net4096 VGND VGND VPWR VPWR _07150_ sky130_fd_sc_hd__nor2_1
X_19953_ net487 _11784_ VGND VGND VPWR VPWR _11785_ sky130_fd_sc_hd__xnor2_1
Xwire5692 net5694 VGND VGND VPWR VPWR net5692 sky130_fd_sc_hd__buf_1
XFILLER_0_120_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14027_ net7646 net1124 VGND VGND VPWR VPWR _06291_ sky130_fd_sc_hd__nand2_1
X_18904_ _10723_ net873 _10744_ VGND VGND VPWR VPWR _10745_ sky130_fd_sc_hd__a21oi_1
Xwire4991 net4992 VGND VGND VPWR VPWR net4991 sky130_fd_sc_hd__buf_1
X_19884_ _11543_ _11553_ _11609_ VGND VGND VPWR VPWR _11717_ sky130_fd_sc_hd__and3_1
X_18835_ net3222 _10677_ VGND VGND VPWR VPWR _10678_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15978_ _07935_ _07938_ _07937_ VGND VGND VPWR VPWR _08046_ sky130_fd_sc_hd__a21o_1
X_18766_ _10608_ _10456_ _10609_ _10564_ _10500_ VGND VGND VPWR VPWR _10611_ sky130_fd_sc_hd__a32o_1
X_17717_ net9200 net1216 net1454 pid_q.curr_int\[8\] VGND VGND VPWR VPWR _00422_ sky130_fd_sc_hd__a22o_1
X_14929_ net6559 net6587 matmul0.matmul_stage_inst.e\[3\] VGND VGND VPWR VPWR _07003_
+ sky130_fd_sc_hd__o21a_1
X_18697_ _10541_ _10542_ VGND VGND VPWR VPWR _10543_ sky130_fd_sc_hd__nand2_1
XFILLER_0_187_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17648_ net6707 net6746 VGND VGND VPWR VPWR _09528_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17579_ _09457_ _09438_ _09460_ VGND VGND VPWR VPWR _09461_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19318_ _11130_ _11154_ VGND VGND VPWR VPWR _11155_ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20590_ net2192 _12372_ VGND VGND VPWR VPWR _12373_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19249_ net6129 _11048_ VGND VGND VPWR VPWR _11086_ sky130_fd_sc_hd__xnor2_1
X_22260_ _02262_ _02263_ VGND VGND VPWR VPWR _02264_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21211_ net1183 _01225_ _01007_ VGND VGND VPWR VPWR _01227_ sky130_fd_sc_hd__a21o_1
XFILLER_0_170_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22191_ net2062 _02193_ _02159_ VGND VGND VPWR VPWR _02196_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21142_ net3816 _01151_ _01150_ VGND VGND VPWR VPWR _01158_ sky130_fd_sc_hd__a21oi_1
Xwire3019 net3020 VGND VGND VPWR VPWR net3019 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2307 net2308 VGND VGND VPWR VPWR net2307 sky130_fd_sc_hd__buf_1
XFILLER_0_158_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21073_ _01036_ _01041_ VGND VGND VPWR VPWR _01089_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2318 net2319 VGND VGND VPWR VPWR net2318 sky130_fd_sc_hd__buf_1
Xwire2329 _04959_ VGND VGND VPWR VPWR net2329 sky130_fd_sc_hd__buf_1
XFILLER_0_67_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24901_ pid_q.ki\[15\] net3711 net3701 net4475 VGND VGND VPWR VPWR _04692_ sky130_fd_sc_hd__a22o_1
X_20024_ net3199 _11798_ _11797_ VGND VGND VPWR VPWR _11854_ sky130_fd_sc_hd__mux2_1
Xwire1606 net1607 VGND VGND VPWR VPWR net1606 sky130_fd_sc_hd__buf_1
X_25881_ clknet_leaf_14_clk _00754_ net8620 VGND VGND VPWR VPWR pid_q.ki\[9\] sky130_fd_sc_hd__dfrtp_1
Xwire1628 _04785_ VGND VGND VPWR VPWR net1628 sky130_fd_sc_hd__buf_1
Xwire1639 _04589_ VGND VGND VPWR VPWR net1639 sky130_fd_sc_hd__clkbuf_1
X_24832_ net7484 net1009 net1017 VGND VGND VPWR VPWR _04649_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24763_ net7990 _04586_ _04587_ net1638 VGND VGND VPWR VPWR _04592_ sky130_fd_sc_hd__a31o_1
XFILLER_0_174_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21975_ _01860_ _01862_ _01982_ VGND VGND VPWR VPWR _01983_ sky130_fd_sc_hd__o21a_1
Xmax_length7036 net7037 VGND VGND VPWR VPWR net7036 sky130_fd_sc_hd__clkbuf_1
X_23714_ _03577_ _03483_ _03579_ VGND VGND VPWR VPWR _03580_ sky130_fd_sc_hd__a21o_1
X_20926_ _00939_ _00940_ _00941_ VGND VGND VPWR VPWR _00942_ sky130_fd_sc_hd__o21ai_1
X_24694_ net8034 net4265 VGND VGND VPWR VPWR _04532_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23645_ net4558 net5023 VGND VGND VPWR VPWR _03512_ sky130_fd_sc_hd__nand2_1
Xmax_length5612 net5613 VGND VGND VPWR VPWR net5612 sky130_fd_sc_hd__buf_1
X_20857_ _00869_ _00870_ net3119 VGND VGND VPWR VPWR _00873_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length5656 net5657 VGND VGND VPWR VPWR net5656 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23576_ _03441_ _03443_ VGND VGND VPWR VPWR _03444_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20788_ _12552_ _12558_ VGND VGND VPWR VPWR _12559_ sky130_fd_sc_hd__xnor2_2
Xmax_length4944 net4940 VGND VGND VPWR VPWR net4944 sky130_fd_sc_hd__buf_1
XFILLER_0_18_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire903 net904 VGND VGND VPWR VPWR net903 sky130_fd_sc_hd__buf_1
XFILLER_0_146_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25315_ clknet_leaf_80_clk _00198_ net8489 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.e\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire914 _05723_ VGND VGND VPWR VPWR net914 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22527_ net5972 net2379 net2046 VGND VGND VPWR VPWR _02526_ sky130_fd_sc_hd__and3_1
XFILLER_0_187_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire925 _04648_ VGND VGND VPWR VPWR net925 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire936 net937 VGND VGND VPWR VPWR net936 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire947 _01517_ VGND VGND VPWR VPWR net947 sky130_fd_sc_hd__buf_1
X_13260_ net7946 net3682 net2294 VGND VGND VPWR VPWR _05533_ sky130_fd_sc_hd__and3_1
Xwire958 net959 VGND VGND VPWR VPWR net958 sky130_fd_sc_hd__buf_1
X_25246_ clknet_leaf_88_clk _00129_ net8443 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.a\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_22458_ net4316 net2488 net205 VGND VGND VPWR VPWR _02460_ sky130_fd_sc_hd__and3_1
Xwire969 net970 VGND VGND VPWR VPWR net969 sky130_fd_sc_hd__clkbuf_1
X_21409_ _01420_ net757 VGND VGND VPWR VPWR _01423_ sky130_fd_sc_hd__nand2_1
X_13191_ _05448_ _05449_ _05463_ VGND VGND VPWR VPWR _05464_ sky130_fd_sc_hd__a21o_1
X_25177_ clknet_leaf_55_clk _00066_ net8728 VGND VGND VPWR VPWR svm0.periodTop\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22389_ pid_d.prev_error\[13\] net5965 VGND VGND VPWR VPWR _02392_ sky130_fd_sc_hd__xor2_1
Xwire4210 _06971_ VGND VGND VPWR VPWR net4210 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4221 net4222 VGND VGND VPWR VPWR net4221 sky130_fd_sc_hd__dlymetal6s2s_1
X_24128_ _03986_ _03989_ VGND VGND VPWR VPWR _03990_ sky130_fd_sc_hd__xnor2_1
Xwire4232 _06532_ VGND VGND VPWR VPWR net4232 sky130_fd_sc_hd__buf_1
Xwire4243 net4244 VGND VGND VPWR VPWR net4243 sky130_fd_sc_hd__clkbuf_1
Xwire4254 net4255 VGND VGND VPWR VPWR net4254 sky130_fd_sc_hd__buf_1
Xwire4265 _04928_ VGND VGND VPWR VPWR net4265 sky130_fd_sc_hd__buf_1
Xwire3520 _07066_ VGND VGND VPWR VPWR net3520 sky130_fd_sc_hd__clkbuf_1
X_24059_ _03824_ _03826_ _03921_ VGND VGND VPWR VPWR _03922_ sky130_fd_sc_hd__a21o_1
X_16950_ net7106 VGND VGND VPWR VPWR _08913_ sky130_fd_sc_hd__inv_2
Xwire3542 net3543 VGND VGND VPWR VPWR net3542 sky130_fd_sc_hd__clkbuf_1
Xwire4287 net4288 VGND VGND VPWR VPWR net4287 sky130_fd_sc_hd__clkbuf_2
Xwire3553 _07043_ VGND VGND VPWR VPWR net3553 sky130_fd_sc_hd__buf_1
Xwire4298 net4299 VGND VGND VPWR VPWR net4298 sky130_fd_sc_hd__buf_1
XFILLER_0_194_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15901_ _07874_ _07968_ _07969_ VGND VGND VPWR VPWR _07970_ sky130_fd_sc_hd__a21o_1
Xwire2830 _07080_ VGND VGND VPWR VPWR net2830 sky130_fd_sc_hd__buf_1
X_16881_ _08822_ _08844_ net6519 VGND VGND VPWR VPWR _08845_ sky130_fd_sc_hd__mux2_1
Xwire3586 _07019_ VGND VGND VPWR VPWR net3586 sky130_fd_sc_hd__buf_1
Xwire2841 net2842 VGND VGND VPWR VPWR net2841 sky130_fd_sc_hd__buf_1
XFILLER_0_95_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3597 _06984_ VGND VGND VPWR VPWR net3597 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2863 _06834_ VGND VGND VPWR VPWR net2863 sky130_fd_sc_hd__clkbuf_1
X_15832_ net2799 net3565 net1846 VGND VGND VPWR VPWR _07902_ sky130_fd_sc_hd__and3_1
X_18620_ net3230 net6957 _10387_ _10466_ VGND VGND VPWR VPWR _10467_ sky130_fd_sc_hd__a31o_1
Xwire2885 _06719_ VGND VGND VPWR VPWR net2885 sky130_fd_sc_hd__buf_1
XFILLER_0_21_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2896 net2897 VGND VGND VPWR VPWR net2896 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_154_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15763_ net1536 _07756_ _07832_ VGND VGND VPWR VPWR _07833_ sky130_fd_sc_hd__o21ai_1
X_18551_ _10398_ _10399_ net6379 VGND VGND VPWR VPWR _10400_ sky130_fd_sc_hd__mux2_1
X_12975_ _05241_ _05247_ net735 VGND VGND VPWR VPWR _05248_ sky130_fd_sc_hd__or3_1
X_17502_ net4067 _09389_ net6659 VGND VGND VPWR VPWR _09390_ sky130_fd_sc_hd__o21a_1
X_14714_ matmul0.sin\[10\] matmul0.sin\[11\] net1908 VGND VGND VPWR VPWR _06855_ sky130_fd_sc_hd__or3_1
X_18482_ net663 net659 _10331_ VGND VGND VPWR VPWR _10332_ sky130_fd_sc_hd__a21oi_2
X_15694_ _07762_ _07764_ VGND VGND VPWR VPWR _07765_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17433_ _09330_ _09331_ _08648_ VGND VGND VPWR VPWR _00390_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_185_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14645_ net7437 matmul0.cos\[4\] _06805_ VGND VGND VPWR VPWR _06807_ sky130_fd_sc_hd__and3_1
XFILLER_0_170_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length6880 net6882 VGND VGND VPWR VPWR net6880 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17364_ net669 VGND VGND VPWR VPWR _09276_ sky130_fd_sc_hd__buf_1
X_14576_ _06741_ _06746_ _06751_ VGND VGND VPWR VPWR _06752_ sky130_fd_sc_hd__a21oi_2
Xmax_length6891 net6887 VGND VGND VPWR VPWR net6891 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19103_ net3190 _10939_ VGND VGND VPWR VPWR _10940_ sky130_fd_sc_hd__xnor2_2
X_16315_ _08308_ _08357_ _08356_ VGND VGND VPWR VPWR _08378_ sky130_fd_sc_hd__a21o_1
X_13527_ _05789_ _05797_ VGND VGND VPWR VPWR _05798_ sky130_fd_sc_hd__xnor2_2
X_17295_ net7806 _09208_ VGND VGND VPWR VPWR _09209_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19034_ _10870_ VGND VGND VPWR VPWR _10871_ sky130_fd_sc_hd__buf_1
XFILLER_0_113_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout6051 cordic0.vec\[0\]\[15\] VGND VGND VPWR VPWR net6051 sky130_fd_sc_hd__buf_1
X_16246_ _08267_ _08293_ _08309_ VGND VGND VPWR VPWR _08310_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_179_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13458_ net7747 net1313 VGND VGND VPWR VPWR _05731_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout6084 net6089 VGND VGND VPWR VPWR net6084 sky130_fd_sc_hd__buf_1
XFILLER_0_51_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16177_ _08226_ _08229_ _08224_ VGND VGND VPWR VPWR _08242_ sky130_fd_sc_hd__a21o_1
X_13389_ net683 net848 VGND VGND VPWR VPWR _05662_ sky130_fd_sc_hd__xor2_2
XFILLER_0_112_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6190 net6185 VGND VGND VPWR VPWR net6190 sky130_fd_sc_hd__clkbuf_1
X_15128_ _07183_ net1278 net1277 VGND VGND VPWR VPWR _07202_ sky130_fd_sc_hd__a21oi_1
Xoutput149 net6682 VGND VGND VPWR VPWR pwmA_out sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15059_ net4105 net4101 VGND VGND VPWR VPWR _07133_ sky130_fd_sc_hd__or2_1
X_19936_ net1410 _11767_ VGND VGND VPWR VPWR _11768_ sky130_fd_sc_hd__xnor2_1
X_19867_ net6033 net6009 net2501 VGND VGND VPWR VPWR _11700_ sky130_fd_sc_hd__mux2_1
X_18818_ _10625_ _10660_ _10652_ VGND VGND VPWR VPWR _10661_ sky130_fd_sc_hd__o21bai_1
X_19798_ net2104 _11046_ _11582_ VGND VGND VPWR VPWR _11632_ sky130_fd_sc_hd__mux2_1
XFILLER_0_179_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18749_ _10541_ _10593_ VGND VGND VPWR VPWR _10594_ sky130_fd_sc_hd__xor2_1
XFILLER_0_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21760_ net5706 net5549 _01768_ _01769_ VGND VGND VPWR VPWR _01770_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20711_ _12472_ _12482_ _12483_ VGND VGND VPWR VPWR _12484_ sky130_fd_sc_hd__a21o_1
X_21691_ _01591_ _01593_ _01701_ VGND VGND VPWR VPWR _01702_ sky130_fd_sc_hd__a21oi_1
Xwire8509 net8505 VGND VGND VPWR VPWR net8509 sky130_fd_sc_hd__buf_1
X_23430_ net1675 net3059 _03196_ VGND VGND VPWR VPWR _03300_ sky130_fd_sc_hd__o21a_1
XFILLER_0_163_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20642_ net1738 _12420_ VGND VGND VPWR VPWR _12421_ sky130_fd_sc_hd__xor2_2
Xwire7808 net7809 VGND VGND VPWR VPWR net7808 sky130_fd_sc_hd__clkbuf_1
Xmax_length3506 net3507 VGND VGND VPWR VPWR net3506 sky130_fd_sc_hd__buf_1
X_23361_ _03183_ _03230_ VGND VGND VPWR VPWR _03231_ sky130_fd_sc_hd__xnor2_1
X_20573_ _12348_ _12349_ _12356_ VGND VGND VPWR VPWR _12357_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_128_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25100_ net232 net1629 _04842_ _04843_ VGND VGND VPWR VPWR _00791_ sky130_fd_sc_hd__a22o_1
X_22312_ net2057 _02315_ VGND VGND VPWR VPWR _02316_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_61_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23292_ _03006_ _03161_ VGND VGND VPWR VPWR _03162_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2827 net2828 VGND VGND VPWR VPWR net2827 sky130_fd_sc_hd__buf_1
XFILLER_0_61_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2849 _07012_ VGND VGND VPWR VPWR net2849 sky130_fd_sc_hd__buf_1
X_25031_ net7473 net2396 VGND VGND VPWR VPWR _04784_ sky130_fd_sc_hd__and2_1
XFILLER_0_132_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22243_ _02245_ _02247_ VGND VGND VPWR VPWR _02248_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22174_ net4367 _02178_ _02179_ VGND VGND VPWR VPWR _02180_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21125_ net5643 net5796 VGND VGND VPWR VPWR _01141_ sky130_fd_sc_hd__nand2_1
Xwire2104 net2105 VGND VGND VPWR VPWR net2104 sky130_fd_sc_hd__clkbuf_2
Xwire2115 net2116 VGND VGND VPWR VPWR net2115 sky130_fd_sc_hd__clkbuf_1
Xwire2126 _10546_ VGND VGND VPWR VPWR net2126 sky130_fd_sc_hd__clkbuf_1
X_25933_ clknet_leaf_25_clk _00806_ net8591 VGND VGND VPWR VPWR pid_d.prev_int\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire2137 _10263_ VGND VGND VPWR VPWR net2137 sky130_fd_sc_hd__clkbuf_1
X_21056_ net3823 _01001_ _01070_ _01071_ _01069_ VGND VGND VPWR VPWR _01072_ sky130_fd_sc_hd__o32a_1
Xwire2148 net2149 VGND VGND VPWR VPWR net2148 sky130_fd_sc_hd__buf_1
Xwire1414 _11685_ VGND VGND VPWR VPWR net1414 sky130_fd_sc_hd__clkbuf_1
Xwire1425 _11067_ VGND VGND VPWR VPWR net1425 sky130_fd_sc_hd__clkbuf_1
X_20007_ _11825_ _11824_ _11836_ VGND VGND VPWR VPWR _11837_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_185_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1436 _10392_ VGND VGND VPWR VPWR net1436 sky130_fd_sc_hd__buf_1
X_25864_ clknet_leaf_16_clk _00737_ net8619 VGND VGND VPWR VPWR pid_q.mult0.a\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1447 _09828_ VGND VGND VPWR VPWR net1447 sky130_fd_sc_hd__clkbuf_2
Xwire1458 net1459 VGND VGND VPWR VPWR net1458 sky130_fd_sc_hd__clkbuf_1
X_24815_ net5189 net1989 _04633_ VGND VGND VPWR VPWR _04638_ sky130_fd_sc_hd__a21oi_1
X_25795_ clknet_leaf_33_clk _00668_ net8678 VGND VGND VPWR VPWR pid_q.curr_int\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_24746_ net5259 VGND VGND VPWR VPWR _04577_ sky130_fd_sc_hd__inv_2
X_12760_ net7850 net1356 VGND VGND VPWR VPWR _05033_ sky130_fd_sc_hd__nand2_1
X_21958_ net5380 _01965_ VGND VGND VPWR VPWR _01966_ sky130_fd_sc_hd__nand2_1
XFILLER_0_185_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8904 net8911 VGND VGND VPWR VPWR net8904 sky130_fd_sc_hd__buf_1
XFILLER_0_178_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20909_ _00921_ _00924_ VGND VGND VPWR VPWR _00925_ sky130_fd_sc_hd__xor2_1
XFILLER_0_189_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24677_ pid_q.curr_error\[10\] net3020 net1645 VGND VGND VPWR VPWR _04521_ sky130_fd_sc_hd__and3_1
X_12691_ net2973 net2972 VGND VGND VPWR VPWR _04964_ sky130_fd_sc_hd__and2_1
X_21889_ _01744_ _01897_ VGND VGND VPWR VPWR _01898_ sky130_fd_sc_hd__nor2_1
XFILLER_0_193_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6176 net6175 VGND VGND VPWR VPWR net6176 sky130_fd_sc_hd__buf_1
X_14430_ _06626_ matmul0.b_in\[9\] net895 VGND VGND VPWR VPWR _06627_ sky130_fd_sc_hd__mux2_1
X_23628_ _03426_ _03427_ VGND VGND VPWR VPWR _03495_ sky130_fd_sc_hd__nor2_1
XFILLER_0_166_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length5475 net5476 VGND VGND VPWR VPWR net5475 sky130_fd_sc_hd__buf_1
XFILLER_0_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14361_ _06573_ VGND VGND VPWR VPWR _00076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23559_ net4664 net4920 VGND VGND VPWR VPWR _03427_ sky130_fd_sc_hd__nand2_1
Xmax_length5497 net5498 VGND VGND VPWR VPWR net5497 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire711 _11367_ VGND VGND VPWR VPWR net711 sky130_fd_sc_hd__clkbuf_1
Xwire722 _08708_ VGND VGND VPWR VPWR net722 sky130_fd_sc_hd__clkbuf_1
Xinput18 currA_in[10] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16100_ net2630 _08165_ _08105_ VGND VGND VPWR VPWR _08166_ sky130_fd_sc_hd__o21ai_1
X_13312_ net7671 net1975 net2311 VGND VGND VPWR VPWR _05585_ sky130_fd_sc_hd__and3_1
Xwire733 _05431_ VGND VGND VPWR VPWR net733 sky130_fd_sc_hd__buf_1
Xwire744 _03561_ VGND VGND VPWR VPWR net744 sky130_fd_sc_hd__buf_1
X_17080_ net1221 _09037_ VGND VGND VPWR VPWR _09038_ sky130_fd_sc_hd__nand2_1
Xinput29 currA_in[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
Xwire755 _03180_ VGND VGND VPWR VPWR net755 sky130_fd_sc_hd__buf_1
X_14292_ net66 _06518_ _06519_ net7711 VGND VGND VPWR VPWR _00061_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire766 _10338_ VGND VGND VPWR VPWR net766 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire777 _08111_ VGND VGND VPWR VPWR net777 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16031_ _08094_ _08097_ VGND VGND VPWR VPWR _08098_ sky130_fd_sc_hd__xnor2_2
Xwire788 _05766_ VGND VGND VPWR VPWR net788 sky130_fd_sc_hd__clkbuf_1
X_13243_ net847 _05515_ VGND VGND VPWR VPWR _05516_ sky130_fd_sc_hd__xor2_1
X_25229_ clknet_leaf_66_clk _00118_ net8647 VGND VGND VPWR VPWR clarke_done sky130_fd_sc_hd__dfrtp_1
Xwire799 _03305_ VGND VGND VPWR VPWR net799 sky130_fd_sc_hd__clkbuf_1
Xmax_length375 _04257_ VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13174_ _05445_ net1137 net1136 VGND VGND VPWR VPWR _05447_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4062 _08824_ VGND VGND VPWR VPWR net4062 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_176_Right_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17982_ _09831_ _09832_ _09825_ VGND VGND VPWR VPWR _09833_ sky130_fd_sc_hd__a21o_1
Xwire4073 _07682_ VGND VGND VPWR VPWR net4073 sky130_fd_sc_hd__clkbuf_1
Xwire4084 net4085 VGND VGND VPWR VPWR net4084 sky130_fd_sc_hd__clkbuf_1
Xwire3350 net3351 VGND VGND VPWR VPWR net3350 sky130_fd_sc_hd__clkbuf_1
Xwire4095 _07351_ VGND VGND VPWR VPWR net4095 sky130_fd_sc_hd__buf_1
Xwire3361 net3362 VGND VGND VPWR VPWR net3361 sky130_fd_sc_hd__clkbuf_1
X_19721_ _11544_ net604 _11553_ VGND VGND VPWR VPWR _11556_ sky130_fd_sc_hd__o21a_1
X_16933_ net6413 _08896_ VGND VGND VPWR VPWR _08897_ sky130_fd_sc_hd__or2_1
Xwire3383 _08663_ VGND VGND VPWR VPWR net3383 sky130_fd_sc_hd__buf_1
Xwire3394 _07688_ VGND VGND VPWR VPWR net3394 sky130_fd_sc_hd__buf_1
Xwire2660 _07724_ VGND VGND VPWR VPWR net2660 sky130_fd_sc_hd__buf_1
X_19652_ net1191 _11472_ _11487_ VGND VGND VPWR VPWR _11488_ sky130_fd_sc_hd__o21ai_2
Xwire2671 _07694_ VGND VGND VPWR VPWR net2671 sky130_fd_sc_hd__buf_1
X_16864_ _08827_ _08828_ net4062 VGND VGND VPWR VPWR _08829_ sky130_fd_sc_hd__mux2_1
Xwire2682 net2683 VGND VGND VPWR VPWR net2682 sky130_fd_sc_hd__clkbuf_2
Xwire2693 net2694 VGND VGND VPWR VPWR net2693 sky130_fd_sc_hd__buf_1
X_18603_ _10441_ net1069 VGND VGND VPWR VPWR _10451_ sky130_fd_sc_hd__xor2_1
Xwire1970 _04926_ VGND VGND VPWR VPWR net1970 sky130_fd_sc_hd__clkbuf_1
X_15815_ _07884_ VGND VGND VPWR VPWR _07885_ sky130_fd_sc_hd__inv_2
Xwire1981 net1985 VGND VGND VPWR VPWR net1981 sky130_fd_sc_hd__clkbuf_1
X_19583_ _11353_ _11361_ VGND VGND VPWR VPWR _11420_ sky130_fd_sc_hd__nand2_1
X_16795_ _08787_ VGND VGND VPWR VPWR _00296_ sky130_fd_sc_hd__clkbuf_1
Xwire1992 net1993 VGND VGND VPWR VPWR net1992 sky130_fd_sc_hd__buf_1
XFILLER_0_88_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15746_ _07804_ _07816_ VGND VGND VPWR VPWR _07817_ sky130_fd_sc_hd__xnor2_2
X_18534_ _10380_ net961 VGND VGND VPWR VPWR _10383_ sky130_fd_sc_hd__xnor2_1
X_12958_ _05214_ net1593 VGND VGND VPWR VPWR _05231_ sky130_fd_sc_hd__xor2_1
XFILLER_0_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18465_ _10221_ net2541 VGND VGND VPWR VPWR _10315_ sky130_fd_sc_hd__nor2_1
X_15677_ net2761 net3399 _07745_ VGND VGND VPWR VPWR _07748_ sky130_fd_sc_hd__o21a_1
X_12889_ net7804 net1610 _05091_ _05090_ VGND VGND VPWR VPWR _05162_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_8_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17416_ _09315_ net615 _09316_ _09318_ VGND VGND VPWR VPWR _00386_ sky130_fd_sc_hd__a31o_1
XFILLER_0_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14628_ _06530_ _06795_ _06796_ VGND VGND VPWR VPWR _00120_ sky130_fd_sc_hd__a21o_1
X_18396_ _10164_ _10179_ _10246_ VGND VGND VPWR VPWR _10247_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17347_ _09212_ _09259_ _09260_ VGND VGND VPWR VPWR _09261_ sky130_fd_sc_hd__mux2_1
X_14559_ net9056 net832 net448 net2886 VGND VGND VPWR VPWR _00111_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17278_ net2984 net154 _09193_ net9111 VGND VGND VPWR VPWR _00372_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19017_ net6209 net6234 VGND VGND VPWR VPWR _10854_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16229_ _08289_ _08293_ VGND VGND VPWR VPWR _08294_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_143_Right_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19919_ net3154 _11749_ _11750_ _11690_ VGND VGND VPWR VPWR _11751_ sky130_fd_sc_hd__or4b_1
XFILLER_0_139_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22930_ net5975 _02812_ net5339 VGND VGND VPWR VPWR _02820_ sky130_fd_sc_hd__a21o_1
XFILLER_0_155_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22861_ _02758_ VGND VGND VPWR VPWR _00637_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24600_ net5169 pid_q.prev_int\[15\] VGND VGND VPWR VPWR _04455_ sky130_fd_sc_hd__xor2_1
X_21812_ _01818_ _01738_ _01820_ VGND VGND VPWR VPWR _01821_ sky130_fd_sc_hd__a21o_1
XFILLER_0_195_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25580_ clknet_leaf_90_clk _00453_ net8425 VGND VGND VPWR VPWR cordic0.cos\[0\] sky130_fd_sc_hd__dfrtp_1
X_22792_ pid_d.kp\[8\] net3072 net1687 VGND VGND VPWR VPWR _02704_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24531_ net4001 _04386_ _04387_ VGND VGND VPWR VPWR _04388_ sky130_fd_sc_hd__or3_1
X_21743_ _01749_ _01752_ VGND VGND VPWR VPWR _01753_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8306 net8307 VGND VGND VPWR VPWR net8306 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24462_ _04319_ VGND VGND VPWR VPWR _04320_ sky130_fd_sc_hd__inv_2
XFILLER_0_176_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21674_ _01677_ _01684_ VGND VGND VPWR VPWR _01685_ sky130_fd_sc_hd__xnor2_2
Xwire8317 net8318 VGND VGND VPWR VPWR net8317 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8339 net8340 VGND VGND VPWR VPWR net8339 sky130_fd_sc_hd__buf_1
X_23413_ net4934 net4679 VGND VGND VPWR VPWR _03283_ sky130_fd_sc_hd__nand2_2
XFILLER_0_136_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20625_ _12405_ VGND VGND VPWR VPWR _00509_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24393_ _04251_ _04180_ pid_q.prev_error\[10\] VGND VGND VPWR VPWR _04252_ sky130_fd_sc_hd__o21ba_1
Xwire7627 net7625 VGND VGND VPWR VPWR net7627 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire7638 net7639 VGND VGND VPWR VPWR net7638 sky130_fd_sc_hd__buf_1
XFILLER_0_7_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6904 net6901 VGND VGND VPWR VPWR net6904 sky130_fd_sc_hd__buf_1
XFILLER_0_190_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23344_ net2429 _03213_ VGND VGND VPWR VPWR _03214_ sky130_fd_sc_hd__xnor2_1
Xmax_length2602 _09004_ VGND VGND VPWR VPWR net2602 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_73_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20556_ net3345 _12339_ _12340_ net6766 _08973_ VGND VGND VPWR VPWR _12341_ sky130_fd_sc_hd__a32o_1
Xmax_length2624 _08040_ VGND VGND VPWR VPWR net2624 sky130_fd_sc_hd__buf_1
XFILLER_0_85_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6948 net6951 VGND VGND VPWR VPWR net6948 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_105_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23275_ _03090_ _03140_ _03143_ _03144_ VGND VGND VPWR VPWR _03145_ sky130_fd_sc_hd__a31o_1
Xmax_length2657 _07759_ VGND VGND VPWR VPWR net2657 sky130_fd_sc_hd__buf_1
XFILLER_0_61_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20487_ net7042 net7010 net6983 net6971 net6514 net6489 VGND VGND VPWR VPWR _12275_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_132_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25014_ net4462 pid_q.curr_int\[3\] VGND VGND VPWR VPWR _04769_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_5_Left_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22226_ net2473 _02230_ VGND VGND VPWR VPWR _02231_ sky130_fd_sc_hd__xnor2_1
X_22157_ _02160_ _02161_ _02162_ VGND VGND VPWR VPWR _02163_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_110_Right_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21108_ _01092_ _01123_ VGND VGND VPWR VPWR _01124_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22088_ _02093_ _02094_ VGND VGND VPWR VPWR _02095_ sky130_fd_sc_hd__or2_1
Xwire1200 net1201 VGND VGND VPWR VPWR net1200 sky130_fd_sc_hd__buf_1
XFILLER_0_121_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1211 _10181_ VGND VGND VPWR VPWR net1211 sky130_fd_sc_hd__buf_1
X_13930_ _06192_ _06195_ VGND VGND VPWR VPWR _06196_ sky130_fd_sc_hd__xnor2_2
Xwire1222 net1223 VGND VGND VPWR VPWR net1222 sky130_fd_sc_hd__clkbuf_1
X_25916_ clknet_leaf_27_clk _00789_ net8651 VGND VGND VPWR VPWR pid_q.out\[12\] sky130_fd_sc_hd__dfrtp_1
X_21039_ net5556 _01053_ net3806 net3823 VGND VGND VPWR VPWR _01055_ sky130_fd_sc_hd__a31o_1
Xwire1233 net1234 VGND VGND VPWR VPWR net1233 sky130_fd_sc_hd__buf_1
Xwire1244 _08515_ VGND VGND VPWR VPWR net1244 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1255 _08183_ VGND VGND VPWR VPWR net1255 sky130_fd_sc_hd__clkbuf_1
Xwire1266 net1267 VGND VGND VPWR VPWR net1266 sky130_fd_sc_hd__buf_1
X_13861_ _06042_ _06126_ _06127_ VGND VGND VPWR VPWR _06128_ sky130_fd_sc_hd__a21o_1
X_25847_ clknet_leaf_20_clk _00720_ net8616 VGND VGND VPWR VPWR pid_q.mult0.b\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1277 _07201_ VGND VGND VPWR VPWR net1277 sky130_fd_sc_hd__buf_1
XFILLER_0_9_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1288 net1289 VGND VGND VPWR VPWR net1288 sky130_fd_sc_hd__clkbuf_1
X_15600_ net3551 net3514 VGND VGND VPWR VPWR _07672_ sky130_fd_sc_hd__nor2_1
Xwire1299 net1300 VGND VGND VPWR VPWR net1299 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_92_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12812_ _04955_ net1343 _04941_ VGND VGND VPWR VPWR _05085_ sky130_fd_sc_hd__a21o_1
X_16580_ _08637_ VGND VGND VPWR VPWR _00231_ sky130_fd_sc_hd__clkbuf_1
X_13792_ _06056_ _06059_ VGND VGND VPWR VPWR _06060_ sky130_fd_sc_hd__xnor2_1
X_25778_ clknet_leaf_74_clk _00651_ net8473 VGND VGND VPWR VPWR matmul0.beta_pass\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_15531_ net2701 net3399 VGND VGND VPWR VPWR _07604_ sky130_fd_sc_hd__nor2_1
X_24729_ net5273 VGND VGND VPWR VPWR _04562_ sky130_fd_sc_hd__inv_2
X_12743_ net7940 net1608 VGND VGND VPWR VPWR _05016_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8712 net8720 VGND VGND VPWR VPWR net8712 sky130_fd_sc_hd__buf_1
X_18250_ _10095_ _10096_ _10098_ net2544 VGND VGND VPWR VPWR _10101_ sky130_fd_sc_hd__nand4_1
XFILLER_0_182_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15462_ net2827 _07012_ net2820 net2686 VGND VGND VPWR VPWR _07536_ sky130_fd_sc_hd__and4_1
XFILLER_0_127_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12674_ _04936_ _04937_ VGND VGND VPWR VPWR _04947_ sky130_fd_sc_hd__xor2_1
XFILLER_0_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8756 net8763 VGND VGND VPWR VPWR net8756 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8767 net8772 VGND VGND VPWR VPWR net8767 sky130_fd_sc_hd__buf_2
X_17201_ net617 _09149_ _09150_ VGND VGND VPWR VPWR _09151_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_127_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14413_ net5272 _06608_ _06603_ net4448 _06613_ VGND VGND VPWR VPWR _06614_ sky130_fd_sc_hd__a221o_1
Xwire8840 net8841 VGND VGND VPWR VPWR net8840 sky130_fd_sc_hd__clkbuf_1
Xfanout8778 net8799 VGND VGND VPWR VPWR net8778 sky130_fd_sc_hd__buf_1
XFILLER_0_181_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18181_ net3346 _09630_ VGND VGND VPWR VPWR _10032_ sky130_fd_sc_hd__xnor2_1
Xwire8851 net8852 VGND VGND VPWR VPWR net8851 sky130_fd_sc_hd__clkbuf_1
X_15393_ _07267_ _07299_ VGND VGND VPWR VPWR _07467_ sky130_fd_sc_hd__xor2_1
X_17132_ _09075_ _09077_ net6932 VGND VGND VPWR VPWR _09087_ sky130_fd_sc_hd__a21o_1
Xwire8884 net131 VGND VGND VPWR VPWR net8884 sky130_fd_sc_hd__clkbuf_1
Xwire530 _06088_ VGND VGND VPWR VPWR net530 sky130_fd_sc_hd__buf_1
X_14344_ net8225 net3645 VGND VGND VPWR VPWR _06560_ sky130_fd_sc_hd__and2_1
Xwire541 net542 VGND VGND VPWR VPWR net541 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire552 _02323_ VGND VGND VPWR VPWR net552 sky130_fd_sc_hd__buf_1
Xmax_length3870 _11271_ VGND VGND VPWR VPWR net3870 sky130_fd_sc_hd__clkbuf_1
Xwire563 net564 VGND VGND VPWR VPWR net563 sky130_fd_sc_hd__clkbuf_1
X_17063_ _09012_ _09021_ VGND VGND VPWR VPWR _09022_ sky130_fd_sc_hd__xnor2_1
Xwire574 net575 VGND VGND VPWR VPWR net574 sky130_fd_sc_hd__buf_1
XFILLER_0_69_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14275_ net51 net2902 net2265 net9011 VGND VGND VPWR VPWR _00046_ sky130_fd_sc_hd__a22o_1
Xwire596 _03939_ VGND VGND VPWR VPWR net596 sky130_fd_sc_hd__clkbuf_1
Xmax_length3892 net3893 VGND VGND VPWR VPWR net3892 sky130_fd_sc_hd__buf_1
XFILLER_0_40_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16014_ _08077_ _08080_ VGND VGND VPWR VPWR _08082_ sky130_fd_sc_hd__or2_1
X_13226_ _05495_ _05498_ VGND VGND VPWR VPWR _05499_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13157_ _05428_ _05429_ VGND VGND VPWR VPWR _05430_ sky130_fd_sc_hd__and2b_1
XFILLER_0_109_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13088_ net919 _05360_ VGND VGND VPWR VPWR _05361_ sky130_fd_sc_hd__xor2_1
X_17965_ _09812_ net2139 VGND VGND VPWR VPWR _09816_ sky130_fd_sc_hd__xor2_1
Xwire3180 net3181 VGND VGND VPWR VPWR net3180 sky130_fd_sc_hd__buf_1
Xwire3191 _10923_ VGND VGND VPWR VPWR net3191 sky130_fd_sc_hd__buf_1
X_19704_ net6012 _11535_ _11536_ _11538_ _11539_ VGND VGND VPWR VPWR _11540_ sky130_fd_sc_hd__o221a_1
XFILLER_0_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16916_ net6369 _08879_ net6396 VGND VGND VPWR VPWR _08880_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_100_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17896_ _09739_ _09745_ _09746_ VGND VGND VPWR VPWR _09747_ sky130_fd_sc_hd__a21boi_2
Xwire2490 _12317_ VGND VGND VPWR VPWR net2490 sky130_fd_sc_hd__clkbuf_1
X_19635_ _11441_ _11471_ VGND VGND VPWR VPWR _11472_ sky130_fd_sc_hd__xnor2_2
X_16847_ _08814_ VGND VGND VPWR VPWR _00321_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_69_Left_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19566_ net3185 net2103 VGND VGND VPWR VPWR _11403_ sky130_fd_sc_hd__xnor2_2
X_16778_ _08778_ VGND VGND VPWR VPWR _00288_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18517_ net2130 _10365_ VGND VGND VPWR VPWR _10366_ sky130_fd_sc_hd__xnor2_1
X_15729_ _07775_ _07799_ VGND VGND VPWR VPWR _07800_ sky130_fd_sc_hd__xnor2_2
X_19497_ _10850_ net3897 net6177 VGND VGND VPWR VPWR _11334_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18448_ net7014 net3253 _10041_ _10241_ VGND VGND VPWR VPWR _10298_ sky130_fd_sc_hd__or4_1
XFILLER_0_145_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18379_ _10221_ _10229_ VGND VGND VPWR VPWR _10230_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_172_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20410_ _12191_ _12197_ VGND VGND VPWR VPWR _12207_ sky130_fd_sc_hd__and2_1
X_21390_ net5456 net2479 net5426 VGND VGND VPWR VPWR _01404_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_141_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_78_Left_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20341_ net1400 _12141_ net8055 VGND VGND VPWR VPWR _12144_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_183_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4809 net4806 VGND VGND VPWR VPWR net4809 sky130_fd_sc_hd__dlymetal6s2s_1
X_23060_ net4913 net4772 _02922_ _02929_ VGND VGND VPWR VPWR _02930_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20272_ _12081_ VGND VGND VPWR VPWR _00480_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22011_ _02016_ _01919_ _02017_ VGND VGND VPWR VPWR _02018_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23962_ _03700_ net1659 _03825_ VGND VGND VPWR VPWR _03826_ sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_87_Left_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25701_ clknet_leaf_5_clk _00574_ net8566 VGND VGND VPWR VPWR pid_d.mult0.b\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_22913_ _02802_ _02803_ VGND VGND VPWR VPWR _02805_ sky130_fd_sc_hd__or2_1
X_23893_ _03679_ _03680_ _03757_ VGND VGND VPWR VPWR _03758_ sky130_fd_sc_hd__a21oi_1
X_25632_ clknet_4_2__leaf_clk _00505_ net8357 VGND VGND VPWR VPWR cordic0.vec\[0\]\[4\]
+ sky130_fd_sc_hd__dfstp_1
X_22844_ _02743_ VGND VGND VPWR VPWR _00635_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_190_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25563_ clknet_leaf_64_clk _00436_ net8664 VGND VGND VPWR VPWR state\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22775_ net2035 VGND VGND VPWR VPWR _02695_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24514_ _04368_ _04370_ VGND VGND VPWR VPWR _04371_ sky130_fd_sc_hd__xnor2_1
X_21726_ pid_d.prev_int\[5\] VGND VGND VPWR VPWR _01736_ sky130_fd_sc_hd__inv_2
Xwire8103 net8104 VGND VGND VPWR VPWR net8103 sky130_fd_sc_hd__clkbuf_1
X_25494_ clknet_leaf_44_clk _00374_ net8786 VGND VGND VPWR VPWR svm0.calc_ready sky130_fd_sc_hd__dfrtp_1
Xwire8114 net8115 VGND VGND VPWR VPWR net8114 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8125 net8126 VGND VGND VPWR VPWR net8125 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24445_ net4555 net4808 _04301_ VGND VGND VPWR VPWR _04303_ sky130_fd_sc_hd__a21oi_1
Xwire8136 net8137 VGND VGND VPWR VPWR net8136 sky130_fd_sc_hd__clkbuf_1
X_21657_ net5718 net5538 VGND VGND VPWR VPWR _01668_ sky130_fd_sc_hd__nand2_1
Xwire7402 net7403 VGND VGND VPWR VPWR net7402 sky130_fd_sc_hd__clkbuf_1
Xwire8147 net8148 VGND VGND VPWR VPWR net8147 sky130_fd_sc_hd__clkbuf_1
Xwire8158 net8159 VGND VGND VPWR VPWR net8158 sky130_fd_sc_hd__clkbuf_1
Xwire7413 matmul0.matmul_stage_inst.c\[5\] VGND VGND VPWR VPWR net7413 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_96_Left_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8169 net8170 VGND VGND VPWR VPWR net8169 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7424 matmul0.matmul_stage_inst.b\[7\] VGND VGND VPWR VPWR net7424 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6701 net6702 VGND VGND VPWR VPWR net6701 sky130_fd_sc_hd__clkbuf_2
X_20608_ _12366_ _12387_ net6195 VGND VGND VPWR VPWR _12389_ sky130_fd_sc_hd__o21a_1
Xmax_length3133 net3134 VGND VGND VPWR VPWR net3133 sky130_fd_sc_hd__clkbuf_1
Xwire7446 net7443 VGND VGND VPWR VPWR net7446 sky130_fd_sc_hd__buf_1
Xwire6712 net6713 VGND VGND VPWR VPWR net6712 sky130_fd_sc_hd__dlymetal6s2s_1
X_24376_ _04233_ _04234_ VGND VGND VPWR VPWR _04235_ sky130_fd_sc_hd__xor2_1
XFILLER_0_145_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21588_ net1721 _01599_ VGND VGND VPWR VPWR _01600_ sky130_fd_sc_hd__xnor2_1
Xwire7457 net7455 VGND VGND VPWR VPWR net7457 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire6723 net6724 VGND VGND VPWR VPWR net6723 sky130_fd_sc_hd__clkbuf_1
Xwire7468 net7466 VGND VGND VPWR VPWR net7468 sky130_fd_sc_hd__buf_1
Xwire6734 net6735 VGND VGND VPWR VPWR net6734 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire6745 svm0.rising VGND VGND VPWR VPWR net6745 sky130_fd_sc_hd__clkbuf_1
X_23327_ net4888 VGND VGND VPWR VPWR _03197_ sky130_fd_sc_hd__inv_2
X_20539_ net6310 net1484 net2082 VGND VGND VPWR VPWR _12324_ sky130_fd_sc_hd__mux2_1
Xwire6756 net6757 VGND VGND VPWR VPWR net6756 sky130_fd_sc_hd__buf_1
Xwire6767 net6768 VGND VGND VPWR VPWR net6767 sky130_fd_sc_hd__buf_1
X_14060_ _06290_ _06309_ _06322_ VGND VGND VPWR VPWR _06323_ sky130_fd_sc_hd__o21ai_4
Xwire6789 net6788 VGND VGND VPWR VPWR net6789 sky130_fd_sc_hd__clkbuf_2
X_23258_ _03124_ _03126_ _03127_ VGND VGND VPWR VPWR _03128_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_104_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13011_ _05280_ _05166_ _05167_ net850 _05283_ VGND VGND VPWR VPWR _05284_ sky130_fd_sc_hd__o32a_1
X_22209_ _02210_ _02213_ VGND VGND VPWR VPWR _02214_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23189_ _03058_ _03039_ VGND VGND VPWR VPWR _03059_ sky130_fd_sc_hd__xor2_1
XFILLER_0_101_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17750_ net6974 net3268 VGND VGND VPWR VPWR _09601_ sky130_fd_sc_hd__xnor2_2
X_14962_ net6634 matmul0.matmul_stage_inst.d\[2\] net7417 net6538 VGND VGND VPWR VPWR
+ _07036_ sky130_fd_sc_hd__a22o_1
Xhold7 matmul0.matmul_stage_inst.a\[0\] VGND VGND VPWR VPWR net8960 sky130_fd_sc_hd__dlygate4sd3_1
Xwire1030 _03321_ VGND VGND VPWR VPWR net1030 sky130_fd_sc_hd__clkbuf_1
Xwire1041 net1042 VGND VGND VPWR VPWR net1041 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_57_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1052 _00818_ VGND VGND VPWR VPWR net1052 sky130_fd_sc_hd__buf_1
X_16701_ _08728_ _08724_ _08729_ VGND VGND VPWR VPWR _08730_ sky130_fd_sc_hd__a21o_1
X_13913_ net1950 _06177_ _06178_ VGND VGND VPWR VPWR _06179_ sky130_fd_sc_hd__a21oi_1
X_17681_ net1791 _09560_ VGND VGND VPWR VPWR _09561_ sky130_fd_sc_hd__nand2_1
Xwire1063 _11205_ VGND VGND VPWR VPWR net1063 sky130_fd_sc_hd__clkbuf_1
X_14893_ net4216 net4214 VGND VGND VPWR VPWR _06967_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1074 net1075 VGND VGND VPWR VPWR net1074 sky130_fd_sc_hd__buf_1
Xwire1085 _08292_ VGND VGND VPWR VPWR net1085 sky130_fd_sc_hd__buf_1
XFILLER_0_96_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19420_ net6265 net3886 VGND VGND VPWR VPWR _11257_ sky130_fd_sc_hd__nor2_1
Xwire1096 _07981_ VGND VGND VPWR VPWR net1096 sky130_fd_sc_hd__clkbuf_1
X_13844_ net839 _06110_ VGND VGND VPWR VPWR _06111_ sky130_fd_sc_hd__xnor2_1
X_16632_ _08670_ VGND VGND VPWR VPWR _00250_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19351_ _11187_ _11134_ net2512 VGND VGND VPWR VPWR _11188_ sky130_fd_sc_hd__o21ai_1
X_13775_ _05965_ _05966_ _05968_ _05969_ VGND VGND VPWR VPWR _06043_ sky130_fd_sc_hd__or4_1
X_16563_ _08600_ _08621_ VGND VGND VPWR VPWR _08622_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_186_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18302_ _10105_ _10100_ _10101_ VGND VGND VPWR VPWR _10153_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_167_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12726_ net1611 _04979_ _04994_ _04997_ VGND VGND VPWR VPWR _04999_ sky130_fd_sc_hd__a211o_1
X_15514_ net1538 _07585_ _07586_ VGND VGND VPWR VPWR _07587_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19282_ net6294 net3213 net3902 VGND VGND VPWR VPWR _11119_ sky130_fd_sc_hd__a21o_1
X_16494_ net1086 net1078 _08553_ VGND VGND VPWR VPWR _08554_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_45_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout8564 net8594 VGND VGND VPWR VPWR net8564 sky130_fd_sc_hd__buf_1
X_18233_ _10077_ _09809_ VGND VGND VPWR VPWR _10084_ sky130_fd_sc_hd__nand2_1
X_15445_ _06974_ net4201 net4092 net4089 VGND VGND VPWR VPWR _07519_ sky130_fd_sc_hd__o22a_1
X_12657_ net2977 VGND VGND VPWR VPWR _04930_ sky130_fd_sc_hd__clkbuf_1
Xfanout8575 net8592 VGND VGND VPWR VPWR net8575 sky130_fd_sc_hd__buf_1
XFILLER_0_167_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8670 net8669 VGND VGND VPWR VPWR net8670 sky130_fd_sc_hd__buf_1
XFILLER_0_4_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18164_ _10001_ _10008_ _10006_ VGND VGND VPWR VPWR _10015_ sky130_fd_sc_hd__or3b_1
X_15376_ _07437_ _07446_ _07449_ _07441_ VGND VGND VPWR VPWR _07450_ sky130_fd_sc_hd__a22o_1
XFILLER_0_182_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12588_ _04871_ VGND VGND VPWR VPWR _00010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17115_ net6470 net6462 VGND VGND VPWR VPWR _09071_ sky130_fd_sc_hd__nor2_1
Xwire360 net361 VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__clkbuf_1
X_14327_ _06547_ VGND VGND VPWR VPWR _00068_ sky130_fd_sc_hd__clkbuf_1
Xwire7980 net7981 VGND VGND VPWR VPWR net7980 sky130_fd_sc_hd__clkbuf_2
X_18095_ net2548 _09944_ _09945_ VGND VGND VPWR VPWR _09946_ sky130_fd_sc_hd__a21oi_1
Xwire7991 net7992 VGND VGND VPWR VPWR net7991 sky130_fd_sc_hd__clkbuf_1
Xwire371 _05681_ VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__clkbuf_1
Xwire382 _10402_ VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__clkbuf_1
Xwire393 net394 VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__clkbuf_1
X_17046_ net6474 net6462 VGND VGND VPWR VPWR _09005_ sky130_fd_sc_hd__or2_1
XFILLER_0_187_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14258_ net6451 VGND VGND VPWR VPWR _06512_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13209_ _05405_ _05481_ VGND VGND VPWR VPWR _05482_ sky130_fd_sc_hd__nand2_1
X_14189_ _06442_ _06448_ VGND VGND VPWR VPWR _06449_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18997_ _10819_ _10833_ VGND VGND VPWR VPWR _10834_ sky130_fd_sc_hd__or2b_1
X_17948_ _09798_ _09676_ net6997 VGND VGND VPWR VPWR _09799_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_136_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17879_ net6844 _09729_ VGND VGND VPWR VPWR _09730_ sky130_fd_sc_hd__xor2_1
XFILLER_0_45_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19618_ net3907 net3868 net6183 VGND VGND VPWR VPWR _11455_ sky130_fd_sc_hd__a21o_1
X_20890_ _00900_ net2481 VGND VGND VPWR VPWR _00906_ sky130_fd_sc_hd__or2_1
X_19549_ net6158 _10944_ _11385_ net3915 _10977_ VGND VGND VPWR VPWR _11386_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22560_ net2459 VGND VGND VPWR VPWR _02544_ sky130_fd_sc_hd__buf_1
XFILLER_0_152_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21511_ net860 _01522_ _01523_ VGND VGND VPWR VPWR _01524_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22491_ _02419_ _02424_ _02491_ VGND VGND VPWR VPWR _02492_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_185_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24230_ net4789 _04090_ VGND VGND VPWR VPWR _04091_ sky130_fd_sc_hd__xnor2_1
X_21442_ net5739 net5542 VGND VGND VPWR VPWR _01455_ sky130_fd_sc_hd__nand2_2
Xwire6019 net6020 VGND VGND VPWR VPWR net6019 sky130_fd_sc_hd__buf_1
XFILLER_0_145_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24161_ _03869_ _03937_ VGND VGND VPWR VPWR _04023_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5307 net5308 VGND VGND VPWR VPWR net5307 sky130_fd_sc_hd__clkbuf_1
X_21373_ _01284_ _01286_ _01282_ VGND VGND VPWR VPWR _01387_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_160_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5318 net5319 VGND VGND VPWR VPWR net5318 sky130_fd_sc_hd__clkbuf_1
Xwire5329 net5330 VGND VGND VPWR VPWR net5329 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23112_ _02973_ _02978_ _02981_ VGND VGND VPWR VPWR _02982_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_142_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4606 net4607 VGND VGND VPWR VPWR net4606 sky130_fd_sc_hd__buf_1
X_20324_ _12126_ _12127_ VGND VGND VPWR VPWR _12128_ sky130_fd_sc_hd__nand2_1
Xwire4617 net4618 VGND VGND VPWR VPWR net4617 sky130_fd_sc_hd__buf_1
X_24092_ pid_q.prev_int\[7\] VGND VGND VPWR VPWR _03954_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4628 net4629 VGND VGND VPWR VPWR net4628 sky130_fd_sc_hd__clkbuf_1
X_23043_ _02909_ _02910_ _02912_ VGND VGND VPWR VPWR _02913_ sky130_fd_sc_hd__a21bo_1
Xwire3905 _10803_ VGND VGND VPWR VPWR net3905 sky130_fd_sc_hd__buf_1
Xwire3916 net3917 VGND VGND VPWR VPWR net3916 sky130_fd_sc_hd__buf_1
X_20255_ _12068_ VGND VGND VPWR VPWR _00476_ sky130_fd_sc_hd__clkbuf_1
Xwire3927 net3931 VGND VGND VPWR VPWR net3927 sky130_fd_sc_hd__buf_1
XFILLER_0_12_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3938 _10045_ VGND VGND VPWR VPWR net3938 sky130_fd_sc_hd__clkbuf_1
Xwire3949 net3950 VGND VGND VPWR VPWR net3949 sky130_fd_sc_hd__dlymetal6s2s_1
X_20186_ _12010_ _12011_ VGND VGND VPWR VPWR _12012_ sky130_fd_sc_hd__or2b_1
X_24994_ net2147 VGND VGND VPWR VPWR _04752_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23945_ net4541 net4972 VGND VGND VPWR VPWR _03809_ sky130_fd_sc_hd__nand2_1
X_23876_ net4729 net3048 _03740_ VGND VGND VPWR VPWR _03741_ sky130_fd_sc_hd__o21a_1
XFILLER_0_168_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length8678 net8679 VGND VGND VPWR VPWR net8678 sky130_fd_sc_hd__buf_1
X_25615_ clknet_leaf_109_clk _00488_ net8346 VGND VGND VPWR VPWR cordic0.slte0.opA\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_22827_ net5366 net5984 net5986 pid_d.out\[0\] VGND VGND VPWR VPWR _02728_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_6_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13560_ _05822_ _05829_ VGND VGND VPWR VPWR _05831_ sky130_fd_sc_hd__nand2_1
X_25546_ clknet_leaf_28_clk _00426_ net8652 VGND VGND VPWR VPWR pid_q.prev_int\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_22758_ _02683_ VGND VGND VPWR VPWR _00609_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21709_ _01612_ _01613_ _01719_ VGND VGND VPWR VPWR _01720_ sky130_fd_sc_hd__o21a_1
X_13491_ net1933 VGND VGND VPWR VPWR _05764_ sky130_fd_sc_hd__clkbuf_1
X_25477_ clknet_leaf_48_clk _00357_ net8762 VGND VGND VPWR VPWR svm0.tB\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22689_ _02634_ VGND VGND VPWR VPWR _00589_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7210 net7212 VGND VGND VPWR VPWR net7210 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15230_ _06992_ net4186 VGND VGND VPWR VPWR _07304_ sky130_fd_sc_hd__or2_1
X_24428_ _04206_ _04211_ _04285_ VGND VGND VPWR VPWR _04286_ sky130_fd_sc_hd__a21o_1
Xwire7221 net7222 VGND VGND VPWR VPWR net7221 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7232 net7233 VGND VGND VPWR VPWR net7232 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7243 net7248 VGND VGND VPWR VPWR net7243 sky130_fd_sc_hd__clkbuf_1
Xfanout6447 state\[1\] VGND VGND VPWR VPWR net6447 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_81_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7254 net7255 VGND VGND VPWR VPWR net7254 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7265 net7266 VGND VGND VPWR VPWR net7265 sky130_fd_sc_hd__buf_1
Xwire6520 net6517 VGND VGND VPWR VPWR net6520 sky130_fd_sc_hd__buf_1
Xfanout5724 net5735 VGND VGND VPWR VPWR net5724 sky130_fd_sc_hd__buf_1
Xfanout6469 cordic0.gm0.iter\[3\] VGND VGND VPWR VPWR net6469 sky130_fd_sc_hd__buf_1
X_15161_ net1886 _07234_ VGND VGND VPWR VPWR _07235_ sky130_fd_sc_hd__or2_1
X_24359_ net2405 _04135_ _04128_ VGND VGND VPWR VPWR _04218_ sky130_fd_sc_hd__o21a_1
Xwire7276 net7277 VGND VGND VPWR VPWR net7276 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6542 net6539 VGND VGND VPWR VPWR net6542 sky130_fd_sc_hd__buf_1
Xwire7287 net7288 VGND VGND VPWR VPWR net7287 sky130_fd_sc_hd__buf_1
Xwire7298 net7299 VGND VGND VPWR VPWR net7298 sky130_fd_sc_hd__clkbuf_1
X_14112_ net1566 VGND VGND VPWR VPWR _06374_ sky130_fd_sc_hd__buf_1
Xwire6564 net6565 VGND VGND VPWR VPWR net6564 sky130_fd_sc_hd__buf_1
Xwire6575 net6578 VGND VGND VPWR VPWR net6575 sky130_fd_sc_hd__buf_1
Xwire5841 net5842 VGND VGND VPWR VPWR net5841 sky130_fd_sc_hd__dlymetal6s2s_1
X_15092_ _07073_ _07165_ VGND VGND VPWR VPWR _07166_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5863 net5864 VGND VGND VPWR VPWR net5863 sky130_fd_sc_hd__clkbuf_1
X_14043_ _06227_ _06232_ _06306_ VGND VGND VPWR VPWR _06307_ sky130_fd_sc_hd__a21oi_2
X_18920_ _10716_ _10738_ VGND VGND VPWR VPWR _10760_ sky130_fd_sc_hd__nor2_1
Xwire5874 net5867 VGND VGND VPWR VPWR net5874 sky130_fd_sc_hd__buf_1
XFILLER_0_120_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5885 net5886 VGND VGND VPWR VPWR net5885 sky130_fd_sc_hd__clkbuf_1
Xwire5896 net5897 VGND VGND VPWR VPWR net5896 sky130_fd_sc_hd__buf_1
XFILLER_0_157_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18851_ _10623_ _10656_ VGND VGND VPWR VPWR _10694_ sky130_fd_sc_hd__nand2b_1
X_17802_ net2562 _09652_ VGND VGND VPWR VPWR _09653_ sky130_fd_sc_hd__and2_1
X_18782_ _10572_ _10593_ _10541_ VGND VGND VPWR VPWR _10626_ sky130_fd_sc_hd__a21bo_1
X_15994_ _08037_ net883 VGND VGND VPWR VPWR _08062_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17733_ net2599 _09589_ VGND VGND VPWR VPWR _00433_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14945_ _07018_ VGND VGND VPWR VPWR _07019_ sky130_fd_sc_hd__buf_1
X_17664_ svm0.counter\[3\] svm0.tA\[3\] VGND VGND VPWR VPWR _09544_ sky130_fd_sc_hd__xor2_1
X_14876_ matmul0.b\[10\] matmul0.matmul_stage_inst.f\[10\] net3604 VGND VGND VPWR
+ VPWR _06956_ sky130_fd_sc_hd__mux2_1
XFILLER_0_187_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19403_ net1192 _11229_ _11239_ VGND VGND VPWR VPWR _11240_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16615_ _08657_ VGND VGND VPWR VPWR _00246_ sky130_fd_sc_hd__clkbuf_1
X_13827_ net7679 net1943 net2292 VGND VGND VPWR VPWR _06094_ sky130_fd_sc_hd__and3_1
X_17595_ net4030 svm0.tB\[15\] _09475_ VGND VGND VPWR VPWR _09476_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_159_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19334_ net6262 net6229 VGND VGND VPWR VPWR _11171_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13758_ _05939_ _05940_ net7741 net1588 VGND VGND VPWR VPWR _06026_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_31_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16546_ net2634 net2631 VGND VGND VPWR VPWR _08605_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12709_ net7883 net2351 net2347 VGND VGND VPWR VPWR _04982_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19265_ _10897_ _11101_ VGND VGND VPWR VPWR _11102_ sky130_fd_sc_hd__xnor2_1
X_13689_ _05900_ _05902_ _05904_ VGND VGND VPWR VPWR _05958_ sky130_fd_sc_hd__o21a_1
X_16477_ net671 _08534_ VGND VGND VPWR VPWR _08538_ sky130_fd_sc_hd__and2b_1
Xfanout8383 net8386 VGND VGND VPWR VPWR net8383 sky130_fd_sc_hd__clkbuf_2
X_18216_ net3232 _10064_ _10066_ VGND VGND VPWR VPWR _10067_ sky130_fd_sc_hd__o21ai_1
Xfanout8394 net8414 VGND VGND VPWR VPWR net8394 sky130_fd_sc_hd__buf_1
Xfanout7660 net7665 VGND VGND VPWR VPWR net7660 sky130_fd_sc_hd__clkbuf_1
X_15428_ _07496_ _07501_ VGND VGND VPWR VPWR _07502_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_171_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19196_ _10903_ _11032_ VGND VGND VPWR VPWR _11033_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18147_ _09872_ net2549 VGND VGND VPWR VPWR _09998_ sky130_fd_sc_hd__or2_1
X_15359_ _07412_ _07415_ _07431_ _07432_ VGND VGND VPWR VPWR _07433_ sky130_fd_sc_hd__nand4_1
XFILLER_0_13_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout6970 net6980 VGND VGND VPWR VPWR net6970 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6981 net6992 VGND VGND VPWR VPWR net6981 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_14_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold204 svm0.tC\[13\] VGND VGND VPWR VPWR net9157 sky130_fd_sc_hd__dlygate4sd3_1
Xwire190 _06270_ VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__buf_1
Xhold215 cordic0.slte0.opA\[5\] VGND VGND VPWR VPWR net9168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 pid_q.prev_error\[13\] VGND VGND VPWR VPWR net9179 sky130_fd_sc_hd__dlygate4sd3_1
X_18078_ _09905_ _09926_ _09928_ VGND VGND VPWR VPWR _09929_ sky130_fd_sc_hd__a21oi_1
Xhold237 svm0.tA\[15\] VGND VGND VPWR VPWR net9190 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold248 pid_q.prev_int\[11\] VGND VGND VPWR VPWR net9201 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold259 pid_q.prev_int\[5\] VGND VGND VPWR VPWR net9212 sky130_fd_sc_hd__dlygate4sd3_1
X_17029_ net5989 _08986_ net2603 _08924_ VGND VGND VPWR VPWR _08989_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20040_ _11850_ _11869_ VGND VGND VPWR VPWR _11870_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21991_ _01892_ _01899_ VGND VGND VPWR VPWR _01999_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23730_ _03526_ _03528_ _03527_ VGND VGND VPWR VPWR _03596_ sky130_fd_sc_hd__o21a_1
X_20942_ _00909_ _00957_ VGND VGND VPWR VPWR _00958_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_178_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23661_ net4598 net4964 VGND VGND VPWR VPWR _03528_ sky130_fd_sc_hd__nand2_1
XFILLER_0_163_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20873_ _12546_ _00888_ VGND VGND VPWR VPWR _00889_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_178_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25400_ clknet_leaf_69_clk _00283_ net8484 VGND VGND VPWR VPWR matmul0.a\[3\] sky130_fd_sc_hd__dfrtp_1
X_22612_ net9043 _02544_ net2042 _02584_ VGND VGND VPWR VPWR _00562_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23592_ _03455_ _03459_ VGND VGND VPWR VPWR _03460_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_118_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25331_ clknet_leaf_76_clk _00214_ net8462 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.f\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_22543_ net5967 net3016 net2048 VGND VGND VPWR VPWR _02534_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25262_ clknet_leaf_76_clk _00145_ net8458 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.b\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_22474_ _02472_ _02473_ net5689 VGND VGND VPWR VPWR _02475_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_161_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24213_ _04067_ _04073_ VGND VGND VPWR VPWR _04074_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_133_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21425_ _01436_ _01437_ VGND VGND VPWR VPWR _01438_ sky130_fd_sc_hd__and2_1
X_25193_ clknet_leaf_58_clk _00082_ net8721 VGND VGND VPWR VPWR matmul0.a_in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire5104 net5105 VGND VGND VPWR VPWR net5104 sky130_fd_sc_hd__buf_1
Xwire5115 net5116 VGND VGND VPWR VPWR net5115 sky130_fd_sc_hd__buf_1
X_24144_ _03909_ _03916_ _03914_ VGND VGND VPWR VPWR _04006_ sky130_fd_sc_hd__o21a_1
Xwire5137 net5138 VGND VGND VPWR VPWR net5137 sky130_fd_sc_hd__clkbuf_1
X_21356_ _01364_ _01369_ VGND VGND VPWR VPWR _01370_ sky130_fd_sc_hd__xnor2_2
Xwire5148 net5149 VGND VGND VPWR VPWR net5148 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4403 net4404 VGND VGND VPWR VPWR net4403 sky130_fd_sc_hd__clkbuf_1
Xwire5159 net5160 VGND VGND VPWR VPWR net5159 sky130_fd_sc_hd__clkbuf_1
Xwire4414 net4415 VGND VGND VPWR VPWR net4414 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4425 net4426 VGND VGND VPWR VPWR net4425 sky130_fd_sc_hd__clkbuf_1
X_20307_ net6479 _12108_ _12111_ VGND VGND VPWR VPWR _12112_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4436 net4437 VGND VGND VPWR VPWR net4436 sky130_fd_sc_hd__clkbuf_1
X_24075_ _03935_ _03937_ VGND VGND VPWR VPWR _03938_ sky130_fd_sc_hd__xor2_1
Xwire3702 net3703 VGND VGND VPWR VPWR net3702 sky130_fd_sc_hd__clkbuf_2
X_21287_ _01276_ _01301_ VGND VGND VPWR VPWR _01302_ sky130_fd_sc_hd__xnor2_1
Xwire3713 net3714 VGND VGND VPWR VPWR net3713 sky130_fd_sc_hd__clkbuf_1
Xwire4458 net4459 VGND VGND VPWR VPWR net4458 sky130_fd_sc_hd__clkbuf_1
Xwire3724 net3725 VGND VGND VPWR VPWR net3724 sky130_fd_sc_hd__clkbuf_1
Xwire4469 net4470 VGND VGND VPWR VPWR net4469 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23026_ net5037 net4684 VGND VGND VPWR VPWR _02896_ sky130_fd_sc_hd__nand2_1
Xwire3735 net3736 VGND VGND VPWR VPWR net3735 sky130_fd_sc_hd__clkbuf_1
Xwire3746 _03456_ VGND VGND VPWR VPWR net3746 sky130_fd_sc_hd__clkbuf_1
X_20238_ net8122 _12054_ VGND VGND VPWR VPWR _12055_ sky130_fd_sc_hd__nor2_1
Xwire3757 _02866_ VGND VGND VPWR VPWR net3757 sky130_fd_sc_hd__buf_1
X_20169_ _11954_ _11992_ _11994_ net868 VGND VGND VPWR VPWR _11995_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_157_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12991_ _05176_ _05181_ _05263_ VGND VGND VPWR VPWR _05264_ sky130_fd_sc_hd__o21a_1
X_24977_ _04743_ VGND VGND VPWR VPWR _00768_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14730_ net3613 net7160 net7163 VGND VGND VPWR VPWR _06866_ sky130_fd_sc_hd__and3_1
X_23928_ net4676 net4799 VGND VGND VPWR VPWR _03792_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14661_ net9021 net2872 _06815_ VGND VGND VPWR VPWR _00134_ sky130_fd_sc_hd__a21o_1
X_23859_ _03622_ _03627_ _03723_ VGND VGND VPWR VPWR _03724_ sky130_fd_sc_hd__a21o_1
XFILLER_0_52_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13612_ net7811 net1578 VGND VGND VPWR VPWR _05882_ sky130_fd_sc_hd__and2_1
X_16400_ net2791 net2621 net2642 net2772 net2245 VGND VGND VPWR VPWR _08462_ sky130_fd_sc_hd__a2111o_1
Xmax_length7785 net7777 VGND VGND VPWR VPWR net7785 sky130_fd_sc_hd__buf_1
X_17380_ net612 _09289_ _09287_ VGND VGND VPWR VPWR _09290_ sky130_fd_sc_hd__a21oi_1
X_14592_ net1989 _06762_ net281 VGND VGND VPWR VPWR _06766_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_184_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13543_ net7747 net1598 _05732_ _05733_ VGND VGND VPWR VPWR _05814_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_137_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16331_ net2626 net2632 net3424 net3421 VGND VGND VPWR VPWR _08394_ sky130_fd_sc_hd__o211a_1
X_25529_ clknet_leaf_45_clk _00409_ net8791 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6200 net6206 VGND VGND VPWR VPWR net6200 sky130_fd_sc_hd__buf_1
X_19050_ net6178 net6220 net6120 _10872_ _10873_ VGND VGND VPWR VPWR _10887_ sky130_fd_sc_hd__a311o_1
X_16262_ net2655 net2632 net3424 net3431 VGND VGND VPWR VPWR _08326_ sky130_fd_sc_hd__o211a_1
X_13474_ _05745_ _05746_ VGND VGND VPWR VPWR _05747_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout6233 cordic0.vec\[0\]\[6\] VGND VGND VPWR VPWR net6233 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18001_ _09847_ _09848_ net3237 VGND VGND VPWR VPWR _09852_ sky130_fd_sc_hd__a21o_1
Xwire7040 net7041 VGND VGND VPWR VPWR net7040 sky130_fd_sc_hd__buf_1
X_15213_ net3513 net3505 VGND VGND VPWR VPWR _07287_ sky130_fd_sc_hd__nor2_1
Xwire7051 net7052 VGND VGND VPWR VPWR net7051 sky130_fd_sc_hd__buf_1
X_16193_ net2670 VGND VGND VPWR VPWR _08258_ sky130_fd_sc_hd__buf_1
Xfanout5532 pid_d.mult0.a\[7\] VGND VGND VPWR VPWR net5532 sky130_fd_sc_hd__clkbuf_1
Xwire7084 net7085 VGND VGND VPWR VPWR net7084 sky130_fd_sc_hd__clkbuf_1
X_15144_ net991 _07213_ _07217_ VGND VGND VPWR VPWR _07218_ sky130_fd_sc_hd__o21ba_1
Xwire7095 net7093 VGND VGND VPWR VPWR net7095 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire6361 net6362 VGND VGND VPWR VPWR net6361 sky130_fd_sc_hd__buf_1
XFILLER_0_11_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6372 cordic0.slte0.opA\[10\] VGND VGND VPWR VPWR net6372 sky130_fd_sc_hd__buf_1
Xwire6383 net6384 VGND VGND VPWR VPWR net6383 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6394 net6395 VGND VGND VPWR VPWR net6394 sky130_fd_sc_hd__clkbuf_1
Xwire5660 net5661 VGND VGND VPWR VPWR net5660 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15075_ net4120 net4115 VGND VGND VPWR VPWR _07149_ sky130_fd_sc_hd__nor2_1
X_19952_ _11782_ _11783_ VGND VGND VPWR VPWR _11784_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5682 net5683 VGND VGND VPWR VPWR net5682 sky130_fd_sc_hd__clkbuf_1
Xfanout4897 net4903 VGND VGND VPWR VPWR net4897 sky130_fd_sc_hd__buf_1
Xwire5693 net5689 VGND VGND VPWR VPWR net5693 sky130_fd_sc_hd__buf_1
X_14026_ _06284_ _06289_ VGND VGND VPWR VPWR _06290_ sky130_fd_sc_hd__xnor2_2
X_18903_ net658 _10664_ _10723_ net873 net657 VGND VGND VPWR VPWR _10744_ sky130_fd_sc_hd__o221a_1
X_19883_ _11661_ net708 VGND VGND VPWR VPWR _11716_ sky130_fd_sc_hd__or2_1
Xwire4992 net4993 VGND VGND VPWR VPWR net4992 sky130_fd_sc_hd__clkbuf_1
X_18834_ net6877 net6796 VGND VGND VPWR VPWR _10677_ sky130_fd_sc_hd__xor2_4
X_18765_ _10608_ _10456_ _10609_ net605 VGND VGND VPWR VPWR _10610_ sky130_fd_sc_hd__o211a_1
XFILLER_0_175_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15977_ _07951_ _07954_ _08044_ VGND VGND VPWR VPWR _08045_ sky130_fd_sc_hd__o21a_1
XFILLER_0_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17716_ net9221 net1216 net1454 net5178 VGND VGND VPWR VPWR _00421_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14928_ net6619 net6644 matmul0.matmul_stage_inst.f\[3\] VGND VGND VPWR VPWR _07002_
+ sky130_fd_sc_hd__o21a_1
X_18696_ net6778 net1760 VGND VGND VPWR VPWR _10542_ sky130_fd_sc_hd__or2_1
X_17647_ net4026 svm0.tA\[8\] VGND VGND VPWR VPWR _09527_ sky130_fd_sc_hd__nor2_1
X_14859_ net7188 matmul0.matmul_stage_inst.f\[2\] _06939_ VGND VGND VPWR VPWR _06947_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17578_ _09434_ _09436_ _09458_ _09459_ VGND VGND VPWR VPWR _09460_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19317_ net2512 _11134_ _11139_ _11153_ VGND VGND VPWR VPWR _11154_ sky130_fd_sc_hd__o22a_1
XFILLER_0_128_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16529_ _08548_ _08588_ VGND VGND VPWR VPWR _08589_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19248_ net6201 _11082_ _11084_ net3178 VGND VGND VPWR VPWR _11085_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19179_ net3187 _10934_ _11015_ VGND VGND VPWR VPWR _11016_ sky130_fd_sc_hd__a21o_1
XFILLER_0_182_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21210_ _01007_ _01224_ _01225_ _01008_ VGND VGND VPWR VPWR _01226_ sky130_fd_sc_hd__o2bb2a_1
X_22190_ _02159_ _02193_ _02194_ VGND VGND VPWR VPWR _02195_ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21141_ net2073 _01156_ VGND VGND VPWR VPWR _01157_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21072_ _01083_ _01084_ _01087_ VGND VGND VPWR VPWR _01088_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2308 net2309 VGND VGND VPWR VPWR net2308 sky130_fd_sc_hd__buf_1
Xwire2319 net2320 VGND VGND VPWR VPWR net2319 sky130_fd_sc_hd__buf_1
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24900_ _04691_ VGND VGND VPWR VPWR _00743_ sky130_fd_sc_hd__clkbuf_1
X_20023_ _11800_ _11851_ _11852_ VGND VGND VPWR VPWR _11853_ sky130_fd_sc_hd__o21ai_1
X_25880_ clknet_leaf_15_clk _00753_ net8622 VGND VGND VPWR VPWR pid_q.ki\[8\] sky130_fd_sc_hd__dfrtp_1
Xwire1607 net1608 VGND VGND VPWR VPWR net1607 sky130_fd_sc_hd__clkbuf_1
Xwire1629 _04780_ VGND VGND VPWR VPWR net1629 sky130_fd_sc_hd__dlymetal6s2s_1
X_24831_ net5043 _04642_ net2000 net924 VGND VGND VPWR VPWR _00717_ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24762_ pid_q.curr_error\[8\] net1368 net1367 net690 VGND VGND VPWR VPWR _00705_
+ sky130_fd_sc_hd__a22o_1
X_21974_ _01860_ _01862_ _01958_ _01981_ VGND VGND VPWR VPWR _01982_ sky130_fd_sc_hd__a211o_1
Xmax_length7026 cordic0.vec\[1\]\[6\] VGND VGND VPWR VPWR net7026 sky130_fd_sc_hd__buf_1
X_23713_ _03577_ _03483_ _03578_ VGND VGND VPWR VPWR _03579_ sky130_fd_sc_hd__o21a_1
XFILLER_0_95_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20925_ net5527 net5905 VGND VGND VPWR VPWR _00941_ sky130_fd_sc_hd__nand2_1
X_24693_ net7490 VGND VGND VPWR VPWR _04531_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length7059 net7060 VGND VGND VPWR VPWR net7059 sky130_fd_sc_hd__clkbuf_1
X_23644_ _03410_ _03421_ _03510_ VGND VGND VPWR VPWR _03511_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_166_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20856_ net3840 VGND VGND VPWR VPWR _00872_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23575_ net2424 _03345_ _03442_ VGND VGND VPWR VPWR _03443_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_14_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20787_ _12555_ _12557_ VGND VGND VPWR VPWR _12558_ sky130_fd_sc_hd__xnor2_1
X_25314_ clknet_leaf_79_clk _00197_ net8490 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.e\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_22526_ pid_d.prev_error\[0\] net1699 _02525_ VGND VGND VPWR VPWR _00535_ sky130_fd_sc_hd__a21o_1
Xwire904 net905 VGND VGND VPWR VPWR net904 sky130_fd_sc_hd__buf_1
Xwire915 _05718_ VGND VGND VPWR VPWR net915 sky130_fd_sc_hd__buf_1
XFILLER_0_91_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire926 _04646_ VGND VGND VPWR VPWR net926 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire937 _03319_ VGND VGND VPWR VPWR net937 sky130_fd_sc_hd__clkbuf_1
X_25245_ clknet_leaf_87_clk _00128_ net8436 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.a\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire948 _01503_ VGND VGND VPWR VPWR net948 sky130_fd_sc_hd__clkbuf_2
X_22457_ _02411_ _02458_ VGND VGND VPWR VPWR _02459_ sky130_fd_sc_hd__xnor2_1
Xwire959 _11597_ VGND VGND VPWR VPWR net959 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_157_Right_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21408_ _01321_ _01323_ _01421_ VGND VGND VPWR VPWR _01422_ sky130_fd_sc_hd__o21a_1
X_25176_ clknet_leaf_54_clk _00065_ net8729 VGND VGND VPWR VPWR svm0.periodTop\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13190_ _05454_ _05462_ VGND VGND VPWR VPWR _05463_ sky130_fd_sc_hd__xnor2_1
X_22388_ _02263_ _02267_ VGND VGND VPWR VPWR _02391_ sky130_fd_sc_hd__nand2_1
Xwire4200 _06976_ VGND VGND VPWR VPWR net4200 sky130_fd_sc_hd__clkbuf_1
X_24127_ _03987_ _03988_ VGND VGND VPWR VPWR _03989_ sky130_fd_sc_hd__xnor2_1
Xwire4211 net4212 VGND VGND VPWR VPWR net4211 sky130_fd_sc_hd__buf_1
X_21339_ _01348_ _01352_ net5638 VGND VGND VPWR VPWR _01353_ sky130_fd_sc_hd__o21ai_1
Xwire4222 _06962_ VGND VGND VPWR VPWR net4222 sky130_fd_sc_hd__buf_1
Xwire4233 net4234 VGND VGND VPWR VPWR net4233 sky130_fd_sc_hd__buf_1
Xwire4244 net4246 VGND VGND VPWR VPWR net4244 sky130_fd_sc_hd__clkbuf_1
Xwire4255 _05347_ VGND VGND VPWR VPWR net4255 sky130_fd_sc_hd__buf_1
Xwire3510 net3513 VGND VGND VPWR VPWR net3510 sky130_fd_sc_hd__buf_1
X_24058_ _03824_ _03826_ _03803_ VGND VGND VPWR VPWR _03921_ sky130_fd_sc_hd__o21ba_1
Xwire4266 net4267 VGND VGND VPWR VPWR net4266 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3532 net3534 VGND VGND VPWR VPWR net3532 sky130_fd_sc_hd__buf_1
Xwire3543 _07048_ VGND VGND VPWR VPWR net3543 sky130_fd_sc_hd__clkbuf_1
Xwire4288 net4289 VGND VGND VPWR VPWR net4288 sky130_fd_sc_hd__clkbuf_1
Xwire3554 net3555 VGND VGND VPWR VPWR net3554 sky130_fd_sc_hd__buf_1
Xwire4299 net4300 VGND VGND VPWR VPWR net4299 sky130_fd_sc_hd__buf_1
X_23009_ _02877_ _02878_ VGND VGND VPWR VPWR _02879_ sky130_fd_sc_hd__xnor2_1
X_15900_ net2732 net2788 _07873_ VGND VGND VPWR VPWR _07969_ sky130_fd_sc_hd__and3_1
Xwire3565 net3566 VGND VGND VPWR VPWR net3565 sky130_fd_sc_hd__clkbuf_1
Xwire2831 net2832 VGND VGND VPWR VPWR net2831 sky130_fd_sc_hd__clkbuf_1
Xwire3576 _07026_ VGND VGND VPWR VPWR net3576 sky130_fd_sc_hd__dlymetal6s2s_1
X_16880_ net6216 net6172 net6504 VGND VGND VPWR VPWR _08844_ sky130_fd_sc_hd__mux2_1
Xwire2842 net2843 VGND VGND VPWR VPWR net2842 sky130_fd_sc_hd__buf_1
Xwire3587 net3588 VGND VGND VPWR VPWR net3587 sky130_fd_sc_hd__buf_1
XFILLER_0_21_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3598 _06973_ VGND VGND VPWR VPWR net3598 sky130_fd_sc_hd__buf_1
Xwire2853 net2854 VGND VGND VPWR VPWR net2853 sky130_fd_sc_hd__buf_1
Xwire2864 _06829_ VGND VGND VPWR VPWR net2864 sky130_fd_sc_hd__clkbuf_1
X_15831_ net2223 _07900_ VGND VGND VPWR VPWR _07901_ sky130_fd_sc_hd__nor2_1
XFILLER_0_189_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18550_ net607 _10398_ _10339_ _10332_ VGND VGND VPWR VPWR _10399_ sky130_fd_sc_hd__a2bb2o_1
X_12974_ _05242_ _05184_ _05185_ VGND VGND VPWR VPWR _05247_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_32_Left_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15762_ net1536 _07756_ _07749_ VGND VGND VPWR VPWR _07832_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_188_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17501_ svm0.delta\[10\] _09388_ VGND VGND VPWR VPWR _09389_ sky130_fd_sc_hd__xnor2_1
X_14713_ net9130 net2861 net2263 net1288 VGND VGND VPWR VPWR _00147_ sky130_fd_sc_hd__a22o_1
X_18481_ net874 _10330_ VGND VGND VPWR VPWR _10331_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_86_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15693_ net2694 _07763_ VGND VGND VPWR VPWR _07764_ sky130_fd_sc_hd__nor2_1
X_17432_ svm0.delta\[15\] _09329_ VGND VGND VPWR VPWR _09331_ sky130_fd_sc_hd__or2_1
X_14644_ net8959 net2880 _06806_ VGND VGND VPWR VPWR _00126_ sky130_fd_sc_hd__a21o_1
XFILLER_0_170_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17363_ _09275_ VGND VGND VPWR VPWR _00376_ sky130_fd_sc_hd__clkbuf_1
X_14575_ net2389 _06737_ _06730_ VGND VGND VPWR VPWR _06751_ sky130_fd_sc_hd__a21oi_1
Xmax_length6881 net6882 VGND VGND VPWR VPWR net6881 sky130_fd_sc_hd__buf_1
XFILLER_0_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19102_ net6147 net6101 VGND VGND VPWR VPWR _10939_ sky130_fd_sc_hd__xnor2_2
X_16314_ _08359_ _08373_ _08375_ _08376_ VGND VGND VPWR VPWR _08377_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_165_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13526_ _05791_ _05796_ VGND VGND VPWR VPWR _05797_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17294_ net7828 _09207_ VGND VGND VPWR VPWR _09208_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19033_ net6105 VGND VGND VPWR VPWR _10870_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout6041 net6047 VGND VGND VPWR VPWR net6041 sky130_fd_sc_hd__buf_1
X_13457_ net1598 VGND VGND VPWR VPWR _05730_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16245_ _08267_ _08293_ _08289_ VGND VGND VPWR VPWR _08309_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_82_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_41_Left_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_124_Right_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout6063 net6076 VGND VGND VPWR VPWR net6063 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6096 net6100 VGND VGND VPWR VPWR net6096 sky130_fd_sc_hd__buf_1
X_13388_ _05405_ _05481_ VGND VGND VPWR VPWR _05661_ sky130_fd_sc_hd__xnor2_1
X_16176_ net385 _08238_ net424 VGND VGND VPWR VPWR _08241_ sky130_fd_sc_hd__o21a_1
XFILLER_0_50_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6191 net6193 VGND VGND VPWR VPWR net6191 sky130_fd_sc_hd__clkbuf_1
X_15127_ net1893 net1892 _07200_ VGND VGND VPWR VPWR _07201_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19935_ net1409 _11766_ VGND VGND VPWR VPWR _11767_ sky130_fd_sc_hd__xor2_1
X_15058_ net6547 net6592 net7389 VGND VGND VPWR VPWR _07132_ sky130_fd_sc_hd__o21a_1
XFILLER_0_195_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14009_ _06214_ _06271_ _06272_ VGND VGND VPWR VPWR _06273_ sky130_fd_sc_hd__a21oi_1
X_19866_ net3130 net6033 net2501 VGND VGND VPWR VPWR _11699_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18817_ _10654_ VGND VGND VPWR VPWR _10660_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_50_Left_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19797_ _11627_ _11629_ _11630_ VGND VGND VPWR VPWR _11631_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_179_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18748_ net1065 _10592_ VGND VGND VPWR VPWR _10593_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_76_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18679_ net3231 net2131 VGND VGND VPWR VPWR _10525_ sky130_fd_sc_hd__nor2_1
X_20710_ net6051 _12475_ VGND VGND VPWR VPWR _12483_ sky130_fd_sc_hd__nor2_1
X_21690_ _01591_ _01593_ _01589_ VGND VGND VPWR VPWR _01701_ sky130_fd_sc_hd__o21a_1
XFILLER_0_176_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20641_ _08992_ _12419_ VGND VGND VPWR VPWR _12420_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7809 net7810 VGND VGND VPWR VPWR net7809 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23360_ _03200_ _03229_ VGND VGND VPWR VPWR _03230_ sky130_fd_sc_hd__xnor2_1
X_20572_ net1742 _12355_ VGND VGND VPWR VPWR _12356_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22311_ _02152_ net1706 _02314_ VGND VGND VPWR VPWR _02315_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23291_ _02984_ _02987_ VGND VGND VPWR VPWR _03161_ sky130_fd_sc_hd__or2b_1
XFILLER_0_6_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25030_ net3739 net1157 VGND VGND VPWR VPWR _04783_ sky130_fd_sc_hd__xnor2_1
X_22242_ _02118_ _02166_ _02246_ VGND VGND VPWR VPWR _02247_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22173_ _02176_ _02177_ VGND VGND VPWR VPWR _02179_ sky130_fd_sc_hd__or2_1
X_21124_ _01133_ _01139_ VGND VGND VPWR VPWR _01140_ sky130_fd_sc_hd__xnor2_1
Xwire2105 _11378_ VGND VGND VPWR VPWR net2105 sky130_fd_sc_hd__clkbuf_1
Xwire2116 _10887_ VGND VGND VPWR VPWR net2116 sky130_fd_sc_hd__clkbuf_1
X_25932_ clknet_leaf_25_clk _00805_ net8579 VGND VGND VPWR VPWR pid_d.prev_int\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire2127 _10481_ VGND VGND VPWR VPWR net2127 sky130_fd_sc_hd__clkbuf_2
X_21055_ net3823 _01001_ _01060_ VGND VGND VPWR VPWR _01071_ sky130_fd_sc_hd__a21oi_1
Xwire2138 _10112_ VGND VGND VPWR VPWR net2138 sky130_fd_sc_hd__buf_1
Xwire2149 net2150 VGND VGND VPWR VPWR net2149 sky130_fd_sc_hd__clkbuf_1
Xwire1404 net1405 VGND VGND VPWR VPWR net1404 sky130_fd_sc_hd__clkbuf_2
Xwire1415 _11510_ VGND VGND VPWR VPWR net1415 sky130_fd_sc_hd__buf_1
Xwire1426 _11007_ VGND VGND VPWR VPWR net1426 sky130_fd_sc_hd__buf_1
X_20006_ _11782_ _11822_ VGND VGND VPWR VPWR _11836_ sky130_fd_sc_hd__nor2_1
X_25863_ clknet_leaf_15_clk _00736_ net8617 VGND VGND VPWR VPWR pid_q.mult0.a\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1437 net1438 VGND VGND VPWR VPWR net1437 sky130_fd_sc_hd__buf_1
Xwire1448 _09628_ VGND VGND VPWR VPWR net1448 sky130_fd_sc_hd__buf_1
Xwire1459 _09509_ VGND VGND VPWR VPWR net1459 sky130_fd_sc_hd__clkbuf_1
X_24814_ net5189 _04635_ _04636_ VGND VGND VPWR VPWR _04637_ sky130_fd_sc_hd__mux2_1
X_25794_ clknet_leaf_33_clk _00667_ net8681 VGND VGND VPWR VPWR pid_q.curr_int\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_24745_ pid_q.curr_error\[6\] net1371 net1366 net738 VGND VGND VPWR VPWR _00703_
+ sky130_fd_sc_hd__a22o_1
X_21957_ net3780 _01964_ VGND VGND VPWR VPWR _01965_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20908_ net5492 net5883 _00867_ _00923_ VGND VGND VPWR VPWR _00924_ sky130_fd_sc_hd__a31oi_2
X_24676_ net9133 _04508_ _04520_ VGND VGND VPWR VPWR _00690_ sky130_fd_sc_hd__a21o_1
X_12690_ net5263 _04856_ net4277 _04889_ svm0.vC\[6\] VGND VGND VPWR VPWR _04963_
+ sky130_fd_sc_hd__a32oi_1
XFILLER_0_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21888_ _01795_ _01895_ VGND VGND VPWR VPWR _01897_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length5410 net5411 VGND VGND VPWR VPWR net5410 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23627_ _03426_ _03427_ VGND VGND VPWR VPWR _03494_ sky130_fd_sc_hd__nand2_1
Xmax_length5432 net5433 VGND VGND VPWR VPWR net5432 sky130_fd_sc_hd__buf_1
X_20839_ _00853_ _00854_ VGND VGND VPWR VPWR _00855_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_182_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length6188 net6189 VGND VGND VPWR VPWR net6188 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14360_ _06571_ matmul0.a_in\[9\] net901 VGND VGND VPWR VPWR _06573_ sky130_fd_sc_hd__mux2_1
X_23558_ net4677 net4900 VGND VGND VPWR VPWR _03426_ sky130_fd_sc_hd__nand2_1
Xmax_length5487 net5488 VGND VGND VPWR VPWR net5487 sky130_fd_sc_hd__buf_1
Xwire701 _01630_ VGND VGND VPWR VPWR net701 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire712 _11252_ VGND VGND VPWR VPWR net712 sky130_fd_sc_hd__clkbuf_1
X_13311_ net7705 net1352 VGND VGND VPWR VPWR _05584_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire723 _08435_ VGND VGND VPWR VPWR net723 sky130_fd_sc_hd__dlymetal6s2s_1
X_22509_ _02451_ _02450_ _02452_ VGND VGND VPWR VPWR _02510_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire734 _05397_ VGND VGND VPWR VPWR net734 sky130_fd_sc_hd__buf_1
Xinput19 currA_in[11] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
Xwire745 net746 VGND VGND VPWR VPWR net745 sky130_fd_sc_hd__clkbuf_2
X_14291_ net80 _06518_ _06519_ net7724 VGND VGND VPWR VPWR _00060_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23489_ net4768 net4826 VGND VGND VPWR VPWR _03358_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire756 _02204_ VGND VGND VPWR VPWR net756 sky130_fd_sc_hd__buf_1
Xwire767 _10256_ VGND VGND VPWR VPWR net767 sky130_fd_sc_hd__clkbuf_1
X_13242_ _05509_ _05514_ VGND VGND VPWR VPWR _05515_ sky130_fd_sc_hd__xnor2_2
Xwire778 _07646_ VGND VGND VPWR VPWR net778 sky130_fd_sc_hd__buf_1
X_16030_ _08095_ _08096_ VGND VGND VPWR VPWR _08097_ sky130_fd_sc_hd__xnor2_1
Xwire789 _05225_ VGND VGND VPWR VPWR net789 sky130_fd_sc_hd__buf_1
X_25228_ clknet_leaf_66_clk _00117_ net8647 VGND VGND VPWR VPWR cordic_done sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25159_ clknet_leaf_45_clk _00048_ net8781 VGND VGND VPWR VPWR pid_q.target\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13173_ net1137 net1136 _05445_ VGND VGND VPWR VPWR _05446_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4030 _09215_ VGND VGND VPWR VPWR net4030 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_20_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17981_ net1214 net1447 _09827_ VGND VGND VPWR VPWR _09832_ sky130_fd_sc_hd__a21o_1
Xwire4063 net4064 VGND VGND VPWR VPWR net4063 sky130_fd_sc_hd__buf_1
Xwire4074 _07602_ VGND VGND VPWR VPWR net4074 sky130_fd_sc_hd__buf_1
X_19720_ net604 _11554_ VGND VGND VPWR VPWR _11555_ sky130_fd_sc_hd__nand2_1
Xwire4085 _07514_ VGND VGND VPWR VPWR net4085 sky130_fd_sc_hd__clkbuf_1
Xwire3351 net3352 VGND VGND VPWR VPWR net3351 sky130_fd_sc_hd__buf_1
X_16932_ net6374 VGND VGND VPWR VPWR _08896_ sky130_fd_sc_hd__inv_2
Xwire4096 net4097 VGND VGND VPWR VPWR net4096 sky130_fd_sc_hd__clkbuf_2
Xwire3362 _08843_ VGND VGND VPWR VPWR net3362 sky130_fd_sc_hd__buf_1
Xwire3373 net3374 VGND VGND VPWR VPWR net3373 sky130_fd_sc_hd__clkbuf_2
Xwire3384 net3385 VGND VGND VPWR VPWR net3384 sky130_fd_sc_hd__buf_1
XFILLER_0_165_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2650 _07763_ VGND VGND VPWR VPWR net2650 sky130_fd_sc_hd__buf_1
X_19651_ net1191 _11472_ _11478_ VGND VGND VPWR VPWR _11487_ sky130_fd_sc_hd__a21bo_1
Xwire2661 net2662 VGND VGND VPWR VPWR net2661 sky130_fd_sc_hd__buf_1
X_16863_ net6172 net6133 net6504 VGND VGND VPWR VPWR _08828_ sky130_fd_sc_hd__mux2_1
Xwire2672 net2673 VGND VGND VPWR VPWR net2672 sky130_fd_sc_hd__buf_1
Xwire2683 net2684 VGND VGND VPWR VPWR net2683 sky130_fd_sc_hd__buf_1
Xwire2694 _07505_ VGND VGND VPWR VPWR net2694 sky130_fd_sc_hd__buf_1
X_18602_ _10442_ _10449_ VGND VGND VPWR VPWR _10450_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1960 _04976_ VGND VGND VPWR VPWR net1960 sky130_fd_sc_hd__buf_1
X_15814_ _07879_ _07880_ _07883_ VGND VGND VPWR VPWR _07884_ sky130_fd_sc_hd__a21o_1
Xwire1971 _04926_ VGND VGND VPWR VPWR net1971 sky130_fd_sc_hd__buf_1
X_19582_ _11373_ _11418_ VGND VGND VPWR VPWR _11419_ sky130_fd_sc_hd__xnor2_1
X_16794_ cordic0.cos\[0\] matmul0.cos\[0\] net3370 VGND VGND VPWR VPWR _08787_ sky130_fd_sc_hd__mux2_1
Xwire1982 net1983 VGND VGND VPWR VPWR net1982 sky130_fd_sc_hd__buf_1
Xwire1993 _04853_ VGND VGND VPWR VPWR net1993 sky130_fd_sc_hd__clkbuf_2
X_18533_ net1766 net1440 _10381_ VGND VGND VPWR VPWR _10382_ sky130_fd_sc_hd__o21ai_1
X_15745_ _07814_ _07815_ VGND VGND VPWR VPWR _07816_ sky130_fd_sc_hd__nor2_1
X_12957_ _04982_ _05229_ _05216_ _05217_ net3689 VGND VGND VPWR VPWR _05230_ sky130_fd_sc_hd__o2111a_1
X_18464_ net3284 net3925 VGND VGND VPWR VPWR _10314_ sky130_fd_sc_hd__xnor2_1
X_15676_ net2699 _07601_ net4071 _07746_ VGND VGND VPWR VPWR _07747_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_169_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12888_ _05104_ _05105_ VGND VGND VPWR VPWR _05161_ sky130_fd_sc_hd__or2_1
Xmax_length7390 matmul0.matmul_stage_inst.e\[9\] VGND VGND VPWR VPWR net7390 sky130_fd_sc_hd__clkbuf_1
X_17415_ net611 _09317_ _09315_ VGND VGND VPWR VPWR _09318_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14627_ matmul0.start _06536_ _06649_ net6453 VGND VGND VPWR VPWR _06796_ sky130_fd_sc_hd__a22o_1
X_18395_ _10164_ _10179_ _10168_ VGND VGND VPWR VPWR _10246_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_23_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17346_ net6703 net7682 VGND VGND VPWR VPWR _09260_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14558_ _06730_ _06735_ VGND VGND VPWR VPWR _06736_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13509_ net2374 net324 net1127 net9152 VGND VGND VPWR VPWR _00017_ sky130_fd_sc_hd__a22o_1
X_17277_ net2983 net155 net2158 net9131 VGND VGND VPWR VPWR _00371_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14489_ _06667_ _06669_ _06672_ VGND VGND VPWR VPWR _06673_ sky130_fd_sc_hd__o21ai_2
X_19016_ net6209 net6248 VGND VGND VPWR VPWR _10853_ sky130_fd_sc_hd__or2b_1
XFILLER_0_141_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16228_ net1091 _08290_ net1085 VGND VGND VPWR VPWR _08293_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_3_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16159_ _08140_ net1256 net1517 VGND VGND VPWR VPWR _08225_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19918_ net3149 _11686_ VGND VGND VPWR VPWR _11750_ sky130_fd_sc_hd__and2_1
XFILLER_0_177_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19849_ net2506 _11639_ _11681_ VGND VGND VPWR VPWR _11682_ sky130_fd_sc_hd__a21oi_1
X_22860_ net8897 _02757_ VGND VGND VPWR VPWR _02758_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21811_ _01818_ _01738_ _01819_ VGND VGND VPWR VPWR _01820_ sky130_fd_sc_hd__o21a_1
X_22791_ _02703_ VGND VGND VPWR VPWR _00622_ sky130_fd_sc_hd__clkbuf_1
X_24530_ net328 _04385_ VGND VGND VPWR VPWR _04387_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21742_ _01750_ _01751_ VGND VGND VPWR VPWR _01752_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_176_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24461_ _04267_ _04318_ VGND VGND VPWR VPWR _04319_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_171_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21673_ _01680_ _01683_ VGND VGND VPWR VPWR _01684_ sky130_fd_sc_hd__xnor2_1
Xwire8307 net8308 VGND VGND VPWR VPWR net8307 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8318 net17 VGND VGND VPWR VPWR net8318 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length4016 _09257_ VGND VGND VPWR VPWR net4016 sky130_fd_sc_hd__buf_1
XFILLER_0_11_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8329 net8331 VGND VGND VPWR VPWR net8329 sky130_fd_sc_hd__buf_1
X_23412_ _03207_ _03212_ _03281_ VGND VGND VPWR VPWR _03282_ sky130_fd_sc_hd__a21o_1
XFILLER_0_163_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20624_ _12403_ _12404_ net6173 VGND VGND VPWR VPWR _12405_ sky130_fd_sc_hd__mux2_1
Xwire7606 net7607 VGND VGND VPWR VPWR net7606 sky130_fd_sc_hd__buf_1
X_24392_ pid_q.curr_error\[10\] VGND VGND VPWR VPWR _04251_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7617 net7618 VGND VGND VPWR VPWR net7617 sky130_fd_sc_hd__buf_1
XFILLER_0_190_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7639 net7640 VGND VGND VPWR VPWR net7639 sky130_fd_sc_hd__clkbuf_1
Xmax_length3326 net3327 VGND VGND VPWR VPWR net3326 sky130_fd_sc_hd__buf_1
X_23343_ _03207_ _03212_ VGND VGND VPWR VPWR _03213_ sky130_fd_sc_hd__xnor2_1
X_20555_ net2600 net3852 net3849 _08970_ _08971_ VGND VGND VPWR VPWR _12340_ sky130_fd_sc_hd__a221o_1
Xwire6916 net6914 VGND VGND VPWR VPWR net6916 sky130_fd_sc_hd__buf_1
XFILLER_0_11_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6927 net6928 VGND VGND VPWR VPWR net6927 sky130_fd_sc_hd__buf_1
Xwire6938 net6936 VGND VGND VPWR VPWR net6938 sky130_fd_sc_hd__buf_1
Xwire6949 net6950 VGND VGND VPWR VPWR net6949 sky130_fd_sc_hd__clkbuf_1
X_23274_ _03130_ _03139_ VGND VGND VPWR VPWR _03144_ sky130_fd_sc_hd__nor2_1
X_20486_ net6853 net6824 net6840 net6790 net6491 net6521 VGND VGND VPWR VPWR _12274_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_89_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25013_ net5179 _04762_ _04767_ VGND VGND VPWR VPWR _04768_ sky130_fd_sc_hd__o21ai_2
X_22225_ net5762 _02227_ _02229_ net3778 VGND VGND VPWR VPWR _02230_ sky130_fd_sc_hd__a211o_1
XFILLER_0_120_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22156_ _02059_ VGND VGND VPWR VPWR _02162_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21107_ net5584 net5880 VGND VGND VPWR VPWR _01123_ sky130_fd_sc_hd__nand2_1
XFILLER_0_196_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22087_ _01986_ _01996_ _01991_ VGND VGND VPWR VPWR _02094_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1201 net1204 VGND VGND VPWR VPWR net1201 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21038_ net5929 net5911 VGND VGND VPWR VPWR _01054_ sky130_fd_sc_hd__or2_1
X_25915_ clknet_leaf_27_clk _00788_ net8648 VGND VGND VPWR VPWR pid_q.out\[11\] sky130_fd_sc_hd__dfrtp_1
Xwire1212 _10007_ VGND VGND VPWR VPWR net1212 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1223 net1224 VGND VGND VPWR VPWR net1223 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_156_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1234 net1235 VGND VGND VPWR VPWR net1234 sky130_fd_sc_hd__buf_1
XFILLER_0_191_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1245 _08509_ VGND VGND VPWR VPWR net1245 sky130_fd_sc_hd__clkbuf_1
Xwire1256 _08145_ VGND VGND VPWR VPWR net1256 sky130_fd_sc_hd__buf_1
X_13860_ net841 _06048_ VGND VGND VPWR VPWR _06127_ sky130_fd_sc_hd__nor2_1
X_25846_ clknet_leaf_20_clk _00719_ net8616 VGND VGND VPWR VPWR pid_q.mult0.b\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1267 _07706_ VGND VGND VPWR VPWR net1267 sky130_fd_sc_hd__clkbuf_1
Xwire1278 net1279 VGND VGND VPWR VPWR net1278 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_69_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1289 _06854_ VGND VGND VPWR VPWR net1289 sky130_fd_sc_hd__clkbuf_1
X_12811_ _05079_ _05083_ VGND VGND VPWR VPWR _05084_ sky130_fd_sc_hd__and2_1
X_13791_ _06057_ _06058_ VGND VGND VPWR VPWR _06059_ sky130_fd_sc_hd__nand2_1
X_22989_ _02862_ VGND VGND VPWR VPWR _00661_ sky130_fd_sc_hd__clkbuf_1
X_25777_ clknet_leaf_81_clk _00650_ net8496 VGND VGND VPWR VPWR matmul0.beta_pass\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_106_Left_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15530_ net4075 net4074 VGND VGND VPWR VPWR _07603_ sky130_fd_sc_hd__nor2_1
X_24728_ pid_q.curr_error\[4\] net1368 net1365 _04561_ VGND VGND VPWR VPWR _00701_
+ sky130_fd_sc_hd__a22o_1
X_12742_ _05014_ VGND VGND VPWR VPWR _05015_ sky130_fd_sc_hd__buf_1
XFILLER_0_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8702 net8731 VGND VGND VPWR VPWR net8702 sky130_fd_sc_hd__buf_1
XFILLER_0_97_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12673_ net7836 net1346 VGND VGND VPWR VPWR _04946_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15461_ net2848 net2820 net2686 net2827 VGND VGND VPWR VPWR _07535_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24659_ net5168 _00011_ net1374 VGND VGND VPWR VPWR _04512_ sky130_fd_sc_hd__and3_1
X_17200_ net617 _09149_ net6841 VGND VGND VPWR VPWR _09150_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_127_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14412_ net8141 net3634 VGND VGND VPWR VPWR _06613_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8830 net8831 VGND VGND VPWR VPWR net8830 sky130_fd_sc_hd__clkbuf_1
X_18180_ net3340 net7142 VGND VGND VPWR VPWR _10031_ sky130_fd_sc_hd__nor2_1
Xwire8841 net8842 VGND VGND VPWR VPWR net8841 sky130_fd_sc_hd__clkbuf_1
X_15392_ _07435_ net779 _07458_ _07461_ _07465_ VGND VGND VPWR VPWR _07466_ sky130_fd_sc_hd__o32ai_1
Xwire8852 net8853 VGND VGND VPWR VPWR net8852 sky130_fd_sc_hd__clkbuf_1
Xwire8863 net8865 VGND VGND VPWR VPWR net8863 sky130_fd_sc_hd__buf_1
XFILLER_0_182_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8874 net8876 VGND VGND VPWR VPWR net8874 sky130_fd_sc_hd__buf_1
X_17131_ _09083_ _09085_ VGND VGND VPWR VPWR _09086_ sky130_fd_sc_hd__xnor2_2
Xwire520 net521 VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14343_ _06559_ VGND VGND VPWR VPWR _00072_ sky130_fd_sc_hd__clkbuf_1
Xwire8885 net128 VGND VGND VPWR VPWR net8885 sky130_fd_sc_hd__clkbuf_1
Xwire531 _06077_ VGND VGND VPWR VPWR net531 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire542 _03384_ VGND VGND VPWR VPWR net542 sky130_fd_sc_hd__clkbuf_1
Xwire553 net554 VGND VGND VPWR VPWR net553 sky130_fd_sc_hd__clkbuf_1
Xmax_length3860 net3861 VGND VGND VPWR VPWR net3860 sky130_fd_sc_hd__buf_1
Xwire564 net565 VGND VGND VPWR VPWR net564 sky130_fd_sc_hd__clkbuf_1
X_14274_ net50 net2914 _06517_ net9078 VGND VGND VPWR VPWR _00045_ sky130_fd_sc_hd__a22o_1
X_17062_ net7039 _09014_ _09016_ _09020_ VGND VGND VPWR VPWR _09021_ sky130_fd_sc_hd__a211o_1
XFILLER_0_40_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire575 net576 VGND VGND VPWR VPWR net575 sky130_fd_sc_hd__clkbuf_1
Xwire586 _04652_ VGND VGND VPWR VPWR net586 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire597 net598 VGND VGND VPWR VPWR net597 sky130_fd_sc_hd__clkbuf_1
X_13225_ _05496_ _05497_ VGND VGND VPWR VPWR _05498_ sky130_fd_sc_hd__xor2_1
XFILLER_0_21_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16013_ _08077_ _08080_ VGND VGND VPWR VPWR _08081_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_115_Left_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13156_ _05426_ _05427_ net917 VGND VGND VPWR VPWR _05429_ sky130_fd_sc_hd__a21o_1
XFILLER_0_176_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13087_ _05357_ net1001 VGND VGND VPWR VPWR _05360_ sky130_fd_sc_hd__xnor2_1
X_17964_ _09690_ net3990 _09813_ _09814_ VGND VGND VPWR VPWR _09815_ sky130_fd_sc_hd__o31a_1
XFILLER_0_100_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3170 net3171 VGND VGND VPWR VPWR net3170 sky130_fd_sc_hd__buf_1
X_19703_ net3291 _11411_ net3864 VGND VGND VPWR VPWR _11539_ sky130_fd_sc_hd__or3_1
Xwire3181 net3182 VGND VGND VPWR VPWR net3181 sky130_fd_sc_hd__clkbuf_1
X_16915_ net6370 net6399 VGND VGND VPWR VPWR _08879_ sky130_fd_sc_hd__or2b_1
Xwire3192 _10919_ VGND VGND VPWR VPWR net3192 sky130_fd_sc_hd__buf_1
X_17895_ _09093_ _09738_ net3242 VGND VGND VPWR VPWR _09746_ sky130_fd_sc_hd__o21ai_1
Xwire2480 _01052_ VGND VGND VPWR VPWR net2480 sky130_fd_sc_hd__buf_1
X_19634_ _11443_ _11470_ VGND VGND VPWR VPWR _11471_ sky130_fd_sc_hd__xor2_1
Xwire2491 _12299_ VGND VGND VPWR VPWR net2491 sky130_fd_sc_hd__clkbuf_1
X_16846_ net6421 matmul0.sin\[11\] net4287 VGND VGND VPWR VPWR _08814_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1790 _09583_ VGND VGND VPWR VPWR net1790 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_124_Left_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19565_ _11400_ _11401_ VGND VGND VPWR VPWR _11402_ sky130_fd_sc_hd__xnor2_1
X_16777_ net7600 matmul0.a\[8\] _08770_ VGND VGND VPWR VPWR _08778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13989_ net7743 net1570 VGND VGND VPWR VPWR _06254_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18516_ _10171_ _10364_ VGND VGND VPWR VPWR _10365_ sky130_fd_sc_hd__xor2_1
X_15728_ net887 _07798_ VGND VGND VPWR VPWR _07799_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19496_ net3168 net3897 VGND VGND VPWR VPWR _11333_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18447_ net6998 _10241_ VGND VGND VPWR VPWR _10297_ sky130_fd_sc_hd__nand2_1
X_15659_ net988 _07729_ VGND VGND VPWR VPWR _07731_ sky130_fd_sc_hd__or2_1
XFILLER_0_173_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18378_ _10225_ net2541 VGND VGND VPWR VPWR _10229_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_173_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17329_ svm0.counter\[3\] VGND VGND VPWR VPWR _09243_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_133_Left_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20340_ cordic0.slte0.opA\[4\] net1400 VGND VGND VPWR VPWR _12143_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20271_ _12080_ cordic0.slte0.opB\[15\] net2531 VGND VGND VPWR VPWR _12081_ sky130_fd_sc_hd__mux2_1
X_22010_ net5977 VGND VGND VPWR VPWR _02017_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23961_ _03700_ net1659 net1660 VGND VGND VPWR VPWR _03825_ sky130_fd_sc_hd__a21bo_1
X_25700_ clknet_leaf_120_clk _00573_ net8414 VGND VGND VPWR VPWR pid_d.mult0.b\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_22912_ _02802_ _02803_ VGND VGND VPWR VPWR _02804_ sky130_fd_sc_hd__nand2_1
X_23892_ _03748_ _03756_ VGND VGND VPWR VPWR _03757_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_169_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25631_ clknet_leaf_106_clk _00504_ net8353 VGND VGND VPWR VPWR cordic0.vec\[0\]\[3\]
+ sky130_fd_sc_hd__dfstp_1
X_22843_ net8897 _02742_ VGND VGND VPWR VPWR _02743_ sky130_fd_sc_hd__and2_1
XFILLER_0_190_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22774_ net8108 net3764 net2434 VGND VGND VPWR VPWR _02694_ sky130_fd_sc_hd__o21ai_1
X_25562_ clknet_leaf_64_clk _00435_ net8670 VGND VGND VPWR VPWR state\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24513_ _04279_ _04307_ _04369_ VGND VGND VPWR VPWR _04370_ sky130_fd_sc_hd__a21o_1
X_21725_ pid_d.curr_int\[5\] net3123 net2078 _01735_ VGND VGND VPWR VPWR _00524_ sky130_fd_sc_hd__a22o_1
X_25493_ clknet_leaf_48_clk _00373_ net8762 VGND VGND VPWR VPWR svm0.tA\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8104 net87 VGND VGND VPWR VPWR net8104 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8115 net8116 VGND VGND VPWR VPWR net8115 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8126 net48 VGND VGND VPWR VPWR net8126 sky130_fd_sc_hd__clkbuf_1
X_24444_ net4565 net4808 _04301_ VGND VGND VPWR VPWR _04302_ sky130_fd_sc_hd__and3_1
X_21656_ net5704 net5550 VGND VGND VPWR VPWR _01667_ sky130_fd_sc_hd__nand2_1
Xwire8137 net8138 VGND VGND VPWR VPWR net8137 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7403 matmul0.matmul_stage_inst.a\[14\] VGND VGND VPWR VPWR net7403 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8148 net8149 VGND VGND VPWR VPWR net8148 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7414 net7415 VGND VGND VPWR VPWR net7414 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8159 net8160 VGND VGND VPWR VPWR net8159 sky130_fd_sc_hd__clkbuf_1
Xfanout6618 net6622 VGND VGND VPWR VPWR net6618 sky130_fd_sc_hd__clkbuf_1
X_20607_ net6195 _12386_ _12387_ _12367_ VGND VGND VPWR VPWR _12388_ sky130_fd_sc_hd__o22a_1
Xwire7425 net7426 VGND VGND VPWR VPWR net7425 sky130_fd_sc_hd__clkbuf_1
X_24375_ net4603 net3044 _04154_ VGND VGND VPWR VPWR _04234_ sky130_fd_sc_hd__or3b_1
XFILLER_0_163_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21587_ _01489_ _01493_ _01598_ VGND VGND VPWR VPWR _01599_ sky130_fd_sc_hd__o21a_1
Xmax_length3134 _11489_ VGND VGND VPWR VPWR net3134 sky130_fd_sc_hd__buf_1
Xwire6713 svm0.counter\[8\] VGND VGND VPWR VPWR net6713 sky130_fd_sc_hd__clkbuf_1
Xmax_length3145 net3146 VGND VGND VPWR VPWR net3145 sky130_fd_sc_hd__buf_1
Xfanout5917 net5925 VGND VGND VPWR VPWR net5917 sky130_fd_sc_hd__clkbuf_1
Xwire6724 net6718 VGND VGND VPWR VPWR net6724 sky130_fd_sc_hd__buf_1
Xwire7469 pid_q.state\[5\] VGND VGND VPWR VPWR net7469 sky130_fd_sc_hd__clkbuf_1
X_23326_ _03190_ _03195_ VGND VGND VPWR VPWR _03196_ sky130_fd_sc_hd__xnor2_1
Xfanout5928 net5933 VGND VGND VPWR VPWR net5928 sky130_fd_sc_hd__buf_1
Xwire6735 svm0.counter\[2\] VGND VGND VPWR VPWR net6735 sky130_fd_sc_hd__buf_1
X_20538_ net1479 _12310_ net6326 VGND VGND VPWR VPWR _12323_ sky130_fd_sc_hd__a21o_1
Xwire6746 svm0.tA\[9\] VGND VGND VPWR VPWR net6746 sky130_fd_sc_hd__buf_1
XFILLER_0_15_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire6757 net6755 VGND VGND VPWR VPWR net6757 sky130_fd_sc_hd__buf_1
XFILLER_0_162_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6768 net6765 VGND VGND VPWR VPWR net6768 sky130_fd_sc_hd__buf_1
XFILLER_0_120_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6779 net6777 VGND VGND VPWR VPWR net6779 sky130_fd_sc_hd__buf_2
X_23257_ _03121_ _03122_ _03123_ VGND VGND VPWR VPWR _03127_ sky130_fd_sc_hd__and3_1
XFILLER_0_162_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20469_ cordic0.slte0.opA\[16\] net1810 _12259_ VGND VGND VPWR VPWR _12260_ sky130_fd_sc_hd__and3_1
XFILLER_0_160_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13010_ _05166_ _05167_ _05281_ _05282_ VGND VGND VPWR VPWR _05283_ sky130_fd_sc_hd__o211a_1
X_22208_ _02211_ _02212_ VGND VGND VPWR VPWR _02213_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23188_ net5116 net4719 VGND VGND VPWR VPWR _03058_ sky130_fd_sc_hd__nand2_1
Xmax_length1787 _09597_ VGND VGND VPWR VPWR net1787 sky130_fd_sc_hd__clkbuf_1
X_22139_ _02139_ _02144_ VGND VGND VPWR VPWR _02145_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_55_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14961_ _07029_ net4132 _07013_ net4151 VGND VGND VPWR VPWR _07035_ sky130_fd_sc_hd__o22a_1
Xwire1020 net1021 VGND VGND VPWR VPWR net1020 sky130_fd_sc_hd__buf_1
Xhold8 matmul0.matmul_stage_inst.a\[5\] VGND VGND VPWR VPWR net8961 sky130_fd_sc_hd__dlygate4sd3_1
Xwire1031 _02986_ VGND VGND VPWR VPWR net1031 sky130_fd_sc_hd__clkbuf_2
X_16700_ _08728_ _08724_ matmul0.matmul_stage_inst.mult2\[11\] VGND VGND VPWR VPWR
+ _08729_ sky130_fd_sc_hd__o21ba_1
X_13912_ _06117_ net1311 net1583 VGND VGND VPWR VPWR _06178_ sky130_fd_sc_hd__and3_1
Xwire1042 net1043 VGND VGND VPWR VPWR net1042 sky130_fd_sc_hd__clkbuf_1
X_17680_ _09543_ _09557_ _09558_ _09559_ VGND VGND VPWR VPWR _09560_ sky130_fd_sc_hd__a22o_1
Xwire1053 _12292_ VGND VGND VPWR VPWR net1053 sky130_fd_sc_hd__buf_1
XFILLER_0_96_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1064 _11011_ VGND VGND VPWR VPWR net1064 sky130_fd_sc_hd__buf_1
X_14892_ net6611 matmul0.matmul_stage_inst.b\[11\] matmul0.matmul_stage_inst.a\[11\]
+ net6581 VGND VGND VPWR VPWR _06966_ sky130_fd_sc_hd__a22o_1
Xwire1075 _10086_ VGND VGND VPWR VPWR net1075 sky130_fd_sc_hd__clkbuf_1
Xwire1086 net1087 VGND VGND VPWR VPWR net1086 sky130_fd_sc_hd__dlymetal6s2s_1
X_16631_ matmul0.alpha_pass\[2\] net2613 net6552 VGND VGND VPWR VPWR _08670_ sky130_fd_sc_hd__mux2_1
X_13843_ _06039_ _06033_ _06034_ VGND VGND VPWR VPWR _06110_ sky130_fd_sc_hd__a21bo_1
X_25829_ clknet_leaf_36_clk _00702_ net8752 VGND VGND VPWR VPWR pid_q.curr_error\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1097 net1098 VGND VGND VPWR VPWR net1097 sky130_fd_sc_hd__buf_1
XFILLER_0_18_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19350_ _11138_ VGND VGND VPWR VPWR _11187_ sky130_fd_sc_hd__inv_2
X_16562_ _08618_ _08620_ VGND VGND VPWR VPWR _08621_ sky130_fd_sc_hd__xnor2_1
X_13774_ _06040_ _06041_ VGND VGND VPWR VPWR _06042_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18301_ _10138_ _10148_ _10150_ _10151_ VGND VGND VPWR VPWR _10152_ sky130_fd_sc_hd__o211a_1
X_15513_ net1861 net1860 VGND VGND VPWR VPWR _07586_ sky130_fd_sc_hd__nor2_1
Xfanout8510 net8525 VGND VGND VPWR VPWR net8510 sky130_fd_sc_hd__buf_1
X_12725_ net1611 _04979_ _04994_ _04997_ VGND VGND VPWR VPWR _04998_ sky130_fd_sc_hd__nand4_1
X_19281_ _11106_ _11108_ net763 VGND VGND VPWR VPWR _11118_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_139_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16493_ net1084 net1078 _08551_ _08552_ VGND VGND VPWR VPWR _08553_ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8554 net8560 VGND VGND VPWR VPWR net8554 sky130_fd_sc_hd__clkbuf_2
X_18232_ _10038_ _10051_ _10052_ net7141 VGND VGND VPWR VPWR _10083_ sky130_fd_sc_hd__a31o_1
XFILLER_0_155_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout7820 net7843 VGND VGND VPWR VPWR net7820 sky130_fd_sc_hd__clkbuf_1
X_15444_ net3597 net3591 net4216 net4214 VGND VGND VPWR VPWR _07518_ sky130_fd_sc_hd__o22a_1
X_12656_ net3693 net4266 VGND VGND VPWR VPWR _04929_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8660 net8658 VGND VGND VPWR VPWR net8660 sky130_fd_sc_hd__buf_1
X_18163_ net1212 _10001_ VGND VGND VPWR VPWR _10014_ sky130_fd_sc_hd__xnor2_1
X_12587_ net8864 net7521 VGND VGND VPWR VPWR _04871_ sky130_fd_sc_hd__and2_1
X_15375_ _07437_ _07447_ VGND VGND VPWR VPWR _07449_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8693 net8694 VGND VGND VPWR VPWR net8693 sky130_fd_sc_hd__buf_1
X_17114_ net3362 _08847_ net2593 VGND VGND VPWR VPWR _09070_ sky130_fd_sc_hd__mux2_1
X_14326_ _06546_ matmul0.a_in\[1\] net902 VGND VGND VPWR VPWR _06547_ sky130_fd_sc_hd__mux2_1
Xwire7970 net7971 VGND VGND VPWR VPWR net7970 sky130_fd_sc_hd__clkbuf_1
X_18094_ _09932_ _09938_ VGND VGND VPWR VPWR _09945_ sky130_fd_sc_hd__and2_1
Xwire361 net362 VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__clkbuf_1
Xwire7981 net7982 VGND VGND VPWR VPWR net7981 sky130_fd_sc_hd__clkbuf_1
Xwire372 net373 VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__buf_1
Xwire7992 net7993 VGND VGND VPWR VPWR net7992 sky130_fd_sc_hd__clkbuf_1
Xwire383 net384 VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17045_ net3334 VGND VGND VPWR VPWR _09004_ sky130_fd_sc_hd__buf_1
Xwire394 net395 VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__clkbuf_1
X_14257_ net3658 VGND VGND VPWR VPWR _06511_ sky130_fd_sc_hd__buf_1
XFILLER_0_123_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13208_ _05471_ _05480_ VGND VGND VPWR VPWR _05481_ sky130_fd_sc_hd__xnor2_1
X_14188_ _06445_ _06447_ VGND VGND VPWR VPWR _06448_ sky130_fd_sc_hd__xor2_1
XFILLER_0_195_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13139_ net7873 net1947 VGND VGND VPWR VPWR _05412_ sky130_fd_sc_hd__nand2_1
X_18996_ net2528 _10832_ VGND VGND VPWR VPWR _10833_ sky130_fd_sc_hd__nand2_1
X_17947_ net6978 net6951 VGND VGND VPWR VPWR _09798_ sky130_fd_sc_hd__nand2_1
X_17878_ net6908 net6948 VGND VGND VPWR VPWR _09729_ sky130_fd_sc_hd__nand2_1
X_19617_ net6087 _11379_ _11452_ _11376_ _11453_ VGND VGND VPWR VPWR _11454_ sky130_fd_sc_hd__a221o_1
X_16829_ _08805_ VGND VGND VPWR VPWR _00312_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19548_ _10944_ _10975_ VGND VGND VPWR VPWR _11385_ sky130_fd_sc_hd__or2b_1
XFILLER_0_75_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19479_ _11308_ _11309_ _11312_ _10986_ _11315_ VGND VGND VPWR VPWR _11316_ sky130_fd_sc_hd__a221o_1
XFILLER_0_159_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21510_ net806 net757 VGND VGND VPWR VPWR _01523_ sky130_fd_sc_hd__and2_1
X_22490_ _02419_ _02424_ _02427_ VGND VGND VPWR VPWR _02491_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_118_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21441_ _01349_ _01354_ _01453_ VGND VGND VPWR VPWR _01454_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_173_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6009 net6010 VGND VGND VPWR VPWR net6009 sky130_fd_sc_hd__buf_1
XFILLER_0_90_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24160_ net694 _04021_ VGND VGND VPWR VPWR _04022_ sky130_fd_sc_hd__xnor2_2
X_21372_ _01377_ _01385_ VGND VGND VPWR VPWR _01386_ sky130_fd_sc_hd__xnor2_1
Xwire5308 net5309 VGND VGND VPWR VPWR net5308 sky130_fd_sc_hd__buf_1
XFILLER_0_71_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5319 pid_d.out\[15\] VGND VGND VPWR VPWR net5319 sky130_fd_sc_hd__clkbuf_1
X_23111_ _02979_ _02980_ VGND VGND VPWR VPWR _02981_ sky130_fd_sc_hd__xnor2_2
X_20323_ net951 _12125_ VGND VGND VPWR VPWR _12127_ sky130_fd_sc_hd__nand2_1
X_24091_ net5178 net3063 net2029 _03953_ VGND VGND VPWR VPWR _00672_ sky130_fd_sc_hd__a22o_1
Xwire4607 net4608 VGND VGND VPWR VPWR net4607 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4618 net4609 VGND VGND VPWR VPWR net4618 sky130_fd_sc_hd__buf_1
XFILLER_0_12_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23042_ _02909_ _02910_ _02911_ VGND VGND VPWR VPWR _02912_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20254_ _12067_ cordic0.slte0.opB\[11\] net2531 VGND VGND VPWR VPWR _12068_ sky130_fd_sc_hd__mux2_1
Xwire3906 _10801_ VGND VGND VPWR VPWR net3906 sky130_fd_sc_hd__buf_1
Xwire3917 _10787_ VGND VGND VPWR VPWR net3917 sky130_fd_sc_hd__buf_1
Xwire3928 net3929 VGND VGND VPWR VPWR net3928 sky130_fd_sc_hd__buf_1
X_20185_ net6004 _11648_ _12006_ _12008_ _12005_ VGND VGND VPWR VPWR _12011_ sky130_fd_sc_hd__a311o_1
X_24993_ _04751_ VGND VGND VPWR VPWR _00776_ sky130_fd_sc_hd__clkbuf_1
X_23944_ net4518 net4986 VGND VGND VPWR VPWR _03808_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23875_ _03617_ _03618_ _03616_ VGND VGND VPWR VPWR _03740_ sky130_fd_sc_hd__a21o_1
Xmax_length8668 net8664 VGND VGND VPWR VPWR net8668 sky130_fd_sc_hd__buf_1
X_25614_ clknet_leaf_108_clk _00487_ net8351 VGND VGND VPWR VPWR cordic0.slte0.opA\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_196_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22826_ net5366 net5984 VGND VGND VPWR VPWR _02727_ sky130_fd_sc_hd__nand2_1
XFILLER_0_168_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25545_ clknet_leaf_28_clk _00425_ net8652 VGND VGND VPWR VPWR pid_q.prev_int\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22757_ pid_d.ki\[10\] net3069 net2037 VGND VGND VPWR VPWR _02683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13490_ net1130 _05643_ VGND VGND VPWR VPWR _05763_ sky130_fd_sc_hd__or2b_1
X_21708_ _01612_ _01613_ _01605_ VGND VGND VPWR VPWR _01719_ sky130_fd_sc_hd__a21bo_1
X_25476_ clknet_leaf_48_clk _00356_ net8762 VGND VGND VPWR VPWR svm0.tB\[14\] sky130_fd_sc_hd__dfrtp_1
X_22688_ _02633_ net5548 net2447 VGND VGND VPWR VPWR _02634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7200 net7202 VGND VGND VPWR VPWR net7200 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24427_ _04206_ _04211_ _04204_ VGND VGND VPWR VPWR _04285_ sky130_fd_sc_hd__o21a_1
Xwire7222 net7223 VGND VGND VPWR VPWR net7222 sky130_fd_sc_hd__clkbuf_1
X_21639_ _01554_ _01615_ VGND VGND VPWR VPWR _01650_ sky130_fd_sc_hd__nand2_1
Xwire7233 net7234 VGND VGND VPWR VPWR net7233 sky130_fd_sc_hd__buf_1
Xwire7244 net7245 VGND VGND VPWR VPWR net7244 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_23_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire7255 net7259 VGND VGND VPWR VPWR net7255 sky130_fd_sc_hd__clkbuf_1
Xwire6510 net6511 VGND VGND VPWR VPWR net6510 sky130_fd_sc_hd__buf_1
Xwire7266 net7267 VGND VGND VPWR VPWR net7266 sky130_fd_sc_hd__clkbuf_1
X_15160_ _07223_ net1884 _07233_ VGND VGND VPWR VPWR _07234_ sky130_fd_sc_hd__o21a_1
X_24358_ net4994 _04214_ _04215_ _04216_ VGND VGND VPWR VPWR _04217_ sky130_fd_sc_hd__o211a_1
Xwire7277 matmul0.alpha_pass\[8\] VGND VGND VPWR VPWR net7277 sky130_fd_sc_hd__clkbuf_1
Xwire6532 net6533 VGND VGND VPWR VPWR net6532 sky130_fd_sc_hd__buf_1
Xwire7288 net7289 VGND VGND VPWR VPWR net7288 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length2241 _07275_ VGND VGND VPWR VPWR net2241 sky130_fd_sc_hd__clkbuf_1
Xwire6554 net6562 VGND VGND VPWR VPWR net6554 sky130_fd_sc_hd__clkbuf_1
X_14111_ _06341_ _06343_ _06372_ VGND VGND VPWR VPWR _06373_ sky130_fd_sc_hd__o21ai_1
Xfanout5758 net5766 VGND VGND VPWR VPWR net5758 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7299 net7300 VGND VGND VPWR VPWR net7299 sky130_fd_sc_hd__buf_1
X_23309_ _03006_ VGND VGND VPWR VPWR _03179_ sky130_fd_sc_hd__inv_2
X_15091_ _07124_ _07164_ VGND VGND VPWR VPWR _07165_ sky130_fd_sc_hd__xnor2_1
Xwire6565 net6566 VGND VGND VPWR VPWR net6565 sky130_fd_sc_hd__clkbuf_1
Xwire5820 net5821 VGND VGND VPWR VPWR net5820 sky130_fd_sc_hd__buf_1
X_24289_ net3041 _04148_ VGND VGND VPWR VPWR _04149_ sky130_fd_sc_hd__xnor2_1
Xmax_length2263 _06825_ VGND VGND VPWR VPWR net2263 sky130_fd_sc_hd__buf_1
Xwire6576 net6577 VGND VGND VPWR VPWR net6576 sky130_fd_sc_hd__clkbuf_1
Xwire5831 net5832 VGND VGND VPWR VPWR net5831 sky130_fd_sc_hd__buf_1
Xwire5842 net5843 VGND VGND VPWR VPWR net5842 sky130_fd_sc_hd__buf_1
Xwire6587 net6588 VGND VGND VPWR VPWR net6587 sky130_fd_sc_hd__buf_1
Xwire6598 net6599 VGND VGND VPWR VPWR net6598 sky130_fd_sc_hd__clkbuf_1
Xwire5853 net5854 VGND VGND VPWR VPWR net5853 sky130_fd_sc_hd__buf_1
Xwire5864 net5865 VGND VGND VPWR VPWR net5864 sky130_fd_sc_hd__buf_1
X_14042_ _06227_ _06232_ _06224_ VGND VGND VPWR VPWR _06306_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_31_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5875 net5876 VGND VGND VPWR VPWR net5875 sky130_fd_sc_hd__clkbuf_1
Xwire5886 net5887 VGND VGND VPWR VPWR net5886 sky130_fd_sc_hd__clkbuf_1
Xwire5897 net5898 VGND VGND VPWR VPWR net5897 sky130_fd_sc_hd__buf_1
X_18850_ _10664_ _10665_ net658 VGND VGND VPWR VPWR _10693_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17801_ net3255 net3258 net3266 _09651_ net7061 VGND VGND VPWR VPWR _09652_ sky130_fd_sc_hd__a311o_1
X_18781_ net526 _10624_ _10602_ VGND VGND VPWR VPWR _10625_ sky130_fd_sc_hd__o21ai_1
X_15993_ _08037_ net883 VGND VGND VPWR VPWR _08061_ sky130_fd_sc_hd__and2_1
X_17732_ net2590 _09588_ VGND VGND VPWR VPWR _09589_ sky130_fd_sc_hd__nor2_1
X_14944_ net6634 net6582 net7404 VGND VGND VPWR VPWR _07018_ sky130_fd_sc_hd__o21a_1
XFILLER_0_173_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17663_ net4007 svm0.tA\[7\] _09542_ VGND VGND VPWR VPWR _09543_ sky130_fd_sc_hd__a21boi_1
X_14875_ _06955_ VGND VGND VPWR VPWR _00208_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19402_ net1192 _11229_ net1061 VGND VGND VPWR VPWR _11239_ sky130_fd_sc_hd__a21o_1
XFILLER_0_159_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16614_ matmul0.matmul_stage_inst.mult2\[14\] net167 net3467 VGND VGND VPWR VPWR
+ _08657_ sky130_fd_sc_hd__mux2_1
X_13826_ net7669 net2308 net1953 VGND VGND VPWR VPWR _06093_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17594_ net4030 svm0.tB\[15\] svm0.tB\[13\] _09426_ _09474_ VGND VGND VPWR VPWR _09475_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_97_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19333_ net6352 net2525 VGND VGND VPWR VPWR _11170_ sky130_fd_sc_hd__and2_1
XFILLER_0_175_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16545_ net2638 _08603_ VGND VGND VPWR VPWR _08604_ sky130_fd_sc_hd__nand2_1
X_13757_ _05939_ _05940_ VGND VGND VPWR VPWR _06025_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12708_ net7826 net2338 net1968 VGND VGND VPWR VPWR _04981_ sky130_fd_sc_hd__and3_2
X_19264_ _11100_ _10893_ VGND VGND VPWR VPWR _11101_ sky130_fd_sc_hd__xnor2_1
X_16476_ _08534_ net671 VGND VGND VPWR VPWR _08537_ sky130_fd_sc_hd__or2b_1
X_13688_ _05878_ _05955_ _05956_ VGND VGND VPWR VPWR _05957_ sky130_fd_sc_hd__a21o_1
Xfanout8362 net8369 VGND VGND VPWR VPWR net8362 sky130_fd_sc_hd__buf_1
X_18215_ _09176_ _10065_ VGND VGND VPWR VPWR _10066_ sky130_fd_sc_hd__xnor2_1
X_15427_ net1273 _07500_ VGND VGND VPWR VPWR _07501_ sky130_fd_sc_hd__xnor2_1
X_12639_ svm0.vC\[3\] net2990 net3694 net4269 VGND VGND VPWR VPWR _04912_ sky130_fd_sc_hd__a22oi_1
X_19195_ _10899_ _11031_ VGND VGND VPWR VPWR _11032_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_170_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18146_ _09872_ net2549 _09873_ _09958_ VGND VGND VPWR VPWR _09997_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_41_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8490 net8491 VGND VGND VPWR VPWR net8490 sky130_fd_sc_hd__buf_1
XFILLER_0_124_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15358_ net1116 _07430_ VGND VGND VPWR VPWR _07432_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14309_ net6450 _06513_ VGND VGND VPWR VPWR _06531_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6993 net7001 VGND VGND VPWR VPWR net6993 sky130_fd_sc_hd__clkbuf_1
Xwire180 _10616_ VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold205 matmul0.a_in\[3\] VGND VGND VPWR VPWR net9158 sky130_fd_sc_hd__dlygate4sd3_1
Xwire191 net192 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__buf_1
X_18077_ _09905_ _09924_ _09925_ _09927_ VGND VGND VPWR VPWR _09928_ sky130_fd_sc_hd__o31a_1
Xhold216 pid_d.curr_int\[10\] VGND VGND VPWR VPWR net9169 sky130_fd_sc_hd__dlygate4sd3_1
X_15289_ _07360_ _07361_ net2794 net2790 _07362_ VGND VGND VPWR VPWR _07363_ sky130_fd_sc_hd__o2111ai_1
Xhold227 svm0.tC\[5\] VGND VGND VPWR VPWR net9180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 cordic0.slte0.opA\[14\] VGND VGND VPWR VPWR net9191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 pid_q.curr_int\[10\] VGND VGND VPWR VPWR net9202 sky130_fd_sc_hd__dlygate4sd3_1
X_17028_ net3362 _08845_ _08987_ _08847_ net3335 net6480 VGND VGND VPWR VPWR _08988_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_22_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18979_ net3213 net3903 _10815_ net6291 VGND VGND VPWR VPWR _10816_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_147_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21990_ _01986_ _01997_ VGND VGND VPWR VPWR _01998_ sky130_fd_sc_hd__xnor2_1
X_20941_ _00900_ net2481 VGND VGND VPWR VPWR _00957_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23660_ net4576 net4998 VGND VGND VPWR VPWR _03527_ sky130_fd_sc_hd__nand2_1
X_20872_ _12541_ _00813_ VGND VGND VPWR VPWR _00888_ sky130_fd_sc_hd__xnor2_1
Xmax_length6518 net6519 VGND VGND VPWR VPWR net6518 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_72_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22611_ net7237 _02579_ VGND VGND VPWR VPWR _02584_ sky130_fd_sc_hd__xnor2_1
X_23591_ _03457_ _03458_ VGND VGND VPWR VPWR _03459_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_147_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_138_Right_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25330_ clknet_leaf_80_clk _00213_ net8488 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.f\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_22542_ net9119 net1701 _02533_ VGND VGND VPWR VPWR _00543_ sky130_fd_sc_hd__a21o_1
XFILLER_0_174_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22473_ net5689 _02472_ _02473_ VGND VGND VPWR VPWR _02474_ sky130_fd_sc_hd__and3_1
X_25261_ clknet_leaf_75_clk _00144_ net8458 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.b\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24212_ net1380 net1379 VGND VGND VPWR VPWR _04073_ sky130_fd_sc_hd__or2b_1
X_21424_ pid_d.prev_int\[2\] _01337_ _01338_ net5983 VGND VGND VPWR VPWR _01437_ sky130_fd_sc_hd__a31o_1
X_25192_ clknet_leaf_58_clk _00081_ net8721 VGND VGND VPWR VPWR matmul0.a_in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire5105 net5106 VGND VGND VPWR VPWR net5105 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5116 net5111 VGND VGND VPWR VPWR net5116 sky130_fd_sc_hd__clkbuf_2
X_24143_ _03892_ _03918_ _04004_ VGND VGND VPWR VPWR _04005_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21355_ _01366_ _01368_ VGND VGND VPWR VPWR _01369_ sky130_fd_sc_hd__xnor2_1
Xwire5138 net5127 VGND VGND VPWR VPWR net5138 sky130_fd_sc_hd__buf_1
XFILLER_0_130_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4404 net4405 VGND VGND VPWR VPWR net4404 sky130_fd_sc_hd__clkbuf_1
Xwire5149 net5155 VGND VGND VPWR VPWR net5149 sky130_fd_sc_hd__clkbuf_2
Xwire4415 net4416 VGND VGND VPWR VPWR net4415 sky130_fd_sc_hd__clkbuf_1
X_20306_ _09054_ _12098_ _12110_ net3313 net6459 VGND VGND VPWR VPWR _12111_ sky130_fd_sc_hd__a221o_1
X_24074_ net1161 _03833_ _03936_ VGND VGND VPWR VPWR _03937_ sky130_fd_sc_hd__o21ai_2
Xwire4426 net4427 VGND VGND VPWR VPWR net4426 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21286_ net1391 net1390 VGND VGND VPWR VPWR _01301_ sky130_fd_sc_hd__xor2_1
Xwire4437 net4438 VGND VGND VPWR VPWR net4437 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4448 net4449 VGND VGND VPWR VPWR net4448 sky130_fd_sc_hd__clkbuf_1
Xwire3703 net3704 VGND VGND VPWR VPWR net3703 sky130_fd_sc_hd__buf_1
Xwire3714 net3715 VGND VGND VPWR VPWR net3714 sky130_fd_sc_hd__clkbuf_1
Xwire4459 net4460 VGND VGND VPWR VPWR net4459 sky130_fd_sc_hd__clkbuf_1
X_23025_ net5015 net4693 VGND VGND VPWR VPWR _02895_ sky130_fd_sc_hd__nand2_1
Xwire3725 net3726 VGND VGND VPWR VPWR net3725 sky130_fd_sc_hd__clkbuf_1
X_20237_ net12 _12050_ VGND VGND VPWR VPWR _12054_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3747 _03456_ VGND VGND VPWR VPWR net3747 sky130_fd_sc_hd__buf_1
Xwire3769 net3770 VGND VGND VPWR VPWR net3769 sky130_fd_sc_hd__buf_1
X_20168_ _11927_ _11955_ _11993_ VGND VGND VPWR VPWR _11994_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_196_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24976_ pid_q.kp\[7\] _04716_ net1358 VGND VGND VPWR VPWR _04743_ sky130_fd_sc_hd__mux2_1
X_12990_ _05176_ _05181_ net1143 VGND VGND VPWR VPWR _05263_ sky130_fd_sc_hd__a21o_1
X_20099_ _11910_ _11920_ net420 _11911_ VGND VGND VPWR VPWR _11927_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_118_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23927_ _03789_ _03790_ VGND VGND VPWR VPWR _03791_ sky130_fd_sc_hd__xor2_2
XFILLER_0_19_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length8443 net8444 VGND VGND VPWR VPWR net8443 sky130_fd_sc_hd__buf_1
XFILLER_0_118_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length7720 net7721 VGND VGND VPWR VPWR net7720 sky130_fd_sc_hd__buf_1
X_14660_ net7446 net7168 net2873 VGND VGND VPWR VPWR _06815_ sky130_fd_sc_hd__and3_1
XFILLER_0_98_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23858_ _03622_ _03627_ _03620_ VGND VGND VPWR VPWR _03723_ sky130_fd_sc_hd__o21a_1
Xmax_length7742 net7743 VGND VGND VPWR VPWR net7742 sky130_fd_sc_hd__buf_1
Xmax_length8487 net8479 VGND VGND VPWR VPWR net8487 sky130_fd_sc_hd__clkbuf_1
Xmax_length8498 net8495 VGND VGND VPWR VPWR net8498 sky130_fd_sc_hd__clkbuf_2
Xmax_length7764 net7765 VGND VGND VPWR VPWR net7764 sky130_fd_sc_hd__clkbuf_1
X_13611_ _05879_ _05880_ VGND VGND VPWR VPWR _05881_ sky130_fd_sc_hd__nor2_1
X_22809_ net4328 pid_d.out_valid net3763 VGND VGND VPWR VPWR _02713_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14591_ net2887 _06764_ _06765_ net892 net8995 VGND VGND VPWR VPWR _00114_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_105_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23789_ _03653_ _03654_ VGND VGND VPWR VPWR _03655_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16330_ _08319_ _08320_ _08392_ VGND VGND VPWR VPWR _08393_ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25528_ clknet_leaf_45_clk net8963 net8791 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__dfrtp_1
X_13542_ _05809_ _05812_ VGND VGND VPWR VPWR _05813_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_138_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16261_ _08270_ _08272_ _08324_ VGND VGND VPWR VPWR _08325_ sky130_fd_sc_hd__a21o_1
X_13473_ net7671 net1982 net2360 VGND VGND VPWR VPWR _05746_ sky130_fd_sc_hd__and3_1
Xfanout6212 cordic0.vec\[0\]\[7\] VGND VGND VPWR VPWR net6212 sky130_fd_sc_hd__clkbuf_2
X_25459_ clknet_leaf_66_clk _00013_ net8662 VGND VGND VPWR VPWR matmul0.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout6223 net6228 VGND VGND VPWR VPWR net6223 sky130_fd_sc_hd__clkbuf_1
X_18000_ _08913_ _09617_ _09644_ _09849_ _09850_ VGND VGND VPWR VPWR _09851_ sky130_fd_sc_hd__a221o_1
Xwire7041 net7039 VGND VGND VPWR VPWR net7041 sky130_fd_sc_hd__buf_1
X_15212_ _07195_ _07284_ _07285_ VGND VGND VPWR VPWR _07286_ sky130_fd_sc_hd__o21a_1
Xwire7052 net7050 VGND VGND VPWR VPWR net7052 sky130_fd_sc_hd__buf_2
X_16192_ net2721 net2707 VGND VGND VPWR VPWR _08257_ sky130_fd_sc_hd__xnor2_1
Xwire7063 net7064 VGND VGND VPWR VPWR net7063 sky130_fd_sc_hd__buf_1
Xwire7074 net7079 VGND VGND VPWR VPWR net7074 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7085 net7080 VGND VGND VPWR VPWR net7085 sky130_fd_sc_hd__clkbuf_1
Xwire6340 net6337 VGND VGND VPWR VPWR net6340 sky130_fd_sc_hd__clkbuf_2
Xfanout4810 net4819 VGND VGND VPWR VPWR net4810 sky130_fd_sc_hd__buf_1
X_15143_ net991 _07215_ _07216_ _07212_ VGND VGND VPWR VPWR _07217_ sky130_fd_sc_hd__o211a_1
Xfanout4821 net4829 VGND VGND VPWR VPWR net4821 sky130_fd_sc_hd__buf_1
XFILLER_0_23_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6362 net6358 VGND VGND VPWR VPWR net6362 sky130_fd_sc_hd__buf_1
Xwire6373 cordic0.slte0.opA\[7\] VGND VGND VPWR VPWR net6373 sky130_fd_sc_hd__buf_1
XFILLER_0_168_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6384 net6385 VGND VGND VPWR VPWR net6384 sky130_fd_sc_hd__clkbuf_1
Xwire6395 cordic0.slte0.opB\[14\] VGND VGND VPWR VPWR net6395 sky130_fd_sc_hd__clkbuf_1
Xwire5661 net5662 VGND VGND VPWR VPWR net5661 sky130_fd_sc_hd__buf_1
X_15074_ net2251 net2790 net2789 _07147_ VGND VGND VPWR VPWR _07148_ sky130_fd_sc_hd__a31o_1
X_19951_ _11780_ _11781_ VGND VGND VPWR VPWR _11783_ sky130_fd_sc_hd__or2_1
Xwire5672 net5669 VGND VGND VPWR VPWR net5672 sky130_fd_sc_hd__buf_1
Xwire5683 net5684 VGND VGND VPWR VPWR net5683 sky130_fd_sc_hd__clkbuf_1
X_14025_ _06287_ _06288_ VGND VGND VPWR VPWR _06289_ sky130_fd_sc_hd__xor2_1
X_18902_ _10741_ _10742_ VGND VGND VPWR VPWR _10743_ sky130_fd_sc_hd__or2b_1
Xwire4960 net4961 VGND VGND VPWR VPWR net4960 sky130_fd_sc_hd__buf_1
Xwire4971 net4972 VGND VGND VPWR VPWR net4971 sky130_fd_sc_hd__buf_1
X_19882_ _11712_ _11714_ VGND VGND VPWR VPWR _11715_ sky130_fd_sc_hd__xor2_2
Xwire4982 net4984 VGND VGND VPWR VPWR net4982 sky130_fd_sc_hd__buf_1
XFILLER_0_140_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18833_ net3298 _10531_ _10675_ VGND VGND VPWR VPWR _10676_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_184_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18764_ _10501_ _10564_ VGND VGND VPWR VPWR _10609_ sky130_fd_sc_hd__and2_1
X_15976_ net2718 net3399 _07953_ VGND VGND VPWR VPWR _08044_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17715_ net9211 net1219 net1453 pid_q.curr_int\[6\] VGND VGND VPWR VPWR _00420_ sky130_fd_sc_hd__a22o_1
X_14927_ net4178 _06998_ net4177 _07000_ VGND VGND VPWR VPWR _07001_ sky130_fd_sc_hd__o22a_1
X_18695_ net6778 net1760 VGND VGND VPWR VPWR _10541_ sky130_fd_sc_hd__nand2_1
XFILLER_0_188_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17646_ net4026 svm0.tA\[8\] VGND VGND VPWR VPWR _09526_ sky130_fd_sc_hd__and2_1
XFILLER_0_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14858_ _06946_ VGND VGND VPWR VPWR _00200_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13809_ net621 _05990_ _06076_ VGND VGND VPWR VPWR _06077_ sky130_fd_sc_hd__a21o_1
XFILLER_0_129_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17577_ svm0.tC\[7\] _09430_ VGND VGND VPWR VPWR _09459_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_109_clk clknet_4_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_109_clk
+ sky130_fd_sc_hd__clkbuf_16
X_14789_ net9057 net3003 net992 VGND VGND VPWR VPWR _00167_ sky130_fd_sc_hd__o21a_1
X_19316_ _11152_ VGND VGND VPWR VPWR _11153_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16528_ _08550_ _08587_ VGND VGND VPWR VPWR _08588_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19247_ _11083_ net6240 _11056_ VGND VGND VPWR VPWR _11084_ sky130_fd_sc_hd__mux2_1
X_16459_ _08510_ _08519_ VGND VGND VPWR VPWR _08520_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_144_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19178_ _11014_ _10910_ net1757 VGND VGND VPWR VPWR _11015_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_170_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18129_ net3339 net3262 net3976 net7092 VGND VGND VPWR VPWR _09980_ sky130_fd_sc_hd__o211a_1
XFILLER_0_143_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21140_ _01126_ _01129_ VGND VGND VPWR VPWR _01156_ sky130_fd_sc_hd__xor2_2
X_21071_ _01083_ _01084_ _01086_ VGND VGND VPWR VPWR _01087_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2309 net2310 VGND VGND VPWR VPWR net2309 sky130_fd_sc_hd__buf_1
XFILLER_0_158_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20022_ net6081 net3199 _11797_ VGND VGND VPWR VPWR _11852_ sky130_fd_sc_hd__or3_1
XFILLER_0_10_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1608 net1609 VGND VGND VPWR VPWR net1608 sky130_fd_sc_hd__buf_1
Xwire1619 net1620 VGND VGND VPWR VPWR net1619 sky130_fd_sc_hd__buf_1
X_24830_ net7480 _04561_ net1383 VGND VGND VPWR VPWR _04648_ sky130_fd_sc_hd__a21o_1
X_24761_ _04588_ _04590_ VGND VGND VPWR VPWR _04591_ sky130_fd_sc_hd__xnor2_1
X_21973_ net1716 net1718 VGND VGND VPWR VPWR _01981_ sky130_fd_sc_hd__and2_1
X_23712_ pid_q.curr_int\[3\] VGND VGND VPWR VPWR _03578_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20924_ net5507 net5935 VGND VGND VPWR VPWR _00940_ sky130_fd_sc_hd__nand2_1
X_24692_ net1643 VGND VGND VPWR VPWR _04530_ sky130_fd_sc_hd__buf_1
Xmax_length7049 cordic0.vec\[1\]\[5\] VGND VGND VPWR VPWR net7049 sky130_fd_sc_hd__buf_1
XFILLER_0_96_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length6315 net6313 VGND VGND VPWR VPWR net6315 sky130_fd_sc_hd__buf_1
XFILLER_0_95_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length6326 net6324 VGND VGND VPWR VPWR net6326 sky130_fd_sc_hd__clkbuf_2
X_23643_ _03410_ _03421_ net1384 VGND VGND VPWR VPWR _03510_ sky130_fd_sc_hd__a21bo_1
X_20855_ net5879 VGND VGND VPWR VPWR _00871_ sky130_fd_sc_hd__inv_2
XFILLER_0_178_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4902 net4897 VGND VGND VPWR VPWR net4902 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23574_ net2424 _03345_ _03341_ VGND VGND VPWR VPWR _03442_ sky130_fd_sc_hd__a21bo_1
X_20786_ net5730 net5740 _12556_ VGND VGND VPWR VPWR _12557_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25313_ clknet_leaf_78_clk _00196_ net8511 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.e\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_22525_ net5973 net2379 net2046 VGND VGND VPWR VPWR _02525_ sky130_fd_sc_hd__and3_1
Xwire916 _05714_ VGND VGND VPWR VPWR net916 sky130_fd_sc_hd__buf_1
Xwire927 _04645_ VGND VGND VPWR VPWR net927 sky130_fd_sc_hd__clkbuf_1
Xwire938 _03303_ VGND VGND VPWR VPWR net938 sky130_fd_sc_hd__buf_1
XFILLER_0_45_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25244_ clknet_leaf_89_clk _00127_ net8443 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.a\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_22456_ _02456_ _02457_ VGND VGND VPWR VPWR _02458_ sky130_fd_sc_hd__nor2_1
Xwire949 net950 VGND VGND VPWR VPWR net949 sky130_fd_sc_hd__buf_1
XFILLER_0_122_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21407_ _01321_ _01323_ _01315_ VGND VGND VPWR VPWR _01421_ sky130_fd_sc_hd__a21bo_1
X_25175_ clknet_leaf_54_clk _00064_ net8730 VGND VGND VPWR VPWR svm0.periodTop\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_22387_ _02337_ _02389_ VGND VGND VPWR VPWR _02390_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4201 net4203 VGND VGND VPWR VPWR net4201 sky130_fd_sc_hd__buf_1
X_24126_ net4553 net4889 VGND VGND VPWR VPWR _03988_ sky130_fd_sc_hd__nand2_1
X_21338_ net5687 _01349_ VGND VGND VPWR VPWR _01352_ sky130_fd_sc_hd__nor2_1
Xwire4212 _06970_ VGND VGND VPWR VPWR net4212 sky130_fd_sc_hd__buf_1
XFILLER_0_102_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4223 _06826_ VGND VGND VPWR VPWR net4223 sky130_fd_sc_hd__clkbuf_1
Xwire4234 _06526_ VGND VGND VPWR VPWR net4234 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4245 net4246 VGND VGND VPWR VPWR net4245 sky130_fd_sc_hd__buf_1
Xwire3500 net3501 VGND VGND VPWR VPWR net3500 sky130_fd_sc_hd__clkbuf_1
Xwire4256 net4257 VGND VGND VPWR VPWR net4256 sky130_fd_sc_hd__buf_1
X_24057_ _03890_ _03919_ VGND VGND VPWR VPWR _03920_ sky130_fd_sc_hd__xnor2_1
Xwire3522 net3523 VGND VGND VPWR VPWR net3522 sky130_fd_sc_hd__buf_1
X_21269_ _00852_ _00853_ _01283_ VGND VGND VPWR VPWR _01284_ sky130_fd_sc_hd__a21oi_2
Xwire4278 _04893_ VGND VGND VPWR VPWR net4278 sky130_fd_sc_hd__buf_1
XFILLER_0_25_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3533 net3535 VGND VGND VPWR VPWR net3533 sky130_fd_sc_hd__clkbuf_1
Xwire3544 _07047_ VGND VGND VPWR VPWR net3544 sky130_fd_sc_hd__clkbuf_2
Xwire4289 net4290 VGND VGND VPWR VPWR net4289 sky130_fd_sc_hd__buf_1
X_23008_ net5133 net4595 VGND VGND VPWR VPWR _02878_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3566 net3567 VGND VGND VPWR VPWR net3566 sky130_fd_sc_hd__buf_1
Xwire2821 net2822 VGND VGND VPWR VPWR net2821 sky130_fd_sc_hd__clkbuf_1
Xwire2832 _07077_ VGND VGND VPWR VPWR net2832 sky130_fd_sc_hd__buf_1
Xwire2843 net2844 VGND VGND VPWR VPWR net2843 sky130_fd_sc_hd__clkbuf_1
Xwire3588 net3589 VGND VGND VPWR VPWR net3588 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire2854 _06914_ VGND VGND VPWR VPWR net2854 sky130_fd_sc_hd__dlymetal6s2s_1
X_15830_ net3425 net2695 VGND VGND VPWR VPWR _07900_ sky130_fd_sc_hd__nand2_1
Xwire3599 net3600 VGND VGND VPWR VPWR net3599 sky130_fd_sc_hd__buf_1
Xwire2865 _06824_ VGND VGND VPWR VPWR net2865 sky130_fd_sc_hd__clkbuf_2
Xwire2876 net2877 VGND VGND VPWR VPWR net2876 sky130_fd_sc_hd__buf_1
Xwire2887 net2888 VGND VGND VPWR VPWR net2887 sky130_fd_sc_hd__clkbuf_2
X_15761_ _07737_ _07827_ _07826_ VGND VGND VPWR VPWR _07831_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_63_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24959_ _04733_ VGND VGND VPWR VPWR _00760_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12973_ _05241_ net735 VGND VGND VPWR VPWR _05246_ sky130_fd_sc_hd__nand2_1
X_17500_ _09307_ _09383_ _09387_ VGND VGND VPWR VPWR _09388_ sky130_fd_sc_hd__a21o_1
X_14712_ matmul0.sin\[11\] _06853_ VGND VGND VPWR VPWR _06854_ sky130_fd_sc_hd__xnor2_1
X_18480_ _10328_ _10329_ VGND VGND VPWR VPWR _10330_ sky130_fd_sc_hd__nand2_1
X_15692_ net3556 VGND VGND VPWR VPWR _07763_ sky130_fd_sc_hd__buf_1
XFILLER_0_170_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17431_ net9213 _09329_ VGND VGND VPWR VPWR _09330_ sky130_fd_sc_hd__nand2_1
X_14643_ net7439 net7181 net2875 VGND VGND VPWR VPWR _06806_ sky130_fd_sc_hd__and3_1
XFILLER_0_185_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17362_ _09271_ _09274_ svm0.delta\[1\] VGND VGND VPWR VPWR _09275_ sky130_fd_sc_hd__mux2_1
Xmax_length6871 cordic0.vec\[1\]\[13\] VGND VGND VPWR VPWR net6871 sky130_fd_sc_hd__clkbuf_1
X_14574_ net2888 _06743_ _06750_ net894 net8967 VGND VGND VPWR VPWR _00112_ sky130_fd_sc_hd__a32o_1
X_19101_ net6162 _10937_ VGND VGND VPWR VPWR _10938_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16313_ net385 net493 net492 _08304_ VGND VGND VPWR VPWR _08376_ sky130_fd_sc_hd__and4b_1
X_13525_ _05792_ _05795_ VGND VGND VPWR VPWR _05796_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17293_ net7890 net7862 _09206_ VGND VGND VPWR VPWR _09207_ sky130_fd_sc_hd__or3_1
XFILLER_0_82_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19032_ _10867_ _10868_ VGND VGND VPWR VPWR _10869_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_153_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout6031 net6038 VGND VGND VPWR VPWR net6031 sky130_fd_sc_hd__buf_1
X_16244_ _08256_ _08295_ _08307_ VGND VGND VPWR VPWR _08308_ sky130_fd_sc_hd__a21o_1
X_13456_ _05727_ _05728_ VGND VGND VPWR VPWR _05729_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout6064 net6068 VGND VGND VPWR VPWR net6064 sky130_fd_sc_hd__clkbuf_1
X_16175_ _08231_ _08233_ _08239_ VGND VGND VPWR VPWR _08240_ sky130_fd_sc_hd__a21o_1
X_13387_ _05565_ _05566_ _05655_ _05659_ VGND VGND VPWR VPWR _05660_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5374 pid_d.mult0.a\[15\] VGND VGND VPWR VPWR net5374 sky130_fd_sc_hd__clkbuf_1
Xwire6170 net6171 VGND VGND VPWR VPWR net6170 sky130_fd_sc_hd__buf_1
XFILLER_0_105_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15126_ net1893 net1892 _07199_ VGND VGND VPWR VPWR _07200_ sky130_fd_sc_hd__a21o_1
Xfanout4673 net4686 VGND VGND VPWR VPWR net4673 sky130_fd_sc_hd__buf_1
X_19934_ _11764_ _11765_ VGND VGND VPWR VPWR _11766_ sky130_fd_sc_hd__and2_1
X_15057_ net6622 net6639 matmul0.matmul_stage_inst.f\[9\] VGND VGND VPWR VPWR _07131_
+ sky130_fd_sc_hd__o21a_1
Xwire5491 net5492 VGND VGND VPWR VPWR net5491 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_189_Left_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14008_ _06265_ _06268_ VGND VGND VPWR VPWR _06272_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4790 net4792 VGND VGND VPWR VPWR net4790 sky130_fd_sc_hd__clkbuf_1
X_19865_ net1412 _11697_ VGND VGND VPWR VPWR _11698_ sky130_fd_sc_hd__xnor2_2
X_18816_ net9098 net2288 net1449 _10659_ VGND VGND VPWR VPWR _00446_ sky130_fd_sc_hd__a31o_1
X_19796_ net6088 net3141 net6016 net2100 VGND VGND VPWR VPWR _11630_ sky130_fd_sc_hd__or4_1
XFILLER_0_37_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15959_ net3460 net2660 VGND VGND VPWR VPWR _08027_ sky130_fd_sc_hd__nor2_1
X_18747_ net1429 _10591_ VGND VGND VPWR VPWR _10592_ sky130_fd_sc_hd__xor2_1
X_18678_ net6893 net3231 net2131 _10523_ VGND VGND VPWR VPWR _10524_ sky130_fd_sc_hd__o31a_1
XFILLER_0_194_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17629_ net3279 svm0.tB\[11\] svm0.tB\[10\] _09393_ VGND VGND VPWR VPWR _09510_ sky130_fd_sc_hd__a31o_1
XFILLER_0_59_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20640_ net1395 _12397_ net1739 VGND VGND VPWR VPWR _12419_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20571_ net1745 _12342_ net1480 VGND VGND VPWR VPWR _12355_ sky130_fd_sc_hd__o21a_1
XFILLER_0_160_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3508 _07096_ VGND VGND VPWR VPWR net3508 sky130_fd_sc_hd__buf_1
XFILLER_0_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22310_ _02152_ net1706 net1712 VGND VGND VPWR VPWR _02314_ sky130_fd_sc_hd__o21a_1
X_23290_ _03145_ _03158_ _03159_ VGND VGND VPWR VPWR _03160_ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22241_ _02118_ _02166_ _02119_ VGND VGND VPWR VPWR _02246_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22172_ _02176_ _02177_ VGND VGND VPWR VPWR _02178_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21123_ _01092_ _01138_ VGND VGND VPWR VPWR _01139_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2106 _11378_ VGND VGND VPWR VPWR net2106 sky130_fd_sc_hd__clkbuf_2
X_25931_ clknet_leaf_26_clk _00804_ net8577 VGND VGND VPWR VPWR pid_d.prev_int\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire2117 net2118 VGND VGND VPWR VPWR net2117 sky130_fd_sc_hd__buf_1
X_21054_ _01060_ _01069_ VGND VGND VPWR VPWR _01070_ sky130_fd_sc_hd__and2b_1
Xwire2128 _10433_ VGND VGND VPWR VPWR net2128 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2139 net2140 VGND VGND VPWR VPWR net2139 sky130_fd_sc_hd__buf_1
Xwire1405 _11857_ VGND VGND VPWR VPWR net1405 sky130_fd_sc_hd__clkbuf_1
X_20005_ _11784_ _11824_ VGND VGND VPWR VPWR _11835_ sky130_fd_sc_hd__or2_1
Xwire1416 _11407_ VGND VGND VPWR VPWR net1416 sky130_fd_sc_hd__buf_1
X_25862_ clknet_leaf_14_clk _00735_ net8617 VGND VGND VPWR VPWR pid_q.mult0.a\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1427 _10759_ VGND VGND VPWR VPWR net1427 sky130_fd_sc_hd__clkbuf_1
Xwire1438 net1439 VGND VGND VPWR VPWR net1438 sky130_fd_sc_hd__buf_1
Xwire1449 _09598_ VGND VGND VPWR VPWR net1449 sky130_fd_sc_hd__buf_1
X_24813_ net7955 _04628_ VGND VGND VPWR VPWR _04636_ sky130_fd_sc_hd__nand2_1
X_25793_ clknet_leaf_32_clk _00666_ net8681 VGND VGND VPWR VPWR pid_q.curr_int\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_193_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24744_ net8002 _04575_ VGND VGND VPWR VPWR _04576_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_190_Right_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21956_ net5841 net5862 VGND VGND VPWR VPWR _01964_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20907_ net5491 _00922_ _00866_ VGND VGND VPWR VPWR _00923_ sky130_fd_sc_hd__a21oi_1
X_24675_ pid_q.curr_error\[9\] net3019 _04510_ VGND VGND VPWR VPWR _04520_ sky130_fd_sc_hd__and3_1
X_21887_ _01795_ _01895_ VGND VGND VPWR VPWR _01896_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23626_ _03489_ _03492_ VGND VGND VPWR VPWR _03493_ sky130_fd_sc_hd__xnor2_2
Xmax_length5433 net5434 VGND VGND VPWR VPWR net5433 sky130_fd_sc_hd__buf_1
X_20838_ net5702 net5626 VGND VGND VPWR VPWR _00854_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23557_ _03336_ _03347_ _03424_ VGND VGND VPWR VPWR _03425_ sky130_fd_sc_hd__o21a_1
XFILLER_0_181_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire702 _01521_ VGND VGND VPWR VPWR net702 sky130_fd_sc_hd__buf_1
X_20769_ _12537_ _12538_ _12539_ VGND VGND VPWR VPWR _12540_ sky130_fd_sc_hd__o21ai_1
Xwire713 _11118_ VGND VGND VPWR VPWR net713 sky130_fd_sc_hd__clkbuf_1
X_13310_ _05495_ _05496_ _05582_ VGND VGND VPWR VPWR _05583_ sky130_fd_sc_hd__o21ai_1
X_22508_ _02498_ _02508_ VGND VGND VPWR VPWR _02509_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire724 _08355_ VGND VGND VPWR VPWR net724 sky130_fd_sc_hd__buf_1
X_14290_ net79 net2901 net2264 net7734 VGND VGND VPWR VPWR _00059_ sky130_fd_sc_hd__a22o_1
Xwire746 net747 VGND VGND VPWR VPWR net746 sky130_fd_sc_hd__clkbuf_1
X_23488_ net4784 net4813 VGND VGND VPWR VPWR _03357_ sky130_fd_sc_hd__nand2_2
XFILLER_0_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire757 _01422_ VGND VGND VPWR VPWR net757 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire768 _10017_ VGND VGND VPWR VPWR net768 sky130_fd_sc_hd__clkbuf_1
X_13241_ _05511_ net1133 VGND VGND VPWR VPWR _05514_ sky130_fd_sc_hd__xor2_1
X_25227_ clknet_leaf_59_clk _00116_ net8694 VGND VGND VPWR VPWR svm0.vC\[15\] sky130_fd_sc_hd__dfrtp_1
X_22439_ net1712 _02152_ VGND VGND VPWR VPWR _02441_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire779 _07452_ VGND VGND VPWR VPWR net779 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25158_ clknet_leaf_54_clk _00047_ net8727 VGND VGND VPWR VPWR pid_q.target\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13172_ _05441_ _05444_ VGND VGND VPWR VPWR _05445_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4020 net4021 VGND VGND VPWR VPWR net4020 sky130_fd_sc_hd__buf_1
Xwire4031 _09215_ VGND VGND VPWR VPWR net4031 sky130_fd_sc_hd__buf_1
XFILLER_0_131_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24109_ _03969_ _03970_ net3742 VGND VGND VPWR VPWR _03971_ sky130_fd_sc_hd__a21oi_1
X_17980_ net3245 net1779 net1447 net1214 VGND VGND VPWR VPWR _09831_ sky130_fd_sc_hd__a211o_1
X_25089_ net4401 _04833_ VGND VGND VPWR VPWR _04834_ sky130_fd_sc_hd__nand2_1
Xwire4053 _08932_ VGND VGND VPWR VPWR net4053 sky130_fd_sc_hd__clkbuf_1
Xwire4064 net4065 VGND VGND VPWR VPWR net4064 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4075 net4076 VGND VGND VPWR VPWR net4075 sky130_fd_sc_hd__dlymetal6s2s_1
X_16931_ net6410 net6373 VGND VGND VPWR VPWR _08895_ sky130_fd_sc_hd__xnor2_1
Xwire4086 _07484_ VGND VGND VPWR VPWR net4086 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3352 net3353 VGND VGND VPWR VPWR net3352 sky130_fd_sc_hd__clkbuf_1
Xwire4097 _07144_ VGND VGND VPWR VPWR net4097 sky130_fd_sc_hd__clkbuf_1
Xwire3363 _08829_ VGND VGND VPWR VPWR net3363 sky130_fd_sc_hd__buf_1
Xwire3374 net3375 VGND VGND VPWR VPWR net3374 sky130_fd_sc_hd__clkbuf_1
Xwire3385 net3386 VGND VGND VPWR VPWR net3385 sky130_fd_sc_hd__clkbuf_1
X_16862_ net6167 net6123 net6501 VGND VGND VPWR VPWR _08827_ sky130_fd_sc_hd__mux2_1
Xwire2651 net2652 VGND VGND VPWR VPWR net2651 sky130_fd_sc_hd__clkbuf_2
X_19650_ net9049 net2122 net1444 _11486_ VGND VGND VPWR VPWR _00453_ sky130_fd_sc_hd__a31o_1
Xwire3396 _07686_ VGND VGND VPWR VPWR net3396 sky130_fd_sc_hd__buf_1
Xwire2662 net2663 VGND VGND VPWR VPWR net2662 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2673 net2674 VGND VGND VPWR VPWR net2673 sky130_fd_sc_hd__clkbuf_1
X_15813_ _07783_ _07881_ _07882_ VGND VGND VPWR VPWR _07883_ sky130_fd_sc_hd__a21o_1
Xwire2684 net2685 VGND VGND VPWR VPWR net2684 sky130_fd_sc_hd__clkbuf_1
X_18601_ _10444_ _10448_ net6831 VGND VGND VPWR VPWR _10449_ sky130_fd_sc_hd__mux2_1
Xwire1950 net1951 VGND VGND VPWR VPWR net1950 sky130_fd_sc_hd__buf_1
X_19581_ _11375_ _11417_ VGND VGND VPWR VPWR _11418_ sky130_fd_sc_hd__xor2_1
Xwire2695 net2696 VGND VGND VPWR VPWR net2695 sky130_fd_sc_hd__buf_1
X_16793_ _08786_ VGND VGND VPWR VPWR _00295_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1972 net1973 VGND VGND VPWR VPWR net1972 sky130_fd_sc_hd__buf_1
Xwire1983 net1984 VGND VGND VPWR VPWR net1983 sky130_fd_sc_hd__buf_1
XFILLER_0_172_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1994 _04787_ VGND VGND VPWR VPWR net1994 sky130_fd_sc_hd__dlymetal6s2s_1
X_18532_ net1766 net1440 net1207 VGND VGND VPWR VPWR _10381_ sky130_fd_sc_hd__a21o_1
X_15744_ net2758 _07812_ net1265 VGND VGND VPWR VPWR _07815_ sky130_fd_sc_hd__nor3_1
XFILLER_0_172_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12956_ net7889 net1350 VGND VGND VPWR VPWR _05229_ sky130_fd_sc_hd__nor2_1
XFILLER_0_181_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18463_ _10310_ _10311_ net6815 VGND VGND VPWR VPWR _10313_ sky130_fd_sc_hd__mux2_1
X_15675_ net2761 _07745_ VGND VGND VPWR VPWR _07746_ sky130_fd_sc_hd__nor2_1
X_12887_ net7906 net1958 _05104_ _05105_ VGND VGND VPWR VPWR _05160_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17414_ net3276 _09316_ VGND VGND VPWR VPWR _09317_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14626_ net6448 net6443 matmul0.start _06794_ VGND VGND VPWR VPWR _06795_ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18394_ net1774 _10244_ VGND VGND VPWR VPWR _10245_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17345_ net7702 _09211_ VGND VGND VPWR VPWR _09259_ sky130_fd_sc_hd__nand2_1
X_14557_ _06733_ _06734_ net1625 VGND VGND VPWR VPWR _06735_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_40_clk clknet_4_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_184_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13508_ net1308 VGND VGND VPWR VPWR _05780_ sky130_fd_sc_hd__clkbuf_1
X_17276_ net2981 net158 net2156 net9143 VGND VGND VPWR VPWR _00370_ sky130_fd_sc_hd__a22o_1
X_14488_ _06667_ _06669_ _06668_ VGND VGND VPWR VPWR _06672_ sky130_fd_sc_hd__a21o_1
X_19015_ _10849_ _10851_ VGND VGND VPWR VPWR _10852_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_141_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16227_ _08291_ VGND VGND VPWR VPWR _08292_ sky130_fd_sc_hd__clkbuf_1
X_13439_ _05707_ _05711_ VGND VGND VPWR VPWR _05712_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16158_ net672 _08223_ VGND VGND VPWR VPWR _08224_ sky130_fd_sc_hd__xor2_1
X_15109_ net1894 _07182_ VGND VGND VPWR VPWR _07183_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16089_ _08153_ _08155_ VGND VGND VPWR VPWR _08156_ sky130_fd_sc_hd__xor2_1
Xfanout4492 pid_q.mult0.a\[15\] VGND VGND VPWR VPWR net4492 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19917_ net3149 _11686_ VGND VGND VPWR VPWR _11749_ sky130_fd_sc_hd__nor2_1
XFILLER_0_177_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19848_ net6157 net2506 VGND VGND VPWR VPWR _11681_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19779_ _11542_ net604 VGND VGND VPWR VPWR _11613_ sky130_fd_sc_hd__nand2_1
X_21810_ net5979 VGND VGND VPWR VPWR _01819_ sky130_fd_sc_hd__inv_2
XFILLER_0_196_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22790_ pid_d.kp\[7\] _02676_ net1681 VGND VGND VPWR VPWR _02703_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21741_ net5567 net5679 VGND VGND VPWR VPWR _01751_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24460_ _04268_ _04317_ VGND VGND VPWR VPWR _04318_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21672_ net5769 net5505 _01681_ _01682_ VGND VGND VPWR VPWR _01683_ sky130_fd_sc_hd__a31o_1
XFILLER_0_114_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8308 net8309 VGND VGND VPWR VPWR net8308 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8319 net8320 VGND VGND VPWR VPWR net8319 sky130_fd_sc_hd__clkbuf_1
X_23411_ _03207_ _03212_ net2429 VGND VGND VPWR VPWR _03281_ sky130_fd_sc_hd__o21a_1
XFILLER_0_190_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20623_ net1494 _12402_ VGND VGND VPWR VPWR _12404_ sky130_fd_sc_hd__nand2_1
Xwire7607 net7609 VGND VGND VPWR VPWR net7607 sky130_fd_sc_hd__buf_1
X_24391_ _04197_ _04249_ VGND VGND VPWR VPWR _04250_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_31_clk clknet_4_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_191_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7618 net7619 VGND VGND VPWR VPWR net7618 sky130_fd_sc_hd__clkbuf_1
Xwire7629 net7631 VGND VGND VPWR VPWR net7629 sky130_fd_sc_hd__buf_1
XFILLER_0_61_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23342_ _03208_ _03211_ VGND VGND VPWR VPWR _03212_ sky130_fd_sc_hd__xnor2_2
X_20554_ net6480 _12338_ VGND VGND VPWR VPWR _12339_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6906 net6907 VGND VGND VPWR VPWR net6906 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6917 net6914 VGND VGND VPWR VPWR net6917 sky130_fd_sc_hd__buf_1
XFILLER_0_190_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length2626 _07936_ VGND VGND VPWR VPWR net2626 sky130_fd_sc_hd__buf_1
X_23273_ _03133_ _03142_ VGND VGND VPWR VPWR _03143_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20485_ net8057 net3170 _12272_ _12273_ VGND VGND VPWR VPWR _00501_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25012_ net5179 _04760_ _04761_ net4466 VGND VGND VPWR VPWR _04767_ sky130_fd_sc_hd__a31o_1
X_22224_ net5762 _02228_ VGND VGND VPWR VPWR _02229_ sky130_fd_sc_hd__nor2_1
X_22155_ net1710 _02057_ VGND VGND VPWR VPWR _02161_ sky130_fd_sc_hd__and2_1
X_21106_ net5605 net5880 _01121_ VGND VGND VPWR VPWR _01122_ sky130_fd_sc_hd__and3_1
X_22086_ _02081_ _02092_ VGND VGND VPWR VPWR _02093_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_196_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_98_clk clknet_4_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_98_clk sky130_fd_sc_hd__clkbuf_16
X_25914_ clknet_leaf_67_clk _00787_ net8648 VGND VGND VPWR VPWR pid_q.out\[10\] sky130_fd_sc_hd__dfrtp_1
X_21037_ net5528 net5950 net5930 net5910 VGND VGND VPWR VPWR _01053_ sky130_fd_sc_hd__a22o_1
Xwire1202 net1203 VGND VGND VPWR VPWR net1202 sky130_fd_sc_hd__buf_1
Xwire1213 _09823_ VGND VGND VPWR VPWR net1213 sky130_fd_sc_hd__buf_1
Xwire1224 net1227 VGND VGND VPWR VPWR net1224 sky130_fd_sc_hd__clkbuf_1
Xwire1235 net1236 VGND VGND VPWR VPWR net1235 sky130_fd_sc_hd__clkbuf_1
Xwire1246 _08463_ VGND VGND VPWR VPWR net1246 sky130_fd_sc_hd__buf_1
X_25845_ clknet_leaf_38_clk _00718_ net8747 VGND VGND VPWR VPWR pid_q.mult0.b\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1257 _08071_ VGND VGND VPWR VPWR net1257 sky130_fd_sc_hd__buf_1
Xwire1268 _07665_ VGND VGND VPWR VPWR net1268 sky130_fd_sc_hd__buf_1
Xwire1279 _07185_ VGND VGND VPWR VPWR net1279 sky130_fd_sc_hd__clkbuf_1
X_12810_ _05081_ _05082_ _04998_ _04972_ VGND VGND VPWR VPWR _05083_ sky130_fd_sc_hd__a2bb2o_1
X_13790_ net7653 net1962 _05975_ VGND VGND VPWR VPWR _06058_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25776_ clknet_leaf_57_clk _00649_ net8711 VGND VGND VPWR VPWR matmul0.beta_pass\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_22988_ net9235 _08738_ net6574 VGND VGND VPWR VPWR _02862_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24727_ net8012 _04560_ VGND VGND VPWR VPWR _04561_ sky130_fd_sc_hd__xor2_1
X_12741_ _04904_ net2989 VGND VGND VPWR VPWR _05014_ sky130_fd_sc_hd__and2_1
X_21939_ _01837_ _01839_ _01838_ VGND VGND VPWR VPWR _01947_ sky130_fd_sc_hd__o21a_1
XFILLER_0_167_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15460_ _07179_ VGND VGND VPWR VPWR _07534_ sky130_fd_sc_hd__clkbuf_1
X_24658_ net9177 net1378 _04511_ VGND VGND VPWR VPWR _00681_ sky130_fd_sc_hd__a21o_1
X_12672_ _04942_ _04943_ _04944_ VGND VGND VPWR VPWR _04945_ sky130_fd_sc_hd__a21o_2
XFILLER_0_195_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8747 net8751 VGND VGND VPWR VPWR net8747 sky130_fd_sc_hd__clkbuf_2
X_14411_ _06612_ VGND VGND VPWR VPWR _00087_ sky130_fd_sc_hd__clkbuf_1
X_23609_ pid_q.prev_error\[2\] pid_q.curr_error\[2\] VGND VGND VPWR VPWR _03477_ sky130_fd_sc_hd__xor2_1
Xwire8820 net8821 VGND VGND VPWR VPWR net8820 sky130_fd_sc_hd__clkbuf_1
Xfanout8769 net8796 VGND VGND VPWR VPWR net8769 sky130_fd_sc_hd__buf_1
Xwire8831 net8839 VGND VGND VPWR VPWR net8831 sky130_fd_sc_hd__clkbuf_1
X_15391_ _07462_ _07463_ _07414_ _07464_ VGND VGND VPWR VPWR _07465_ sky130_fd_sc_hd__o22a_1
XFILLER_0_38_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8842 net8843 VGND VGND VPWR VPWR net8842 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24589_ net263 _04444_ VGND VGND VPWR VPWR _04445_ sky130_fd_sc_hd__xor2_1
XFILLER_0_38_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8853 net8854 VGND VGND VPWR VPWR net8853 sky130_fd_sc_hd__clkbuf_1
X_17130_ net1221 _09084_ VGND VGND VPWR VPWR _09085_ sky130_fd_sc_hd__nand2_1
XFILLER_0_181_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8864 net8865 VGND VGND VPWR VPWR net8864 sky130_fd_sc_hd__buf_1
Xwire510 _04177_ VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__buf_1
X_14342_ _06558_ matmul0.a_in\[5\] net902 VGND VGND VPWR VPWR _06559_ sky130_fd_sc_hd__mux2_1
Xwire521 _02415_ VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8886 net127 VGND VGND VPWR VPWR net8886 sky130_fd_sc_hd__clkbuf_1
Xwire532 _06075_ VGND VGND VPWR VPWR net532 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_123_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8897 net8898 VGND VGND VPWR VPWR net8897 sky130_fd_sc_hd__clkbuf_2
Xwire543 net544 VGND VGND VPWR VPWR net543 sky130_fd_sc_hd__clkbuf_1
Xmax_length3850 _12269_ VGND VGND VPWR VPWR net3850 sky130_fd_sc_hd__buf_1
XFILLER_0_80_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17061_ _09019_ VGND VGND VPWR VPWR _09020_ sky130_fd_sc_hd__inv_2
Xwire554 net555 VGND VGND VPWR VPWR net554 sky130_fd_sc_hd__clkbuf_1
X_14273_ net2922 VGND VGND VPWR VPWR _06517_ sky130_fd_sc_hd__clkbuf_2
Xwire565 net566 VGND VGND VPWR VPWR net565 sky130_fd_sc_hd__clkbuf_1
Xwire576 _07556_ VGND VGND VPWR VPWR net576 sky130_fd_sc_hd__clkbuf_1
Xwire587 _04248_ VGND VGND VPWR VPWR net587 sky130_fd_sc_hd__buf_1
X_16012_ _07997_ _08078_ _08079_ VGND VGND VPWR VPWR _08080_ sky130_fd_sc_hd__a21oi_1
Xwire598 _02454_ VGND VGND VPWR VPWR net598 sky130_fd_sc_hd__clkbuf_1
X_13224_ net7674 net2350 net2346 VGND VGND VPWR VPWR _05497_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13155_ net917 _05426_ _05427_ VGND VGND VPWR VPWR _05428_ sky130_fd_sc_hd__and3_1
XFILLER_0_176_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13086_ _05269_ _05358_ _05275_ VGND VGND VPWR VPWR _05359_ sky130_fd_sc_hd__a21oi_1
X_17963_ _09690_ _09633_ VGND VGND VPWR VPWR _09814_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3160 _11293_ VGND VGND VPWR VPWR net3160 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_89_clk clknet_4_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_89_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_109_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3171 net3172 VGND VGND VPWR VPWR net3171 sky130_fd_sc_hd__clkbuf_1
X_19702_ _11380_ _11384_ _11537_ VGND VGND VPWR VPWR _11538_ sky130_fd_sc_hd__a21oi_1
Xwire3182 _11037_ VGND VGND VPWR VPWR net3182 sky130_fd_sc_hd__clkbuf_1
X_16914_ net6410 _08872_ _08873_ net9247 VGND VGND VPWR VPWR _08878_ sky130_fd_sc_hd__o211a_1
Xwire3193 net3194 VGND VGND VPWR VPWR net3193 sky130_fd_sc_hd__buf_1
X_17894_ _09742_ net2553 _09744_ VGND VGND VPWR VPWR _09745_ sky130_fd_sc_hd__o21a_1
Xwire2470 _02362_ VGND VGND VPWR VPWR net2470 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_189_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19633_ _11458_ _11469_ VGND VGND VPWR VPWR _11470_ sky130_fd_sc_hd__xnor2_2
Xwire2481 _00905_ VGND VGND VPWR VPWR net2481 sky130_fd_sc_hd__buf_1
Xwire2492 _12278_ VGND VGND VPWR VPWR net2492 sky130_fd_sc_hd__buf_1
X_16845_ _08813_ VGND VGND VPWR VPWR _00320_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1780 _09714_ VGND VGND VPWR VPWR net1780 sky130_fd_sc_hd__buf_1
Xwire1791 _09538_ VGND VGND VPWR VPWR net1791 sky130_fd_sc_hd__buf_1
X_19564_ _11190_ _11191_ VGND VGND VPWR VPWR _11401_ sky130_fd_sc_hd__and2_1
X_16776_ _08777_ VGND VGND VPWR VPWR _00287_ sky130_fd_sc_hd__clkbuf_1
X_13988_ _06192_ _06194_ _06252_ VGND VGND VPWR VPWR _06253_ sky130_fd_sc_hd__o21a_1
XFILLER_0_189_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15727_ _07792_ _07797_ VGND VGND VPWR VPWR _07798_ sky130_fd_sc_hd__xnor2_2
X_18515_ net7013 net6915 VGND VGND VPWR VPWR _10364_ sky130_fd_sc_hd__xnor2_2
X_12939_ net7917 net1350 VGND VGND VPWR VPWR _05212_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19495_ _11331_ VGND VGND VPWR VPWR _11332_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15658_ net988 _07729_ VGND VGND VPWR VPWR _07730_ sky130_fd_sc_hd__nand2_1
X_18446_ net7014 _10295_ _10041_ VGND VGND VPWR VPWR _10296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14609_ _06768_ _06777_ VGND VGND VPWR VPWR _06782_ sky130_fd_sc_hd__nor2_1
X_18377_ net6927 _10226_ _10227_ net3311 _10043_ VGND VGND VPWR VPWR _10228_ sky130_fd_sc_hd__a221o_1
XFILLER_0_69_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15589_ net1859 _07582_ _07576_ VGND VGND VPWR VPWR _07661_ sky130_fd_sc_hd__a21o_1
XFILLER_0_84_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_13_clk clknet_4_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_16
X_17328_ net4028 net7608 _09239_ _09241_ VGND VGND VPWR VPWR _09242_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_154_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17259_ net7606 net2960 net153 net2163 net9214 VGND VGND VPWR VPWR _00357_ sky130_fd_sc_hd__a32o_1
XFILLER_0_4_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20270_ net5 _12079_ VGND VGND VPWR VPWR _12080_ sky130_fd_sc_hd__xor2_1
XFILLER_0_70_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23960_ _03806_ _03823_ VGND VGND VPWR VPWR _03824_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_166_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22911_ net5340 pid_d.curr_int\[11\] VGND VGND VPWR VPWR _02803_ sky130_fd_sc_hd__xnor2_1
Xmax_length8806 net8803 VGND VGND VPWR VPWR net8806 sky130_fd_sc_hd__buf_1
X_23891_ _03754_ _03755_ VGND VGND VPWR VPWR _03756_ sky130_fd_sc_hd__nor2_1
XFILLER_0_190_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25630_ clknet_leaf_108_clk _00503_ net8351 VGND VGND VPWR VPWR cordic0.vec\[0\]\[2\]
+ sky130_fd_sc_hd__dfstp_1
X_22842_ pid_d.out\[3\] _02741_ net3065 VGND VGND VPWR VPWR _02742_ sky130_fd_sc_hd__mux2_1
X_25561_ clknet_leaf_115_clk _00434_ net8336 VGND VGND VPWR VPWR cordic0.gm0.iter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_22773_ _02693_ VGND VGND VPWR VPWR _00614_ sky130_fd_sc_hd__clkbuf_1
X_24512_ _04279_ _04307_ _04270_ VGND VGND VPWR VPWR _04369_ sky130_fd_sc_hd__o21a_1
X_21724_ net4385 _01648_ net524 net4318 net946 VGND VGND VPWR VPWR _01735_ sky130_fd_sc_hd__a221o_1
X_25492_ clknet_leaf_48_clk _00372_ net8759 VGND VGND VPWR VPWR svm0.tA\[14\] sky130_fd_sc_hd__dfrtp_1
Xwire8105 net85 VGND VGND VPWR VPWR net8105 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8116 net8117 VGND VGND VPWR VPWR net8116 sky130_fd_sc_hd__clkbuf_1
X_24443_ _04299_ _04300_ VGND VGND VPWR VPWR _04301_ sky130_fd_sc_hd__xor2_1
XFILLER_0_93_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21655_ net5744 net5516 VGND VGND VPWR VPWR _01666_ sky130_fd_sc_hd__nand2_1
Xwire8127 net8128 VGND VGND VPWR VPWR net8127 sky130_fd_sc_hd__clkbuf_1
Xwire8138 net8139 VGND VGND VPWR VPWR net8138 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7404 matmul0.matmul_stage_inst.a\[3\] VGND VGND VPWR VPWR net7404 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8149 net8150 VGND VGND VPWR VPWR net8149 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7415 net7416 VGND VGND VPWR VPWR net7415 sky130_fd_sc_hd__clkbuf_1
X_20606_ net1480 net1396 VGND VGND VPWR VPWR _12387_ sky130_fd_sc_hd__nand2_1
Xwire7426 matmul0.matmul_stage_inst.b\[6\] VGND VGND VPWR VPWR net7426 sky130_fd_sc_hd__clkbuf_1
X_24374_ _04231_ _04232_ net4589 VGND VGND VPWR VPWR _04233_ sky130_fd_sc_hd__mux2_1
Xwire7437 net7438 VGND VGND VPWR VPWR net7437 sky130_fd_sc_hd__buf_1
XFILLER_0_145_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21586_ _01489_ _01493_ _01487_ VGND VGND VPWR VPWR _01598_ sky130_fd_sc_hd__a21o_1
Xwire6703 net6704 VGND VGND VPWR VPWR net6703 sky130_fd_sc_hd__buf_1
XFILLER_0_61_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6714 net6715 VGND VGND VPWR VPWR net6714 sky130_fd_sc_hd__buf_1
Xwire6725 net6726 VGND VGND VPWR VPWR net6725 sky130_fd_sc_hd__clkbuf_1
X_23325_ _03193_ _03194_ VGND VGND VPWR VPWR _03195_ sky130_fd_sc_hd__xnor2_1
Xwire6736 svm0.counter\[2\] VGND VGND VPWR VPWR net6736 sky130_fd_sc_hd__buf_1
Xmax_length3168 _11132_ VGND VGND VPWR VPWR net3168 sky130_fd_sc_hd__clkbuf_1
X_20537_ net1398 _12321_ _12322_ net6306 net8056 VGND VGND VPWR VPWR _00504_ sky130_fd_sc_hd__o32a_1
Xwire6747 svm0.tB\[13\] VGND VGND VPWR VPWR net6747 sky130_fd_sc_hd__buf_1
XFILLER_0_105_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6758 net6755 VGND VGND VPWR VPWR net6758 sky130_fd_sc_hd__clkbuf_1
X_23256_ _03097_ _03125_ VGND VGND VPWR VPWR _03126_ sky130_fd_sc_hd__xnor2_2
Xmax_length2467 net2468 VGND VGND VPWR VPWR net2467 sky130_fd_sc_hd__buf_1
X_20468_ _12133_ _12258_ VGND VGND VPWR VPWR _12259_ sky130_fd_sc_hd__xnor2_1
X_22207_ net5690 net5466 VGND VGND VPWR VPWR _02212_ sky130_fd_sc_hd__nand2_1
X_23187_ net5139 net4698 VGND VGND VPWR VPWR _03057_ sky130_fd_sc_hd__nand2_1
X_20399_ cordic0.slte0.opA\[8\] net865 VGND VGND VPWR VPWR _12197_ sky130_fd_sc_hd__nand2_1
X_22138_ _02141_ _02143_ VGND VGND VPWR VPWR _02144_ sky130_fd_sc_hd__xnor2_1
X_14960_ _07018_ net4146 net4139 _07027_ VGND VGND VPWR VPWR _07034_ sky130_fd_sc_hd__o22a_1
XFILLER_0_100_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22069_ net1716 _01967_ VGND VGND VPWR VPWR _02076_ sky130_fd_sc_hd__and2_1
Xwire1010 _04549_ VGND VGND VPWR VPWR net1010 sky130_fd_sc_hd__buf_1
Xhold9 net150 VGND VGND VPWR VPWR net8962 sky130_fd_sc_hd__dlygate4sd3_1
Xwire1021 net1022 VGND VGND VPWR VPWR net1021 sky130_fd_sc_hd__clkbuf_1
Xwire1032 _02921_ VGND VGND VPWR VPWR net1032 sky130_fd_sc_hd__buf_1
X_13911_ net7632 net7611 VGND VGND VPWR VPWR _06177_ sky130_fd_sc_hd__and2_1
Xwire1043 _02051_ VGND VGND VPWR VPWR net1043 sky130_fd_sc_hd__clkbuf_1
X_14891_ net6631 matmul0.matmul_stage_inst.d\[11\] net7405 net6533 VGND VGND VPWR
+ VPWR _06965_ sky130_fd_sc_hd__a22o_1
Xwire1054 _12145_ VGND VGND VPWR VPWR net1054 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1065 _10578_ VGND VGND VPWR VPWR net1065 sky130_fd_sc_hd__clkbuf_2
Xwire1076 net1077 VGND VGND VPWR VPWR net1076 sky130_fd_sc_hd__buf_1
X_16630_ _08667_ _08668_ VGND VGND VPWR VPWR _08669_ sky130_fd_sc_hd__xnor2_1
X_13842_ _06056_ _06107_ _06108_ VGND VGND VPWR VPWR _06109_ sky130_fd_sc_hd__a21o_1
X_25828_ clknet_leaf_36_clk _00701_ net8753 VGND VGND VPWR VPWR pid_q.curr_error\[4\]
+ sky130_fd_sc_hd__dfrtp_2
Xwire1087 _08290_ VGND VGND VPWR VPWR net1087 sky130_fd_sc_hd__clkbuf_2
Xwire1098 _07758_ VGND VGND VPWR VPWR net1098 sky130_fd_sc_hd__clkbuf_1
X_16561_ _08529_ _08572_ _08619_ VGND VGND VPWR VPWR _08620_ sky130_fd_sc_hd__o21a_1
X_13773_ _06039_ _06033_ _06034_ VGND VGND VPWR VPWR _06041_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25759_ clknet_leaf_95_clk _00632_ net8402 VGND VGND VPWR VPWR pid_d.out\[0\] sky130_fd_sc_hd__dfrtp_2
X_15512_ net1861 net1860 VGND VGND VPWR VPWR _07585_ sky130_fd_sc_hd__nand2_1
X_18300_ net815 _10147_ _10137_ _10149_ VGND VGND VPWR VPWR _10151_ sky130_fd_sc_hd__nand4_1
X_12724_ _04985_ _04995_ _04996_ VGND VGND VPWR VPWR _04997_ sky130_fd_sc_hd__a21o_2
X_19280_ _11111_ _11113_ _11115_ _11116_ VGND VGND VPWR VPWR _11117_ sky130_fd_sc_hd__a22o_1
X_16492_ _08522_ net975 VGND VGND VPWR VPWR _08552_ sky130_fd_sc_hd__or2_1
XFILLER_0_183_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18231_ _10053_ _10080_ _10081_ VGND VGND VPWR VPWR _10082_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15443_ net3602 net3419 VGND VGND VPWR VPWR _07517_ sky130_fd_sc_hd__nor2_1
XFILLER_0_182_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12655_ net6751 net6600 net5308 VGND VGND VPWR VPWR _04928_ sky130_fd_sc_hd__and3_1
Xfanout8555 net8590 VGND VGND VPWR VPWR net8555 sky130_fd_sc_hd__buf_1
Xwire8650 net8649 VGND VGND VPWR VPWR net8650 sky130_fd_sc_hd__clkbuf_2
X_18162_ _10001_ _10006_ _10008_ _10009_ _10012_ VGND VGND VPWR VPWR _10013_ sky130_fd_sc_hd__a311oi_1
XFILLER_0_108_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15374_ _07441_ _07446_ _07447_ VGND VGND VPWR VPWR _07448_ sky130_fd_sc_hd__a21o_1
X_12586_ net3019 VGND VGND VPWR VPWR _00011_ sky130_fd_sc_hd__buf_1
XFILLER_0_68_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8672 net8669 VGND VGND VPWR VPWR net8672 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire8683 net8680 VGND VGND VPWR VPWR net8683 sky130_fd_sc_hd__dlymetal6s2s_1
X_17113_ net3332 VGND VGND VPWR VPWR _09069_ sky130_fd_sc_hd__buf_1
XFILLER_0_154_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8694 net8695 VGND VGND VPWR VPWR net8694 sky130_fd_sc_hd__clkbuf_2
Xwire340 net341 VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__clkbuf_1
X_14325_ net7356 net1299 net2896 pid_d.out\[1\] _06545_ VGND VGND VPWR VPWR _06546_
+ sky130_fd_sc_hd__a221o_1
Xwire7960 pid_q.target\[14\] VGND VGND VPWR VPWR net7960 sky130_fd_sc_hd__clkbuf_1
X_18093_ _09932_ _09938_ VGND VGND VPWR VPWR _09944_ sky130_fd_sc_hd__or2_1
Xwire351 _11735_ VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__buf_1
XFILLER_0_167_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7971 net7972 VGND VGND VPWR VPWR net7971 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7982 net7983 VGND VGND VPWR VPWR net7982 sky130_fd_sc_hd__clkbuf_1
Xwire362 net363 VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__clkbuf_1
Xwire373 _04617_ VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7993 net7994 VGND VGND VPWR VPWR net7993 sky130_fd_sc_hd__clkbuf_1
X_17044_ net3328 net1231 _09001_ _09003_ VGND VGND VPWR VPWR _00329_ sky130_fd_sc_hd__a31o_1
Xwire384 _08730_ VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14256_ net6451 _06497_ VGND VGND VPWR VPWR _06510_ sky130_fd_sc_hd__nor2_1
Xwire395 _08010_ VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__clkbuf_1
X_13207_ _05475_ _05479_ VGND VGND VPWR VPWR _05480_ sky130_fd_sc_hd__xnor2_1
Xmax_length2990 net2991 VGND VGND VPWR VPWR net2990 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_110_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14187_ _05972_ _06446_ VGND VGND VPWR VPWR _06447_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13138_ _05388_ _05389_ _05393_ _05410_ net1585 VGND VGND VPWR VPWR _05411_ sky130_fd_sc_hd__a32o_1
XFILLER_0_29_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18995_ _10827_ net3212 _10829_ _10831_ net6266 VGND VGND VPWR VPWR _10832_ sky130_fd_sc_hd__a311o_1
XFILLER_0_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13069_ _05338_ _05341_ VGND VGND VPWR VPWR _05342_ sky130_fd_sc_hd__xnor2_2
X_17946_ net3956 _09676_ _09796_ VGND VGND VPWR VPWR _09797_ sky130_fd_sc_hd__o21bai_1
Xclkbuf_leaf_2_clk clknet_4_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_174_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_119_Right_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17877_ net1780 _09722_ _09727_ VGND VGND VPWR VPWR _09728_ sky130_fd_sc_hd__o21ba_1
X_19616_ net6087 net6102 VGND VGND VPWR VPWR _11453_ sky130_fd_sc_hd__nor2_1
X_16828_ cordic0.sin\[2\] matmul0.sin\[2\] net3365 VGND VGND VPWR VPWR _08805_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19547_ net6105 _11328_ _11381_ net3151 _11383_ VGND VGND VPWR VPWR _11384_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16759_ _08768_ VGND VGND VPWR VPWR _00279_ sky130_fd_sc_hd__clkbuf_1
X_19478_ _11310_ _11313_ _11314_ net6359 VGND VGND VPWR VPWR _11315_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_75_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18429_ net6785 net3283 VGND VGND VPWR VPWR _10279_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21440_ _01349_ _01354_ _01348_ VGND VGND VPWR VPWR _01453_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_185_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21371_ _01379_ _01384_ VGND VGND VPWR VPWR _01385_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5309 net5310 VGND VGND VPWR VPWR net5309 sky130_fd_sc_hd__clkbuf_1
X_23110_ _02900_ _02901_ VGND VGND VPWR VPWR _02980_ sky130_fd_sc_hd__xnor2_1
X_20322_ net951 _12125_ VGND VGND VPWR VPWR _12126_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24090_ net7523 _03865_ net329 net7462 net741 VGND VGND VPWR VPWR _03953_ sky130_fd_sc_hd__a221o_1
Xwire4608 net4602 VGND VGND VPWR VPWR net4608 sky130_fd_sc_hd__buf_1
XFILLER_0_141_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4619 net4620 VGND VGND VPWR VPWR net4619 sky130_fd_sc_hd__buf_1
X_23041_ net5142 net4610 VGND VGND VPWR VPWR _02911_ sky130_fd_sc_hd__nand2_1
X_20253_ net16 _12066_ VGND VGND VPWR VPWR _12067_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3918 net3919 VGND VGND VPWR VPWR net3918 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_177_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3929 net3930 VGND VGND VPWR VPWR net3929 sky130_fd_sc_hd__buf_1
XFILLER_0_122_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20184_ net2580 _11648_ _12005_ _12009_ VGND VGND VPWR VPWR _12010_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_177_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24992_ net4475 _04732_ _04734_ VGND VGND VPWR VPWR _04751_ sky130_fd_sc_hd__mux2_1
X_23943_ net4559 net4951 VGND VGND VPWR VPWR _03807_ sky130_fd_sc_hd__nand2_2
XFILLER_0_192_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23874_ net3747 VGND VGND VPWR VPWR _03739_ sky130_fd_sc_hd__clkbuf_1
Xmax_length7924 net7925 VGND VGND VPWR VPWR net7924 sky130_fd_sc_hd__clkbuf_1
X_25613_ clknet_leaf_109_clk _00486_ net8352 VGND VGND VPWR VPWR cordic0.slte0.opA\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xmax_length7935 net7936 VGND VGND VPWR VPWR net7935 sky130_fd_sc_hd__clkbuf_1
X_22825_ net5366 net3065 _02726_ net8897 VGND VGND VPWR VPWR _00633_ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25544_ clknet_leaf_30_clk net9203 net8676 VGND VGND VPWR VPWR pid_q.prev_int\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_22756_ net4303 net8092 VGND VGND VPWR VPWR _02682_ sky130_fd_sc_hd__and2_1
XFILLER_0_165_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21707_ _01654_ _01717_ VGND VGND VPWR VPWR _01718_ sky130_fd_sc_hd__xnor2_2
Xfanout7106 net7117 VGND VGND VPWR VPWR net7106 sky130_fd_sc_hd__buf_1
X_25475_ clknet_leaf_47_clk _00355_ net8775 VGND VGND VPWR VPWR svm0.tB\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22687_ pid_d.ki\[6\] net2440 net2993 pid_d.kp\[6\] VGND VGND VPWR VPWR _02633_ sky130_fd_sc_hd__a22o_1
Xfanout7139 net7145 VGND VGND VPWR VPWR net7139 sky130_fd_sc_hd__buf_1
X_24426_ net1651 net1650 VGND VGND VPWR VPWR _04284_ sky130_fd_sc_hd__xor2_4
XFILLER_0_118_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7212 net7213 VGND VGND VPWR VPWR net7212 sky130_fd_sc_hd__buf_1
X_21638_ net600 _01631_ _01632_ VGND VGND VPWR VPWR _01649_ sky130_fd_sc_hd__a21o_1
XFILLER_0_180_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7223 net7224 VGND VGND VPWR VPWR net7223 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7234 net7235 VGND VGND VPWR VPWR net7234 sky130_fd_sc_hd__buf_1
Xwire6500 net6498 VGND VGND VPWR VPWR net6500 sky130_fd_sc_hd__buf_1
XFILLER_0_62_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire7256 net7258 VGND VGND VPWR VPWR net7256 sky130_fd_sc_hd__clkbuf_1
Xwire6511 net6506 VGND VGND VPWR VPWR net6511 sky130_fd_sc_hd__buf_1
XFILLER_0_35_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24357_ net4960 net4937 net3041 VGND VGND VPWR VPWR _04216_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21569_ _01575_ _01580_ VGND VGND VPWR VPWR _01581_ sky130_fd_sc_hd__xnor2_1
Xwire7267 net7268 VGND VGND VPWR VPWR net7267 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7278 net7279 VGND VGND VPWR VPWR net7278 sky130_fd_sc_hd__clkbuf_2
Xwire6533 net6531 VGND VGND VPWR VPWR net6533 sky130_fd_sc_hd__clkbuf_2
X_14110_ _06341_ _06343_ _06342_ VGND VGND VPWR VPWR _06372_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_62_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7289 net7290 VGND VGND VPWR VPWR net7289 sky130_fd_sc_hd__clkbuf_1
X_23308_ _02965_ _03176_ _03177_ net1677 VGND VGND VPWR VPWR _03178_ sky130_fd_sc_hd__a2bb2o_1
Xwire6555 net6556 VGND VGND VPWR VPWR net6555 sky130_fd_sc_hd__clkbuf_1
Xwire5810 net5811 VGND VGND VPWR VPWR net5810 sky130_fd_sc_hd__buf_1
XFILLER_0_132_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15090_ net1280 net1117 VGND VGND VPWR VPWR _07164_ sky130_fd_sc_hd__xnor2_1
Xwire6566 matmul0.matmul_stage_inst.state\[6\] VGND VGND VPWR VPWR net6566 sky130_fd_sc_hd__buf_1
Xwire5821 net5822 VGND VGND VPWR VPWR net5821 sky130_fd_sc_hd__clkbuf_2
X_24288_ net4937 _04146_ _04147_ VGND VGND VPWR VPWR _04148_ sky130_fd_sc_hd__a21o_1
Xwire5832 net5836 VGND VGND VPWR VPWR net5832 sky130_fd_sc_hd__buf_1
Xwire6577 net6578 VGND VGND VPWR VPWR net6577 sky130_fd_sc_hd__clkbuf_1
Xwire6588 net6590 VGND VGND VPWR VPWR net6588 sky130_fd_sc_hd__buf_1
Xwire5843 net5844 VGND VGND VPWR VPWR net5843 sky130_fd_sc_hd__buf_1
X_14041_ _06295_ _06304_ VGND VGND VPWR VPWR _06305_ sky130_fd_sc_hd__xnor2_2
Xwire6599 net6600 VGND VGND VPWR VPWR net6599 sky130_fd_sc_hd__buf_1
Xwire5854 net5855 VGND VGND VPWR VPWR net5854 sky130_fd_sc_hd__clkbuf_1
X_23239_ _03093_ _03095_ _03094_ VGND VGND VPWR VPWR _03109_ sky130_fd_sc_hd__o21a_1
Xwire5865 net5866 VGND VGND VPWR VPWR net5865 sky130_fd_sc_hd__buf_1
Xwire5876 net5877 VGND VGND VPWR VPWR net5876 sky130_fd_sc_hd__clkbuf_1
Xwire5898 net5895 VGND VGND VPWR VPWR net5898 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_152_Left_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17800_ net3263 _09650_ net7132 VGND VGND VPWR VPWR _09651_ sky130_fd_sc_hd__a21oi_1
X_15992_ _08049_ _08059_ VGND VGND VPWR VPWR _08060_ sky130_fd_sc_hd__xor2_1
X_18780_ _10565_ _10601_ VGND VGND VPWR VPWR _10624_ sky130_fd_sc_hd__nand2_1
X_17731_ net6475 _09588_ VGND VGND VPWR VPWR _00432_ sky130_fd_sc_hd__xnor2_1
X_14943_ _07012_ _07016_ VGND VGND VPWR VPWR _07017_ sky130_fd_sc_hd__nand2_1
X_17662_ net4007 svm0.tA\[7\] svm0.tA\[5\] net4021 _09541_ VGND VGND VPWR VPWR _09542_
+ sky130_fd_sc_hd__o221a_1
X_14874_ matmul0.b\[9\] matmul0.matmul_stage_inst.f\[9\] net3604 VGND VGND VPWR VPWR
+ _06955_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19401_ _11155_ _11203_ _11233_ _11237_ VGND VGND VPWR VPWR _11238_ sky130_fd_sc_hd__a31o_1
X_13825_ net7708 net1307 VGND VGND VPWR VPWR _06092_ sky130_fd_sc_hd__nand2_1
X_16613_ _08656_ VGND VGND VPWR VPWR _00245_ sky130_fd_sc_hd__clkbuf_1
X_17593_ _09472_ _09473_ VGND VGND VPWR VPWR _09474_ sky130_fd_sc_hd__nor2_1
X_19332_ net6352 net2525 VGND VGND VPWR VPWR _11169_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16544_ _08559_ _08601_ _08602_ net2791 VGND VGND VPWR VPWR _08603_ sky130_fd_sc_hd__a22o_1
X_13756_ _05961_ _06022_ _06023_ VGND VGND VPWR VPWR _06024_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_161_Left_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12707_ net7854 net1974 net1971 VGND VGND VPWR VPWR _04980_ sky130_fd_sc_hd__and3_2
X_19263_ _10904_ net1758 VGND VGND VPWR VPWR _11100_ sky130_fd_sc_hd__nand2_1
X_16475_ _08467_ _08472_ _08535_ VGND VGND VPWR VPWR _08536_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_167_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13687_ _05881_ _05886_ VGND VGND VPWR VPWR _05956_ sky130_fd_sc_hd__and2b_1
XFILLER_0_31_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15426_ net1543 net2703 _07499_ VGND VGND VPWR VPWR _07500_ sky130_fd_sc_hd__a21oi_1
X_18214_ net6894 net6856 VGND VGND VPWR VPWR _10065_ sky130_fd_sc_hd__nand2_1
X_12638_ net6750 net6600 net5284 VGND VGND VPWR VPWR _04911_ sky130_fd_sc_hd__and3_1
X_19194_ _10898_ _10813_ VGND VGND VPWR VPWR _11031_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8385 net8393 VGND VGND VPWR VPWR net8385 sky130_fd_sc_hd__buf_1
XFILLER_0_54_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8480 net8481 VGND VGND VPWR VPWR net8480 sky130_fd_sc_hd__clkbuf_1
Xfanout7684 net7699 VGND VGND VPWR VPWR net7684 sky130_fd_sc_hd__buf_1
X_18145_ _09985_ _09986_ _09992_ _09995_ VGND VGND VPWR VPWR _09996_ sky130_fd_sc_hd__or4_1
X_15357_ net1116 _07430_ VGND VGND VPWR VPWR _07431_ sky130_fd_sc_hd__nand2_1
X_12569_ net2388 VGND VGND VPWR VPWR _04859_ sky130_fd_sc_hd__buf_1
Xwire8491 net8488 VGND VGND VPWR VPWR net8491 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout6961 cordic0.vec\[1\]\[8\] VGND VGND VPWR VPWR net6961 sky130_fd_sc_hd__buf_1
XFILLER_0_41_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14308_ net6453 VGND VGND VPWR VPWR _06530_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire170 net171 VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_1
Xwire7790 net7786 VGND VGND VPWR VPWR net7790 sky130_fd_sc_hd__buf_1
XFILLER_0_25_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18076_ net3987 net3942 VGND VGND VPWR VPWR _09927_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold206 pid_d.prev_error\[13\] VGND VGND VPWR VPWR net9159 sky130_fd_sc_hd__dlygate4sd3_1
X_15288_ net2757 net3483 VGND VGND VPWR VPWR _07362_ sky130_fd_sc_hd__nor2_1
Xwire181 net182 VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__buf_1
Xwire192 _06152_ VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__buf_1
XFILLER_0_124_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold217 _00803_ VGND VGND VPWR VPWR net9170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 pid_d.prev_error\[11\] VGND VGND VPWR VPWR net9181 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17027_ net4048 net4237 VGND VGND VPWR VPWR _08987_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14239_ net7606 net2373 net153 _05779_ net9194 VGND VGND VPWR VPWR _00032_ sky130_fd_sc_hd__a32o_1
Xhold239 matmul0.op_in\[0\] VGND VGND VPWR VPWR net9192 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_170_Left_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18978_ net3902 _10814_ net6260 VGND VGND VPWR VPWR _10815_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17929_ net2145 net2143 VGND VGND VPWR VPWR _09780_ sky130_fd_sc_hd__nor2_1
X_20940_ _00952_ _00955_ VGND VGND VPWR VPWR _00956_ sky130_fd_sc_hd__nand2_1
X_20871_ _00880_ net2482 VGND VGND VPWR VPWR _00887_ sky130_fd_sc_hd__and2_1
XFILLER_0_178_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22610_ _02583_ VGND VGND VPWR VPWR _00561_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23590_ net4768 net4813 VGND VGND VPWR VPWR _03458_ sky130_fd_sc_hd__nand2_1
XFILLER_0_163_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22541_ pid_d.curr_error\[8\] net2381 net2048 VGND VGND VPWR VPWR _02533_ sky130_fd_sc_hd__and3_1
X_25260_ clknet_leaf_76_clk _00143_ net8458 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.b\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_22472_ net5713 net5732 net5753 VGND VGND VPWR VPWR _02473_ sky130_fd_sc_hd__or3_1
XFILLER_0_9_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24211_ _04069_ _04070_ VGND VGND VPWR VPWR _04072_ sky130_fd_sc_hd__or2_1
X_21423_ _01337_ _01338_ pid_d.prev_int\[2\] VGND VGND VPWR VPWR _01436_ sky130_fd_sc_hd__a21o_1
X_25191_ clknet_leaf_61_clk _00080_ net8721 VGND VGND VPWR VPWR matmul0.a_in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5106 net5107 VGND VGND VPWR VPWR net5106 sky130_fd_sc_hd__clkbuf_1
X_24142_ _03892_ _03918_ _03890_ VGND VGND VPWR VPWR _04004_ sky130_fd_sc_hd__o21a_1
XFILLER_0_115_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21354_ _01278_ _01279_ _01367_ VGND VGND VPWR VPWR _01368_ sky130_fd_sc_hd__a21oi_2
Xwire5128 net5129 VGND VGND VPWR VPWR net5128 sky130_fd_sc_hd__clkbuf_1
Xwire4405 pid_q.out\[13\] VGND VGND VPWR VPWR net4405 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4416 net4417 VGND VGND VPWR VPWR net4416 sky130_fd_sc_hd__clkbuf_1
X_20305_ net6467 _12109_ net1808 VGND VGND VPWR VPWR _12110_ sky130_fd_sc_hd__mux2_1
X_24073_ net1161 _03833_ _03742_ VGND VGND VPWR VPWR _03936_ sky130_fd_sc_hd__a21bo_1
Xwire4427 net4428 VGND VGND VPWR VPWR net4427 sky130_fd_sc_hd__clkbuf_1
X_21285_ _01288_ _01299_ VGND VGND VPWR VPWR _01300_ sky130_fd_sc_hd__xnor2_1
Xwire4438 net4439 VGND VGND VPWR VPWR net4438 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4449 net4450 VGND VGND VPWR VPWR net4449 sky130_fd_sc_hd__clkbuf_1
Xwire3704 _04877_ VGND VGND VPWR VPWR net3704 sky130_fd_sc_hd__buf_1
X_23024_ _02890_ _02893_ VGND VGND VPWR VPWR _02894_ sky130_fd_sc_hd__xnor2_2
Xwire3715 _04869_ VGND VGND VPWR VPWR net3715 sky130_fd_sc_hd__buf_1
XFILLER_0_40_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3726 _04867_ VGND VGND VPWR VPWR net3726 sky130_fd_sc_hd__clkbuf_1
X_20236_ _12053_ VGND VGND VPWR VPWR _00472_ sky130_fd_sc_hd__clkbuf_1
Xwire3737 _04038_ VGND VGND VPWR VPWR net3737 sky130_fd_sc_hd__buf_1
Xwire3759 net3760 VGND VGND VPWR VPWR net3759 sky130_fd_sc_hd__buf_1
X_20167_ _11927_ _11955_ _11991_ VGND VGND VPWR VPWR _11993_ sky130_fd_sc_hd__a21o_1
X_24975_ _04742_ VGND VGND VPWR VPWR _00767_ sky130_fd_sc_hd__clkbuf_1
X_20098_ net487 _11835_ _11873_ VGND VGND VPWR VPWR _11926_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_196_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23926_ net4635 net4855 VGND VGND VPWR VPWR _03790_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length8433 net8434 VGND VGND VPWR VPWR net8433 sky130_fd_sc_hd__clkbuf_1
Xmax_length8455 net8456 VGND VGND VPWR VPWR net8455 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_98_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length8466 net8467 VGND VGND VPWR VPWR net8466 sky130_fd_sc_hd__clkbuf_2
X_23857_ _03713_ _03721_ VGND VGND VPWR VPWR _03722_ sky130_fd_sc_hd__xnor2_2
Xmax_length7732 net7733 VGND VGND VPWR VPWR net7732 sky130_fd_sc_hd__clkbuf_1
Xmax_length8477 net8478 VGND VGND VPWR VPWR net8477 sky130_fd_sc_hd__clkbuf_2
X_13610_ _05786_ _05787_ VGND VGND VPWR VPWR _05880_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22808_ net4381 net4317 net4350 net4373 VGND VGND VPWR VPWR _02712_ sky130_fd_sc_hd__or4_1
Xmax_length7776 net7771 VGND VGND VPWR VPWR net7776 sky130_fd_sc_hd__clkbuf_1
X_14590_ net2882 _06763_ net281 VGND VGND VPWR VPWR _06765_ sky130_fd_sc_hd__o21ai_1
X_23788_ net1165 _03553_ _03552_ VGND VGND VPWR VPWR _03654_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_196_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25527_ clknet_leaf_45_clk net9001 net8788 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__dfrtp_1
X_13541_ _05810_ _05811_ VGND VGND VPWR VPWR _05812_ sky130_fd_sc_hd__xor2_1
X_22739_ pid_d.ki\[4\] _02670_ net1689 VGND VGND VPWR VPWR _02671_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16260_ _08270_ _08272_ _08271_ VGND VGND VPWR VPWR _08324_ sky130_fd_sc_hd__o21ba_1
X_13472_ net7655 net1975 net2311 VGND VGND VPWR VPWR _05745_ sky130_fd_sc_hd__and3_1
X_25458_ clknet_leaf_100_clk _00341_ net8389 VGND VGND VPWR VPWR cordic0.vec\[1\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7020 net7022 VGND VGND VPWR VPWR net7020 sky130_fd_sc_hd__buf_1
XFILLER_0_82_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15211_ net2828 net3453 _07195_ _07284_ VGND VGND VPWR VPWR _07285_ sky130_fd_sc_hd__a22o_1
X_24409_ _04264_ _04266_ VGND VGND VPWR VPWR _04267_ sky130_fd_sc_hd__nand2_1
Xwire7031 net7033 VGND VGND VPWR VPWR net7031 sky130_fd_sc_hd__buf_1
Xwire7042 net7039 VGND VGND VPWR VPWR net7042 sky130_fd_sc_hd__buf_1
XFILLER_0_30_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16191_ _08249_ _08255_ VGND VGND VPWR VPWR _08256_ sky130_fd_sc_hd__xnor2_2
Xfanout5512 pid_d.mult0.a\[8\] VGND VGND VPWR VPWR net5512 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25389_ clknet_leaf_74_clk _00272_ net8466 VGND VGND VPWR VPWR matmul0.b\[8\] sky130_fd_sc_hd__dfrtp_1
Xfanout5523 net5533 VGND VGND VPWR VPWR net5523 sky130_fd_sc_hd__clkbuf_1
Xwire7064 net7065 VGND VGND VPWR VPWR net7064 sky130_fd_sc_hd__buf_1
XFILLER_0_140_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout6268 net6282 VGND VGND VPWR VPWR net6268 sky130_fd_sc_hd__clkbuf_2
Xwire6330 net6331 VGND VGND VPWR VPWR net6330 sky130_fd_sc_hd__buf_1
Xwire7075 net7077 VGND VGND VPWR VPWR net7075 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15142_ _07202_ _07203_ _07214_ VGND VGND VPWR VPWR _07216_ sky130_fd_sc_hd__or3_1
Xfanout5556 net5569 VGND VGND VPWR VPWR net5556 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire6352 net6351 VGND VGND VPWR VPWR net6352 sky130_fd_sc_hd__buf_2
Xwire7097 net7096 VGND VGND VPWR VPWR net7097 sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_length2050 _02521_ VGND VGND VPWR VPWR net2050 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6363 net6364 VGND VGND VPWR VPWR net6363 sky130_fd_sc_hd__buf_1
XFILLER_0_51_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6374 cordic0.slte0.opA\[6\] VGND VGND VPWR VPWR net6374 sky130_fd_sc_hd__clkbuf_2
Xwire5640 net5644 VGND VGND VPWR VPWR net5640 sky130_fd_sc_hd__clkbuf_1
Xwire6385 cordic0.domain\[1\] VGND VGND VPWR VPWR net6385 sky130_fd_sc_hd__clkbuf_1
Xmax_length2072 _01434_ VGND VGND VPWR VPWR net2072 sky130_fd_sc_hd__clkbuf_1
Xwire6396 net6397 VGND VGND VPWR VPWR net6396 sky130_fd_sc_hd__buf_1
X_15073_ net2780 net2776 _07146_ VGND VGND VPWR VPWR _07147_ sky130_fd_sc_hd__and3_1
X_19950_ _11780_ _11781_ VGND VGND VPWR VPWR _11782_ sky130_fd_sc_hd__nand2_2
XFILLER_0_61_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5651 net5652 VGND VGND VPWR VPWR net5651 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire5662 net5663 VGND VGND VPWR VPWR net5662 sky130_fd_sc_hd__clkbuf_1
X_14024_ net7718 net1567 VGND VGND VPWR VPWR _06288_ sky130_fd_sc_hd__nand2_1
Xwire5684 pid_d.mult0.b\[14\] VGND VGND VPWR VPWR net5684 sky130_fd_sc_hd__clkbuf_1
X_18901_ _10735_ _10740_ VGND VGND VPWR VPWR _10742_ sky130_fd_sc_hd__or2_1
Xwire4950 net4951 VGND VGND VPWR VPWR net4950 sky130_fd_sc_hd__clkbuf_1
Xwire5695 net5696 VGND VGND VPWR VPWR net5695 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4961 net4956 VGND VGND VPWR VPWR net4961 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19881_ _11655_ _11659_ _11713_ VGND VGND VPWR VPWR _11714_ sky130_fd_sc_hd__o21ai_2
Xwire4972 net4973 VGND VGND VPWR VPWR net4972 sky130_fd_sc_hd__buf_1
Xwire4983 net4984 VGND VGND VPWR VPWR net4983 sky130_fd_sc_hd__buf_1
Xwire4994 net4995 VGND VGND VPWR VPWR net4994 sky130_fd_sc_hd__buf_1
X_18832_ net6896 net6829 net2588 VGND VGND VPWR VPWR _10675_ sky130_fd_sc_hd__and3_1
XFILLER_0_184_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18763_ net714 VGND VGND VPWR VPWR _10608_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15975_ _08038_ _08042_ VGND VGND VPWR VPWR _08043_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17714_ net9212 net1219 net1453 pid_q.curr_int\[5\] VGND VGND VPWR VPWR _00419_ sky130_fd_sc_hd__a22o_1
X_14926_ net6609 net7424 matmul0.matmul_stage_inst.a\[7\] net6585 VGND VGND VPWR VPWR
+ _07000_ sky130_fd_sc_hd__a22o_1
X_18694_ net6820 _10276_ _10285_ _10538_ _10539_ VGND VGND VPWR VPWR _10540_ sky130_fd_sc_hd__a221o_1
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17645_ net6701 svm0.tA\[12\] VGND VGND VPWR VPWR _09525_ sky130_fd_sc_hd__xor2_1
X_14857_ net7190 matmul0.matmul_stage_inst.f\[1\] net3608 VGND VGND VPWR VPWR _06946_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13808_ net621 _05990_ _05984_ VGND VGND VPWR VPWR _06076_ sky130_fd_sc_hd__o21a_1
XFILLER_0_129_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17576_ svm0.tC\[7\] _09430_ net4006 VGND VGND VPWR VPWR _09458_ sky130_fd_sc_hd__a21o_1
X_14788_ net9146 net3003 net992 VGND VGND VPWR VPWR _00166_ sky130_fd_sc_hd__o21a_1
XFILLER_0_133_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19315_ net2108 _11151_ VGND VGND VPWR VPWR _11152_ sky130_fd_sc_hd__xor2_1
X_13739_ net322 _06007_ VGND VGND VPWR VPWR _06008_ sky130_fd_sc_hd__nand2_1
X_16527_ _08554_ _08586_ VGND VGND VPWR VPWR _08587_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19246_ net6201 net6240 VGND VGND VPWR VPWR _11083_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16458_ net1244 _08518_ VGND VGND VPWR VPWR _08519_ sky130_fd_sc_hd__xor2_2
XFILLER_0_27_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout7470 pid_q.state\[4\] VGND VGND VPWR VPWR net7470 sky130_fd_sc_hd__buf_1
XFILLER_0_60_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15409_ net6621 net6640 matmul0.matmul_stage_inst.f\[13\] VGND VGND VPWR VPWR _07483_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_115_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19177_ net3187 VGND VGND VPWR VPWR _11014_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16389_ net2635 net2622 VGND VGND VPWR VPWR _08451_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18128_ net3347 net3265 _09978_ net3256 VGND VGND VPWR VPWR _09979_ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6780 net6783 VGND VGND VPWR VPWR net6780 sky130_fd_sc_hd__clkbuf_1
X_18059_ net7067 net7111 VGND VGND VPWR VPWR _09910_ sky130_fd_sc_hd__nand2_1
X_21070_ _01039_ _01085_ VGND VGND VPWR VPWR _01086_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_111_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20021_ net6081 _11797_ net3199 VGND VGND VPWR VPWR _11851_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_171_Right_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1609 _05015_ VGND VGND VPWR VPWR net1609 sky130_fd_sc_hd__clkbuf_1
X_24760_ net7990 net1638 VGND VGND VPWR VPWR _04590_ sky130_fd_sc_hd__xnor2_1
X_21972_ _01973_ _01979_ VGND VGND VPWR VPWR _01980_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_174_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23711_ pid_q.prev_int\[3\] VGND VGND VPWR VPWR _03577_ sky130_fd_sc_hd__inv_2
X_20923_ net5491 net5954 VGND VGND VPWR VPWR _00939_ sky130_fd_sc_hd__nand2_2
X_24691_ _04528_ VGND VGND VPWR VPWR _04529_ sky130_fd_sc_hd__buf_1
Xmax_length6305 net6301 VGND VGND VPWR VPWR net6305 sky130_fd_sc_hd__buf_1
XFILLER_0_95_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23642_ _03503_ _03508_ VGND VGND VPWR VPWR _03509_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_7_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20854_ net5473 _00868_ VGND VGND VPWR VPWR _00870_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23573_ net2420 _03361_ _03440_ VGND VGND VPWR VPWR _03441_ sky130_fd_sc_hd__a21o_1
X_20785_ net5636 net5625 VGND VGND VPWR VPWR _12556_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25312_ clknet_leaf_80_clk _00195_ net8511 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.e\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22524_ _02523_ VGND VGND VPWR VPWR _02524_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire906 _06199_ VGND VGND VPWR VPWR net906 sky130_fd_sc_hd__buf_1
Xwire917 _05411_ VGND VGND VPWR VPWR net917 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire928 _04311_ VGND VGND VPWR VPWR net928 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25243_ clknet_leaf_87_clk _00126_ net8442 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.a\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_22455_ net520 net597 VGND VGND VPWR VPWR _02457_ sky130_fd_sc_hd__and2_1
Xwire939 net940 VGND VGND VPWR VPWR net939 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21406_ net806 _01419_ VGND VGND VPWR VPWR _01420_ sky130_fd_sc_hd__xnor2_1
X_25174_ clknet_leaf_54_clk _00063_ net8730 VGND VGND VPWR VPWR svm0.periodTop\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_161_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22386_ _02387_ _02388_ VGND VGND VPWR VPWR _02389_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24125_ net4534 net4928 VGND VGND VPWR VPWR _03987_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21337_ _01348_ _01350_ VGND VGND VPWR VPWR _01351_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4213 _06969_ VGND VGND VPWR VPWR net4213 sky130_fd_sc_hd__buf_1
XFILLER_0_163_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4246 net4247 VGND VGND VPWR VPWR net4246 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3501 _07106_ VGND VGND VPWR VPWR net3501 sky130_fd_sc_hd__buf_1
X_24056_ _03892_ _03918_ VGND VGND VPWR VPWR _03919_ sky130_fd_sc_hd__xor2_1
Xwire3512 _07095_ VGND VGND VPWR VPWR net3512 sky130_fd_sc_hd__buf_1
Xwire4257 net4258 VGND VGND VPWR VPWR net4257 sky130_fd_sc_hd__clkbuf_1
X_21268_ _00852_ _00853_ _00854_ VGND VGND VPWR VPWR _01283_ sky130_fd_sc_hd__o21a_1
Xwire4268 _04911_ VGND VGND VPWR VPWR net4268 sky130_fd_sc_hd__clkbuf_1
Xwire3523 net3524 VGND VGND VPWR VPWR net3523 sky130_fd_sc_hd__buf_1
Xwire4279 net4280 VGND VGND VPWR VPWR net4279 sky130_fd_sc_hd__clkbuf_1
X_23007_ net5141 net4571 VGND VGND VPWR VPWR _02877_ sky130_fd_sc_hd__nand2_1
Xwire2800 net2801 VGND VGND VPWR VPWR net2800 sky130_fd_sc_hd__buf_1
Xwire3545 net3549 VGND VGND VPWR VPWR net3545 sky130_fd_sc_hd__buf_1
X_20219_ net8953 net8119 net8 net8120 VGND VGND VPWR VPWR _12040_ sky130_fd_sc_hd__a31o_1
Xwire3556 net3557 VGND VGND VPWR VPWR net3556 sky130_fd_sc_hd__buf_1
Xwire2811 net2813 VGND VGND VPWR VPWR net2811 sky130_fd_sc_hd__buf_1
XFILLER_0_159_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2822 net2823 VGND VGND VPWR VPWR net2822 sky130_fd_sc_hd__buf_1
Xwire3567 net3568 VGND VGND VPWR VPWR net3567 sky130_fd_sc_hd__buf_1
X_21199_ _01144_ _01147_ _01213_ _01214_ VGND VGND VPWR VPWR _01215_ sky130_fd_sc_hd__o22a_1
Xwire2833 _07077_ VGND VGND VPWR VPWR net2833 sky130_fd_sc_hd__buf_1
Xwire3578 net3579 VGND VGND VPWR VPWR net3578 sky130_fd_sc_hd__buf_1
Xwire2844 net2845 VGND VGND VPWR VPWR net2844 sky130_fd_sc_hd__clkbuf_1
Xwire3589 _06989_ VGND VGND VPWR VPWR net3589 sky130_fd_sc_hd__clkbuf_1
Xwire2855 _06911_ VGND VGND VPWR VPWR net2855 sky130_fd_sc_hd__buf_1
Xwire2877 _06802_ VGND VGND VPWR VPWR net2877 sky130_fd_sc_hd__buf_1
Xwire2888 _06653_ VGND VGND VPWR VPWR net2888 sky130_fd_sc_hd__buf_1
Xwire2899 net2900 VGND VGND VPWR VPWR net2899 sky130_fd_sc_hd__buf_1
X_15760_ _07830_ VGND VGND VPWR VPWR _00218_ sky130_fd_sc_hd__clkbuf_1
X_24958_ pid_q.ki\[15\] _04732_ _04701_ VGND VGND VPWR VPWR _04733_ sky130_fd_sc_hd__mux2_1
X_12972_ _05243_ _05244_ _05202_ VGND VGND VPWR VPWR _05245_ sky130_fd_sc_hd__nor3b_1
X_14711_ matmul0.sin\[10\] net1908 net7456 VGND VGND VPWR VPWR _06853_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23909_ _03770_ _03673_ _03772_ VGND VGND VPWR VPWR _03773_ sky130_fd_sc_hd__a21o_1
X_15691_ net2724 _07761_ VGND VGND VPWR VPWR _07762_ sky130_fd_sc_hd__nor2_1
X_24889_ pid_q.ki\[11\] net2398 net3700 pid_q.kp\[11\] VGND VGND VPWR VPWR _04684_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_185_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17430_ svm0.delta\[14\] _09325_ _09273_ VGND VGND VPWR VPWR _09329_ sky130_fd_sc_hd__o21ai_1
X_14642_ net3697 VGND VGND VPWR VPWR _06805_ sky130_fd_sc_hd__clkbuf_1
X_17361_ net7377 net2579 net667 VGND VGND VPWR VPWR _09274_ sky130_fd_sc_hd__o21ai_1
X_14573_ net2884 _06749_ VGND VGND VPWR VPWR _06750_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19100_ net6204 net6178 VGND VGND VPWR VPWR _10937_ sky130_fd_sc_hd__and2b_1
X_13524_ _05793_ _05794_ VGND VGND VPWR VPWR _05795_ sky130_fd_sc_hd__xor2_1
X_16312_ _08359_ _08373_ _08374_ _08303_ VGND VGND VPWR VPWR _08375_ sky130_fd_sc_hd__a22o_1
Xmax_length6894 net6892 VGND VGND VPWR VPWR net6894 sky130_fd_sc_hd__buf_1
X_17292_ net7943 net7919 VGND VGND VPWR VPWR _09206_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19031_ _10860_ _10793_ VGND VGND VPWR VPWR _10868_ sky130_fd_sc_hd__xnor2_1
X_16243_ _08256_ _08295_ _08247_ VGND VGND VPWR VPWR _08307_ sky130_fd_sc_hd__o21a_1
X_13455_ _05699_ _05726_ _05725_ VGND VGND VPWR VPWR _05728_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_179_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16174_ net572 _08157_ _08231_ _08233_ VGND VGND VPWR VPWR _08239_ sky130_fd_sc_hd__o2bb2a_1
X_13386_ _05656_ _05657_ _05658_ _05558_ _05654_ VGND VGND VPWR VPWR _05659_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_51_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6160 net6161 VGND VGND VPWR VPWR net6160 sky130_fd_sc_hd__clkbuf_1
X_15125_ _07174_ _07198_ VGND VGND VPWR VPWR _07199_ sky130_fd_sc_hd__xnor2_1
Xfanout4630 pid_q.mult0.a\[7\] VGND VGND VPWR VPWR net4630 sky130_fd_sc_hd__buf_1
Xwire6171 net6169 VGND VGND VPWR VPWR net6171 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6193 cordic0.vec\[0\]\[8\] VGND VGND VPWR VPWR net6193 sky130_fd_sc_hd__buf_1
Xwire5470 pid_d.mult0.a\[11\] VGND VGND VPWR VPWR net5470 sky130_fd_sc_hd__clkbuf_1
Xwire5481 net5487 VGND VGND VPWR VPWR net5481 sky130_fd_sc_hd__buf_1
X_15056_ net2794 VGND VGND VPWR VPWR _07130_ sky130_fd_sc_hd__clkbuf_1
X_19933_ net6007 net2498 VGND VGND VPWR VPWR _11765_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5492 net5493 VGND VGND VPWR VPWR net5492 sky130_fd_sc_hd__buf_1
X_14007_ _06265_ _06268_ VGND VGND VPWR VPWR _06271_ sky130_fd_sc_hd__nand2_1
Xwire4780 net4781 VGND VGND VPWR VPWR net4780 sky130_fd_sc_hd__buf_1
X_19864_ net2097 _11696_ VGND VGND VPWR VPWR _11697_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18815_ _10657_ _10658_ net2132 VGND VGND VPWR VPWR _10659_ sky130_fd_sc_hd__o21a_1
X_19795_ net6008 net2100 _11628_ net6043 net3130 VGND VGND VPWR VPWR _11629_ sky130_fd_sc_hd__o221a_1
XFILLER_0_128_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18746_ _10589_ _10590_ VGND VGND VPWR VPWR _10591_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15958_ net2803 net2633 VGND VGND VPWR VPWR _08026_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14909_ net6614 net7423 matmul0.matmul_stage_inst.a\[8\] net6585 VGND VGND VPWR VPWR
+ _06983_ sky130_fd_sc_hd__a22o_1
X_18677_ _10521_ _10522_ _10475_ VGND VGND VPWR VPWR _10523_ sky130_fd_sc_hd__mux2_1
X_15889_ _07949_ _07957_ VGND VGND VPWR VPWR _07958_ sky130_fd_sc_hd__or2_1
X_17628_ _09482_ _09506_ _09494_ _09481_ _09508_ VGND VGND VPWR VPWR _09509_ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17559_ _09439_ _09440_ VGND VGND VPWR VPWR _09441_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20570_ _09008_ _12350_ _12352_ net3333 _12353_ VGND VGND VPWR VPWR _12354_ sky130_fd_sc_hd__o221a_1
XFILLER_0_128_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19229_ net6240 _11048_ net2519 net6139 VGND VGND VPWR VPWR _11066_ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2808 _07108_ VGND VGND VPWR VPWR net2808 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22240_ _02199_ _02244_ VGND VGND VPWR VPWR _02245_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_147_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22171_ pid_d.prev_error\[10\] pid_d.curr_error\[10\] VGND VGND VPWR VPWR _02177_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21122_ _01136_ _01137_ _00871_ VGND VGND VPWR VPWR _01138_ sky130_fd_sc_hd__a21oi_1
Xwire2107 _11157_ VGND VGND VPWR VPWR net2107 sky130_fd_sc_hd__buf_1
X_25930_ clknet_leaf_26_clk net9170 net8573 VGND VGND VPWR VPWR pid_d.prev_int\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_21053_ net3805 _01068_ VGND VGND VPWR VPWR _01069_ sky130_fd_sc_hd__or2_1
Xwire2118 net2119 VGND VGND VPWR VPWR net2118 sky130_fd_sc_hd__clkbuf_1
Xwire2129 _10368_ VGND VGND VPWR VPWR net2129 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_185_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1406 net1407 VGND VGND VPWR VPWR net1406 sky130_fd_sc_hd__clkbuf_2
X_20004_ net8975 net2122 net1444 _11834_ VGND VGND VPWR VPWR _00459_ sky130_fd_sc_hd__a31o_1
X_25861_ clknet_leaf_15_clk _00734_ net8617 VGND VGND VPWR VPWR pid_q.mult0.a\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1417 _11399_ VGND VGND VPWR VPWR net1417 sky130_fd_sc_hd__buf_1
XFILLER_0_185_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1428 _10674_ VGND VGND VPWR VPWR net1428 sky130_fd_sc_hd__buf_1
Xwire1439 _10344_ VGND VGND VPWR VPWR net1439 sky130_fd_sc_hd__buf_1
X_24812_ net5194 net5189 VGND VGND VPWR VPWR _04635_ sky130_fd_sc_hd__nand2_1
XFILLER_0_193_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25792_ clknet_leaf_32_clk _00665_ net8681 VGND VGND VPWR VPWR pid_q.curr_int\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_24743_ net1988 _04574_ VGND VGND VPWR VPWR _04575_ sky130_fd_sc_hd__nand2_1
X_21955_ net5858 net3787 _01962_ VGND VGND VPWR VPWR _01963_ sky130_fd_sc_hd__a21o_1
XFILLER_0_139_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20906_ net5906 _00865_ net5883 VGND VGND VPWR VPWR _00922_ sky130_fd_sc_hd__a21o_1
X_24674_ net9142 net1378 _04519_ VGND VGND VPWR VPWR _00689_ sky130_fd_sc_hd__a21o_1
X_21886_ net2068 _01794_ VGND VGND VPWR VPWR _01895_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_178_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6135 net6136 VGND VGND VPWR VPWR net6135 sky130_fd_sc_hd__buf_1
X_23625_ _03490_ _03491_ VGND VGND VPWR VPWR _03492_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_167_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20837_ net5731 net5615 VGND VGND VPWR VPWR _00853_ sky130_fd_sc_hd__nand2_1
XFILLER_0_193_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6168 net6164 VGND VGND VPWR VPWR net6168 sky130_fd_sc_hd__clkbuf_2
Xmax_length4700 net4692 VGND VGND VPWR VPWR net4700 sky130_fd_sc_hd__buf_1
X_23556_ _03336_ _03347_ _03335_ VGND VGND VPWR VPWR _03424_ sky130_fd_sc_hd__a21o_1
Xmax_length4722 net4723 VGND VGND VPWR VPWR net4722 sky130_fd_sc_hd__clkbuf_1
X_20768_ net5627 net5760 VGND VGND VPWR VPWR _12539_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire703 net704 VGND VGND VPWR VPWR net703 sky130_fd_sc_hd__buf_1
X_22507_ _02447_ _02500_ _02503_ _02507_ VGND VGND VPWR VPWR _02508_ sky130_fd_sc_hd__a211o_1
Xwire714 _10409_ VGND VGND VPWR VPWR net714 sky130_fd_sc_hd__buf_2
XFILLER_0_91_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire725 _07466_ VGND VGND VPWR VPWR net725 sky130_fd_sc_hd__clkbuf_1
X_23487_ _03241_ _03242_ _03355_ VGND VGND VPWR VPWR _03356_ sky130_fd_sc_hd__a21bo_1
Xwire736 _05123_ VGND VGND VPWR VPWR net736 sky130_fd_sc_hd__buf_1
XFILLER_0_52_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20699_ net6763 _09144_ _12313_ _09096_ VGND VGND VPWR VPWR _12473_ sky130_fd_sc_hd__a22o_1
Xmax_length323 net324 VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__clkbuf_1
Xwire747 net748 VGND VGND VPWR VPWR net747 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25226_ clknet_leaf_59_clk _00115_ net8694 VGND VGND VPWR VPWR svm0.vC\[14\] sky130_fd_sc_hd__dfrtp_1
X_13240_ _05441_ _05443_ _05512_ VGND VGND VPWR VPWR _05513_ sky130_fd_sc_hd__o21a_1
Xwire758 _01327_ VGND VGND VPWR VPWR net758 sky130_fd_sc_hd__buf_1
XFILLER_0_91_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire769 _09471_ VGND VGND VPWR VPWR net769 sky130_fd_sc_hd__clkbuf_1
X_22438_ _02438_ _02439_ VGND VGND VPWR VPWR _02440_ sky130_fd_sc_hd__xor2_1
XFILLER_0_134_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25157_ clknet_leaf_54_clk _00046_ net8727 VGND VGND VPWR VPWR pid_q.target\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13171_ _05442_ _05443_ VGND VGND VPWR VPWR _05444_ sky130_fd_sc_hd__xnor2_1
X_22369_ net5841 net5862 net2067 net2051 VGND VGND VPWR VPWR _02372_ sky130_fd_sc_hd__a31o_1
XFILLER_0_103_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4010 net4011 VGND VGND VPWR VPWR net4010 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4021 _09230_ VGND VGND VPWR VPWR net4021 sky130_fd_sc_hd__buf_1
XFILLER_0_62_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24108_ net5059 net5028 VGND VGND VPWR VPWR _03970_ sky130_fd_sc_hd__nand2_1
Xwire4032 net4033 VGND VGND VPWR VPWR net4032 sky130_fd_sc_hd__buf_1
X_25088_ net1627 _04832_ net1633 VGND VGND VPWR VPWR _04833_ sky130_fd_sc_hd__a21o_1
Xwire4043 net4044 VGND VGND VPWR VPWR net4043 sky130_fd_sc_hd__buf_1
Xwire4054 _08900_ VGND VGND VPWR VPWR net4054 sky130_fd_sc_hd__buf_1
Xwire3320 net3321 VGND VGND VPWR VPWR net3320 sky130_fd_sc_hd__clkbuf_1
Xwire4065 net4066 VGND VGND VPWR VPWR net4065 sky130_fd_sc_hd__clkbuf_1
Xwire3331 _08985_ VGND VGND VPWR VPWR net3331 sky130_fd_sc_hd__buf_1
X_24039_ _03900_ _03901_ VGND VGND VPWR VPWR _03902_ sky130_fd_sc_hd__xor2_1
X_16930_ net6416 _08890_ _08892_ _08893_ VGND VGND VPWR VPWR _08894_ sky130_fd_sc_hd__a22o_1
Xwire4076 _07601_ VGND VGND VPWR VPWR net4076 sky130_fd_sc_hd__buf_1
Xwire3342 _08948_ VGND VGND VPWR VPWR net3342 sky130_fd_sc_hd__buf_1
Xwire4087 net4088 VGND VGND VPWR VPWR net4087 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3353 net3354 VGND VGND VPWR VPWR net3353 sky130_fd_sc_hd__buf_1
Xwire4098 net4099 VGND VGND VPWR VPWR net4098 sky130_fd_sc_hd__buf_1
Xwire3364 _08826_ VGND VGND VPWR VPWR net3364 sky130_fd_sc_hd__clkbuf_1
Xwire2630 _07933_ VGND VGND VPWR VPWR net2630 sky130_fd_sc_hd__buf_1
Xwire3375 net3376 VGND VGND VPWR VPWR net3375 sky130_fd_sc_hd__clkbuf_1
Xwire3386 _08647_ VGND VGND VPWR VPWR net3386 sky130_fd_sc_hd__buf_1
Xwire2641 net2642 VGND VGND VPWR VPWR net2641 sky130_fd_sc_hd__buf_1
X_16861_ _08820_ _08821_ _08822_ _08823_ net4062 _08825_ VGND VGND VPWR VPWR _08826_
+ sky130_fd_sc_hd__mux4_1
Xwire2652 _07761_ VGND VGND VPWR VPWR net2652 sky130_fd_sc_hd__buf_1
XFILLER_0_74_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3397 _07684_ VGND VGND VPWR VPWR net3397 sky130_fd_sc_hd__buf_1
Xwire2663 net2664 VGND VGND VPWR VPWR net2663 sky130_fd_sc_hd__clkbuf_1
X_18600_ _10445_ _10446_ net6793 _10447_ VGND VGND VPWR VPWR _10448_ sky130_fd_sc_hd__o2bb2a_1
Xwire2674 net2675 VGND VGND VPWR VPWR net2674 sky130_fd_sc_hd__clkbuf_1
Xwire1940 net1941 VGND VGND VPWR VPWR net1940 sky130_fd_sc_hd__buf_1
X_15812_ _07785_ _07790_ VGND VGND VPWR VPWR _07882_ sky130_fd_sc_hd__nor2_1
Xwire2685 net2686 VGND VGND VPWR VPWR net2685 sky130_fd_sc_hd__buf_1
X_19580_ _11405_ _11416_ VGND VGND VPWR VPWR _11417_ sky130_fd_sc_hd__xnor2_2
Xwire2696 _07489_ VGND VGND VPWR VPWR net2696 sky130_fd_sc_hd__buf_1
Xwire1962 net1965 VGND VGND VPWR VPWR net1962 sky130_fd_sc_hd__buf_1
X_16792_ net7577 matmul0.a\[15\] net3373 VGND VGND VPWR VPWR _08786_ sky130_fd_sc_hd__mux2_1
Xwire1973 _04924_ VGND VGND VPWR VPWR net1973 sky130_fd_sc_hd__buf_1
Xwire1984 net1986 VGND VGND VPWR VPWR net1984 sky130_fd_sc_hd__clkbuf_1
X_18531_ net1197 _10379_ VGND VGND VPWR VPWR _10380_ sky130_fd_sc_hd__xnor2_2
Xwire1995 _04787_ VGND VGND VPWR VPWR net1995 sky130_fd_sc_hd__buf_1
X_12955_ _05002_ _05226_ VGND VGND VPWR VPWR _05228_ sky130_fd_sc_hd__or2_1
X_15743_ _07813_ VGND VGND VPWR VPWR _07814_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18462_ _10310_ _10311_ net3284 VGND VGND VPWR VPWR _10312_ sky130_fd_sc_hd__mux2_1
X_12886_ _05155_ _05158_ VGND VGND VPWR VPWR _05159_ sky130_fd_sc_hd__xnor2_2
X_15674_ net2701 net3526 VGND VGND VPWR VPWR _07745_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17413_ svm0.delta\[10\] _09312_ VGND VGND VPWR VPWR _09316_ sky130_fd_sc_hd__or2_1
X_14625_ net6448 _06541_ VGND VGND VPWR VPWR _06794_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18393_ net1773 _10243_ VGND VGND VPWR VPWR _10244_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17344_ net4016 VGND VGND VPWR VPWR _09258_ sky130_fd_sc_hd__buf_1
X_14556_ _06731_ _06732_ VGND VGND VPWR VPWR _06734_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13507_ _05778_ VGND VGND VPWR VPWR _05779_ sky130_fd_sc_hd__clkbuf_2
X_17275_ net2982 net157 net2157 net9232 VGND VGND VPWR VPWR _00369_ sky130_fd_sc_hd__a22o_1
X_14487_ net9051 net832 net1292 _06671_ VGND VGND VPWR VPWR _00104_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19014_ net6181 _10850_ VGND VGND VPWR VPWR _10851_ sky130_fd_sc_hd__xnor2_4
X_13438_ _05708_ _05710_ VGND VGND VPWR VPWR _05711_ sky130_fd_sc_hd__xnor2_1
X_16226_ net2206 net1513 VGND VGND VPWR VPWR _08291_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16157_ _08212_ _08222_ VGND VGND VPWR VPWR _08223_ sky130_fd_sc_hd__xor2_1
X_13369_ svm0.vC\[15\] net2378 _05641_ net3028 VGND VGND VPWR VPWR _05642_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15108_ _07176_ _07181_ VGND VGND VPWR VPWR _07182_ sky130_fd_sc_hd__xor2_1
X_16088_ _08068_ net1257 _08154_ VGND VGND VPWR VPWR _08155_ sky130_fd_sc_hd__o21a_1
Xfanout4482 net4489 VGND VGND VPWR VPWR net4482 sky130_fd_sc_hd__buf_1
X_19916_ net6110 net3149 _11686_ _11747_ VGND VGND VPWR VPWR _11748_ sky130_fd_sc_hd__o31a_1
X_15039_ net4195 net4193 net4205 net4204 VGND VGND VPWR VPWR _07113_ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19847_ _11642_ _11678_ _11679_ VGND VGND VPWR VPWR _11680_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19778_ net1767 _11610_ _11611_ _11612_ VGND VGND VPWR VPWR _00455_ sky130_fd_sc_hd__a31o_1
XFILLER_0_155_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18729_ net6877 _10534_ VGND VGND VPWR VPWR _10574_ sky130_fd_sc_hd__or2_1
XFILLER_0_189_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21740_ net5686 net5551 VGND VGND VPWR VPWR _01750_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21671_ _01571_ _01573_ VGND VGND VPWR VPWR _01682_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8309 net8310 VGND VGND VPWR VPWR net8309 sky130_fd_sc_hd__clkbuf_1
X_23410_ _03269_ _03279_ VGND VGND VPWR VPWR _03280_ sky130_fd_sc_hd__xor2_1
XFILLER_0_15_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length4018 net4019 VGND VGND VPWR VPWR net4018 sky130_fd_sc_hd__buf_1
X_20622_ net2191 _12402_ net8054 VGND VGND VPWR VPWR _12403_ sky130_fd_sc_hd__o21a_1
XFILLER_0_191_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24390_ net588 net587 VGND VGND VPWR VPWR _04249_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7619 net7614 VGND VGND VPWR VPWR net7619 sky130_fd_sc_hd__buf_1
XFILLER_0_184_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23341_ _03209_ _03210_ VGND VGND VPWR VPWR _03211_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20553_ net3854 net3853 net3335 VGND VGND VPWR VPWR _12338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6907 net6908 VGND VGND VPWR VPWR net6907 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6929 net6930 VGND VGND VPWR VPWR net6929 sky130_fd_sc_hd__buf_1
X_23272_ _03134_ _03141_ VGND VGND VPWR VPWR _03142_ sky130_fd_sc_hd__xnor2_1
Xmax_length2627 _07936_ VGND VGND VPWR VPWR net2627 sky130_fd_sc_hd__buf_1
X_20484_ net1237 net2087 net3170 VGND VGND VPWR VPWR _12273_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_171_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25011_ net4466 net1631 net2394 _04766_ VGND VGND VPWR VPWR _00779_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22223_ net5785 net5800 VGND VGND VPWR VPWR _02228_ sky130_fd_sc_hd__or2_2
XFILLER_0_89_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22154_ net1710 _02057_ VGND VGND VPWR VPWR _02160_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21105_ _01117_ _01118_ _01120_ VGND VGND VPWR VPWR _01121_ sky130_fd_sc_hd__a21oi_1
X_22085_ _02090_ _02091_ VGND VGND VPWR VPWR _02092_ sky130_fd_sc_hd__and2b_1
XFILLER_0_100_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_1__f_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_4_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_25913_ clknet_leaf_66_clk _00786_ net8659 VGND VGND VPWR VPWR pid_q.out\[9\] sky130_fd_sc_hd__dfrtp_1
X_21036_ _01050_ _01051_ VGND VGND VPWR VPWR _01052_ sky130_fd_sc_hd__and2b_1
Xwire1203 _10343_ VGND VGND VPWR VPWR net1203 sky130_fd_sc_hd__buf_1
Xwire1225 net1226 VGND VGND VPWR VPWR net1225 sky130_fd_sc_hd__clkbuf_1
Xwire1236 _08917_ VGND VGND VPWR VPWR net1236 sky130_fd_sc_hd__clkbuf_1
X_25844_ clknet_leaf_38_clk _00717_ net8747 VGND VGND VPWR VPWR pid_q.mult0.b\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1247 _08419_ VGND VGND VPWR VPWR net1247 sky130_fd_sc_hd__buf_1
Xwire1258 net1259 VGND VGND VPWR VPWR net1258 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1269 _07662_ VGND VGND VPWR VPWR net1269 sky130_fd_sc_hd__buf_1
XFILLER_0_92_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22987_ _02861_ VGND VGND VPWR VPWR _00660_ sky130_fd_sc_hd__clkbuf_1
X_25775_ clknet_leaf_64_clk _00648_ net8662 VGND VGND VPWR VPWR matmul0.beta_pass\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12740_ net7916 net1342 VGND VGND VPWR VPWR _05013_ sky130_fd_sc_hd__nand2_1
XFILLER_0_195_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24726_ _04558_ _04559_ net1988 VGND VGND VPWR VPWR _04560_ sky130_fd_sc_hd__o21a_1
X_21938_ _01942_ _01945_ VGND VGND VPWR VPWR _01946_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_167_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24657_ pid_q.curr_error\[0\] _00011_ net1374 VGND VGND VPWR VPWR _04511_ sky130_fd_sc_hd__and3_1
X_12671_ _04942_ _04943_ net7853 net1615 VGND VGND VPWR VPWR _04944_ sky130_fd_sc_hd__o211a_1
X_21869_ net1047 _01877_ VGND VGND VPWR VPWR _01878_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_127_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14410_ _06611_ matmul0.b_in\[4\] net897 VGND VGND VPWR VPWR _06612_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23608_ pid_q.prev_error\[1\] net5168 pid_q.prev_error\[0\] pid_q.curr_error\[0\]
+ VGND VGND VPWR VPWR _03476_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_139_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15390_ _07453_ _07327_ net990 VGND VGND VPWR VPWR _07464_ sky130_fd_sc_hd__mux2_1
Xwire8821 net8822 VGND VGND VPWR VPWR net8821 sky130_fd_sc_hd__buf_1
X_24588_ _04441_ net631 VGND VGND VPWR VPWR _04444_ sky130_fd_sc_hd__xnor2_1
Xmax_length5253 net5254 VGND VGND VPWR VPWR net5253 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8832 net8833 VGND VGND VPWR VPWR net8832 sky130_fd_sc_hd__clkbuf_1
Xwire8843 net8814 VGND VGND VPWR VPWR net8843 sky130_fd_sc_hd__clkbuf_1
Xmax_length4530 net4531 VGND VGND VPWR VPWR net4530 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8854 net8855 VGND VGND VPWR VPWR net8854 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire500 net501 VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__clkbuf_1
X_14341_ net7309 net1299 net2896 pid_d.out\[5\] _06557_ VGND VGND VPWR VPWR _06558_
+ sky130_fd_sc_hd__a221o_1
X_23539_ _03405_ _03406_ VGND VGND VPWR VPWR _03407_ sky130_fd_sc_hd__or2b_1
Xwire8865 net8862 VGND VGND VPWR VPWR net8865 sky130_fd_sc_hd__buf_1
XFILLER_0_163_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire511 _03846_ VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__buf_1
Xwire8876 net8877 VGND VGND VPWR VPWR net8876 sky130_fd_sc_hd__buf_1
Xwire522 _02106_ VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__buf_1
XFILLER_0_80_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire533 _05847_ VGND VGND VPWR VPWR net533 sky130_fd_sc_hd__buf_1
XFILLER_0_150_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire544 net545 VGND VGND VPWR VPWR net544 sky130_fd_sc_hd__clkbuf_1
Xwire8898 net8895 VGND VGND VPWR VPWR net8898 sky130_fd_sc_hd__buf_1
X_17060_ _08977_ _09018_ VGND VGND VPWR VPWR _09019_ sky130_fd_sc_hd__or2_1
X_14272_ net3657 VGND VGND VPWR VPWR _06516_ sky130_fd_sc_hd__clkbuf_1
Xwire555 net556 VGND VGND VPWR VPWR net555 sky130_fd_sc_hd__buf_1
XFILLER_0_69_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3873 _11164_ VGND VGND VPWR VPWR net3873 sky130_fd_sc_hd__clkbuf_1
Xwire566 _01331_ VGND VGND VPWR VPWR net566 sky130_fd_sc_hd__clkbuf_1
Xwire577 _05835_ VGND VGND VPWR VPWR net577 sky130_fd_sc_hd__buf_1
XFILLER_0_122_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16011_ _07999_ _08001_ VGND VGND VPWR VPWR _08079_ sky130_fd_sc_hd__and2b_1
XFILLER_0_33_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13223_ net7640 net2339 net1967 VGND VGND VPWR VPWR _05496_ sky130_fd_sc_hd__and3_1
Xwire588 _04246_ VGND VGND VPWR VPWR net588 sky130_fd_sc_hd__buf_1
X_25209_ clknet_leaf_62_clk _00098_ net8672 VGND VGND VPWR VPWR matmul0.b_in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire599 _01903_ VGND VGND VPWR VPWR net599 sky130_fd_sc_hd__buf_1
XFILLER_0_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13154_ _05424_ _05425_ _05416_ VGND VGND VPWR VPWR _05427_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13085_ _05270_ _05271_ _05272_ _05273_ VGND VGND VPWR VPWR _05358_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_29_Left_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17962_ net7090 _09620_ VGND VGND VPWR VPWR _09813_ sky130_fd_sc_hd__nor2_1
Xwire3150 net3151 VGND VGND VPWR VPWR net3150 sky130_fd_sc_hd__buf_1
X_19701_ _11380_ _11384_ _11386_ VGND VGND VPWR VPWR _11537_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16913_ _08862_ net6371 _08874_ _08875_ _08876_ VGND VGND VPWR VPWR _08877_ sky130_fd_sc_hd__a2111oi_1
Xwire3161 _11273_ VGND VGND VPWR VPWR net3161 sky130_fd_sc_hd__clkbuf_2
Xwire3172 net3173 VGND VGND VPWR VPWR net3172 sky130_fd_sc_hd__clkbuf_1
Xwire3183 _11027_ VGND VGND VPWR VPWR net3183 sky130_fd_sc_hd__buf_1
X_17893_ _09742_ net2553 _09695_ VGND VGND VPWR VPWR _09744_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3194 net3195 VGND VGND VPWR VPWR net3194 sky130_fd_sc_hd__clkbuf_1
Xwire2460 net2461 VGND VGND VPWR VPWR net2460 sky130_fd_sc_hd__buf_1
Xwire2471 _02301_ VGND VGND VPWR VPWR net2471 sky130_fd_sc_hd__dlymetal6s2s_1
X_19632_ net1749 net2101 VGND VGND VPWR VPWR _11469_ sky130_fd_sc_hd__xnor2_1
X_16844_ net6422 matmul0.sin\[10\] net3365 VGND VGND VPWR VPWR _08813_ sky130_fd_sc_hd__mux2_1
Xwire2482 _00886_ VGND VGND VPWR VPWR net2482 sky130_fd_sc_hd__buf_1
Xwire2493 _11893_ VGND VGND VPWR VPWR net2493 sky130_fd_sc_hd__buf_1
XFILLER_0_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1770 net1771 VGND VGND VPWR VPWR net1770 sky130_fd_sc_hd__buf_1
X_19563_ _11076_ _11075_ net3177 VGND VGND VPWR VPWR _11400_ sky130_fd_sc_hd__mux2_1
Xwire1781 _09658_ VGND VGND VPWR VPWR net1781 sky130_fd_sc_hd__buf_1
XFILLER_0_189_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16775_ matmul0.a_in\[7\] matmul0.a\[7\] _08770_ VGND VGND VPWR VPWR _08777_ sky130_fd_sc_hd__mux2_1
Xwire1792 net1793 VGND VGND VPWR VPWR net1792 sky130_fd_sc_hd__clkbuf_1
X_13987_ _06192_ _06194_ _06193_ VGND VGND VPWR VPWR _06252_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_34_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18514_ net3331 _09791_ _10303_ net6970 VGND VGND VPWR VPWR _10363_ sky130_fd_sc_hd__a22o_1
X_15726_ _07794_ _07796_ VGND VGND VPWR VPWR _07797_ sky130_fd_sc_hd__xnor2_1
X_12938_ _05152_ _05210_ VGND VGND VPWR VPWR _05211_ sky130_fd_sc_hd__xnor2_1
X_19494_ _11328_ _11330_ VGND VGND VPWR VPWR _11331_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18445_ net7017 net7099 VGND VGND VPWR VPWR _10295_ sky130_fd_sc_hd__nor2_1
X_15657_ _07584_ _07588_ _07728_ VGND VGND VPWR VPWR _07729_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_38_Left_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12869_ _05126_ net791 VGND VGND VPWR VPWR _05142_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14608_ _06768_ _06777_ VGND VGND VPWR VPWR _06781_ sky130_fd_sc_hd__and2_1
X_18376_ net3936 _09634_ VGND VGND VPWR VPWR _10227_ sky130_fd_sc_hd__nand2_1
X_15588_ _07651_ _07659_ VGND VGND VPWR VPWR _07660_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17327_ _09206_ _09240_ VGND VGND VPWR VPWR _09241_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14539_ net5247 _06710_ _06711_ VGND VGND VPWR VPWR _06718_ sky130_fd_sc_hd__nor3_1
XFILLER_0_172_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17258_ net2960 net154 _09189_ net9096 VGND VGND VPWR VPWR _00356_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_183_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16209_ _08270_ _08273_ VGND VGND VPWR VPWR _08274_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17189_ net2932 _09138_ net4245 VGND VGND VPWR VPWR _09140_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_47_Left_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22910_ _02183_ _02797_ _02801_ VGND VGND VPWR VPWR _02802_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23890_ _03750_ _03752_ VGND VGND VPWR VPWR _03755_ sky130_fd_sc_hd__nor2_1
X_22841_ net4335 _02739_ _02740_ net415 net4354 VGND VGND VPWR VPWR _02741_ sky130_fd_sc_hd__a32o_1
XFILLER_0_155_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25560_ clknet_leaf_115_clk _00433_ net8335 VGND VGND VPWR VPWR cordic0.gm0.iter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_22772_ pid_d.ki\[15\] _02692_ net2039 VGND VGND VPWR VPWR _02693_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_56_Left_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24511_ _04272_ _04276_ _04367_ VGND VGND VPWR VPWR _04368_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_66_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21723_ net4358 _01732_ _01733_ VGND VGND VPWR VPWR _01734_ sky130_fd_sc_hd__and3_1
X_25491_ clknet_leaf_47_clk _00371_ net8775 VGND VGND VPWR VPWR svm0.tA\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8106 net83 VGND VGND VPWR VPWR net8106 sky130_fd_sc_hd__clkbuf_1
X_24442_ net4516 net4844 VGND VGND VPWR VPWR _04300_ sky130_fd_sc_hd__nand2_1
Xwire8117 net81 VGND VGND VPWR VPWR net8117 sky130_fd_sc_hd__clkbuf_1
X_21654_ _01661_ _01664_ VGND VGND VPWR VPWR _01665_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_163_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8128 net8129 VGND VGND VPWR VPWR net8128 sky130_fd_sc_hd__clkbuf_1
Xwire8139 net8140 VGND VGND VPWR VPWR net8139 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7405 matmul0.matmul_stage_inst.c\[11\] VGND VGND VPWR VPWR net7405 sky130_fd_sc_hd__clkbuf_1
X_20605_ _12385_ net1396 VGND VGND VPWR VPWR _12386_ sky130_fd_sc_hd__nor2_1
Xfanout6609 net6623 VGND VGND VPWR VPWR net6609 sky130_fd_sc_hd__clkbuf_1
X_24373_ net4804 _04126_ _04230_ VGND VGND VPWR VPWR _04232_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire7416 matmul0.matmul_stage_inst.c\[4\] VGND VGND VPWR VPWR net7416 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21585_ _01472_ _01474_ _01596_ VGND VGND VPWR VPWR _01597_ sky130_fd_sc_hd__o21a_1
Xwire7427 net7428 VGND VGND VPWR VPWR net7427 sky130_fd_sc_hd__clkbuf_1
Xmax_length3125 _11754_ VGND VGND VPWR VPWR net3125 sky130_fd_sc_hd__clkbuf_2
Xwire6704 svm0.counter\[11\] VGND VGND VPWR VPWR net6704 sky130_fd_sc_hd__buf_1
Xwire7449 net7452 VGND VGND VPWR VPWR net7449 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6715 net6716 VGND VGND VPWR VPWR net6715 sky130_fd_sc_hd__clkbuf_1
X_23324_ net4850 net4771 VGND VGND VPWR VPWR _03194_ sky130_fd_sc_hd__nand2_1
X_20536_ _12305_ _12320_ _12309_ VGND VGND VPWR VPWR _12322_ sky130_fd_sc_hd__and3_1
Xwire6726 svm0.counter\[6\] VGND VGND VPWR VPWR net6726 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6737 svm0.counter\[1\] VGND VGND VPWR VPWR net6737 sky130_fd_sc_hd__buf_1
Xwire6748 net6749 VGND VGND VPWR VPWR net6748 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23255_ net2430 _03100_ VGND VGND VPWR VPWR _03125_ sky130_fd_sc_hd__xor2_1
X_20467_ _12252_ _12256_ _12257_ VGND VGND VPWR VPWR _12258_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_65_Left_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22206_ net5489 net5675 VGND VGND VPWR VPWR _02211_ sky130_fd_sc_hd__nand2_1
X_23186_ _03054_ _03055_ VGND VGND VPWR VPWR _03056_ sky130_fd_sc_hd__xor2_2
Xmax_length1767 net1768 VGND VGND VPWR VPWR net1767 sky130_fd_sc_hd__buf_1
X_20398_ net6458 _12195_ VGND VGND VPWR VPWR _12196_ sky130_fd_sc_hd__nor2_1
X_22137_ _02039_ _02041_ _02142_ VGND VGND VPWR VPWR _02143_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22068_ net1716 _01967_ VGND VGND VPWR VPWR _02075_ sky130_fd_sc_hd__nor2_1
Xwire1000 _05446_ VGND VGND VPWR VPWR net1000 sky130_fd_sc_hd__buf_1
Xwire1011 _04539_ VGND VGND VPWR VPWR net1011 sky130_fd_sc_hd__buf_1
Xwire1022 net1023 VGND VGND VPWR VPWR net1022 sky130_fd_sc_hd__clkbuf_1
X_13910_ net7632 net1583 _06175_ net1965 VGND VGND VPWR VPWR _06176_ sky130_fd_sc_hd__o22a_1
X_21019_ _01033_ _01034_ VGND VGND VPWR VPWR _01035_ sky130_fd_sc_hd__xnor2_1
Xwire1033 net1034 VGND VGND VPWR VPWR net1033 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1044 _01983_ VGND VGND VPWR VPWR net1044 sky130_fd_sc_hd__buf_1
X_14890_ net4221 net4219 VGND VGND VPWR VPWR _06964_ sky130_fd_sc_hd__nor2_1
Xwire1055 _11951_ VGND VGND VPWR VPWR net1055 sky130_fd_sc_hd__buf_1
Xwire1066 net1067 VGND VGND VPWR VPWR net1066 sky130_fd_sc_hd__buf_1
X_13841_ _06057_ _06058_ _06106_ VGND VGND VPWR VPWR _06108_ sky130_fd_sc_hd__a21oi_1
X_25827_ clknet_leaf_36_clk _00700_ net8748 VGND VGND VPWR VPWR pid_q.curr_error\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1077 _08992_ VGND VGND VPWR VPWR net1077 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1088 _08219_ VGND VGND VPWR VPWR net1088 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_74_Left_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1099 net1100 VGND VGND VPWR VPWR net1099 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_57_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13772_ _06033_ _06034_ _06039_ VGND VGND VPWR VPWR _06040_ sky130_fd_sc_hd__a21oi_1
X_16560_ _08529_ _08572_ net1243 VGND VGND VPWR VPWR _08619_ sky130_fd_sc_hd__a21bo_1
X_25758_ clknet_leaf_27_clk _00631_ net8645 VGND VGND VPWR VPWR pid_d.out_valid sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15511_ _07576_ _07583_ VGND VGND VPWR VPWR _07584_ sky130_fd_sc_hd__xnor2_2
X_24709_ net5299 net8028 VGND VGND VPWR VPWR _04545_ sky130_fd_sc_hd__and2b_1
X_12723_ _04986_ _04987_ VGND VGND VPWR VPWR _04996_ sky130_fd_sc_hd__and2_1
Xfanout8501 net8505 VGND VGND VPWR VPWR net8501 sky130_fd_sc_hd__clkbuf_1
X_16491_ _08522_ net975 VGND VGND VPWR VPWR _08551_ sky130_fd_sc_hd__nand2_1
XFILLER_0_167_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25689_ clknet_leaf_3_clk _00562_ net8569 VGND VGND VPWR VPWR pid_d.curr_error\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_18230_ net7063 _10034_ _10038_ VGND VGND VPWR VPWR _10081_ sky130_fd_sc_hd__mux2_1
X_12654_ net7797 _04924_ _04926_ VGND VGND VPWR VPWR _04927_ sky130_fd_sc_hd__and3_1
Xfanout7800 net7813 VGND VGND VPWR VPWR net7800 sky130_fd_sc_hd__buf_1
X_15442_ net4083 net4081 VGND VGND VPWR VPWR _07516_ sky130_fd_sc_hd__nor2_1
XFILLER_0_183_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8640 net8641 VGND VGND VPWR VPWR net8640 sky130_fd_sc_hd__clkbuf_1
Xfanout7844 net7857 VGND VGND VPWR VPWR net7844 sky130_fd_sc_hd__clkbuf_1
X_18161_ _10010_ _10011_ VGND VGND VPWR VPWR _10012_ sky130_fd_sc_hd__xnor2_1
X_12585_ net3716 VGND VGND VPWR VPWR _04870_ sky130_fd_sc_hd__clkbuf_1
Xwire8651 net8652 VGND VGND VPWR VPWR net8651 sky130_fd_sc_hd__buf_1
XFILLER_0_52_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15373_ _07443_ _07445_ VGND VGND VPWR VPWR _07447_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8662 net8661 VGND VGND VPWR VPWR net8662 sky130_fd_sc_hd__clkbuf_2
X_17112_ net1813 VGND VGND VPWR VPWR _09068_ sky130_fd_sc_hd__buf_1
Xwire7950 net7951 VGND VGND VPWR VPWR net7950 sky130_fd_sc_hd__clkbuf_1
Xfanout7888 svm0.periodTop\[2\] VGND VGND VPWR VPWR net7888 sky130_fd_sc_hd__buf_1
Xwire330 _03945_ VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14324_ net8271 net3642 VGND VGND VPWR VPWR _06545_ sky130_fd_sc_hd__and2_1
Xwire8695 net8692 VGND VGND VPWR VPWR net8695 sky130_fd_sc_hd__buf_1
XFILLER_0_135_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire341 _02172_ VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__clkbuf_1
X_18092_ _09901_ _09942_ VGND VGND VPWR VPWR _09943_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7961 net7962 VGND VGND VPWR VPWR net7961 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_108_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire352 _10693_ VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_83_Left_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire7972 net7973 VGND VGND VPWR VPWR net7972 sky130_fd_sc_hd__clkbuf_1
Xwire363 net364 VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__clkbuf_1
Xwire7983 net7984 VGND VGND VPWR VPWR net7983 sky130_fd_sc_hd__clkbuf_1
Xwire374 net375 VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__clkbuf_1
Xwire7994 net7995 VGND VGND VPWR VPWR net7994 sky130_fd_sc_hd__clkbuf_1
X_17043_ net3328 _09002_ VGND VGND VPWR VPWR _09003_ sky130_fd_sc_hd__nor2_1
X_14255_ net2285 net1554 VGND VGND VPWR VPWR _00034_ sky130_fd_sc_hd__nand2_1
Xwire385 net386 VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__buf_1
Xwire396 net397 VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__buf_1
XFILLER_0_187_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13206_ _05477_ _05478_ VGND VGND VPWR VPWR _05479_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14186_ net1304 VGND VGND VPWR VPWR _06446_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13137_ _05388_ _05389_ _05391_ _05392_ VGND VGND VPWR VPWR _05410_ sky130_fd_sc_hd__a211o_1
X_18994_ _10811_ _10830_ net6356 VGND VGND VPWR VPWR _10831_ sky130_fd_sc_hd__a21oi_1
X_13068_ _05339_ _05340_ VGND VGND VPWR VPWR _05341_ sky130_fd_sc_hd__xnor2_1
X_17945_ net6978 net6951 VGND VGND VPWR VPWR _09796_ sky130_fd_sc_hd__nor2_1
X_17876_ _09725_ net1780 net2141 _09726_ VGND VGND VPWR VPWR _09727_ sky130_fd_sc_hd__a22o_1
Xwire2290 _06502_ VGND VGND VPWR VPWR net2290 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19615_ _11379_ _11451_ VGND VGND VPWR VPWR _11452_ sky130_fd_sc_hd__or2b_1
X_16827_ _08804_ VGND VGND VPWR VPWR _00311_ sky130_fd_sc_hd__clkbuf_1
X_19546_ net6116 net6097 VGND VGND VPWR VPWR _11383_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16758_ net7553 matmul0.b\[15\] net3382 VGND VGND VPWR VPWR _08768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15709_ net3454 VGND VGND VPWR VPWR _07780_ sky130_fd_sc_hd__clkbuf_1
X_19477_ _10985_ net3895 _11265_ VGND VGND VPWR VPWR _11314_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16689_ _08718_ _08719_ VGND VGND VPWR VPWR _08720_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18428_ net3929 net6801 VGND VGND VPWR VPWR _10278_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18359_ _10207_ _10208_ _10209_ VGND VGND VPWR VPWR _10210_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_161_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21370_ _01380_ _01383_ VGND VGND VPWR VPWR _01384_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20321_ _12102_ _12113_ _12123_ _12124_ VGND VGND VPWR VPWR _12125_ sky130_fd_sc_hd__a31o_1
XFILLER_0_82_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23040_ net5087 net4647 VGND VGND VPWR VPWR _02910_ sky130_fd_sc_hd__nand2_1
X_20252_ net8121 _12065_ VGND VGND VPWR VPWR _12066_ sky130_fd_sc_hd__nor2_1
Xwire3908 net3909 VGND VGND VPWR VPWR net3908 sky130_fd_sc_hd__buf_1
X_20183_ net6004 _12006_ _12008_ VGND VGND VPWR VPWR _12009_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24991_ _04750_ VGND VGND VPWR VPWR _00775_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23942_ net3741 _03805_ VGND VGND VPWR VPWR _03806_ sky130_fd_sc_hd__nor2_1
X_23873_ net4674 net4704 _03373_ VGND VGND VPWR VPWR _03738_ sky130_fd_sc_hd__nand3_1
XFILLER_0_168_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25612_ clknet_leaf_111_clk _00485_ net8349 VGND VGND VPWR VPWR cordic0.slte0.opA\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_22824_ net4360 net560 _02725_ net4335 net2463 VGND VGND VPWR VPWR _02726_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22755_ _02681_ VGND VGND VPWR VPWR _00608_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25543_ clknet_leaf_32_clk _00423_ net8679 VGND VGND VPWR VPWR pid_q.prev_int\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_165_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21706_ _01708_ _01716_ VGND VGND VPWR VPWR _01717_ sky130_fd_sc_hd__xor2_1
X_25474_ clknet_leaf_47_clk _00354_ net8776 VGND VGND VPWR VPWR svm0.tB\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22686_ _02632_ VGND VGND VPWR VPWR _00588_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout7118 net7127 VGND VGND VPWR VPWR net7118 sky130_fd_sc_hd__buf_1
X_24425_ net4485 _04282_ VGND VGND VPWR VPWR _04283_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7202 matmul0.alpha_pass\[15\] VGND VGND VPWR VPWR net7202 sky130_fd_sc_hd__buf_1
X_21637_ _01646_ _01647_ VGND VGND VPWR VPWR _01648_ sky130_fd_sc_hd__xnor2_1
Xwire7213 matmul0.alpha_pass\[14\] VGND VGND VPWR VPWR net7213 sky130_fd_sc_hd__buf_1
XFILLER_0_34_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7235 net7236 VGND VGND VPWR VPWR net7235 sky130_fd_sc_hd__clkbuf_1
X_24356_ net4937 _03605_ _04078_ net3742 VGND VGND VPWR VPWR _04215_ sky130_fd_sc_hd__a31oi_1
Xwire7246 net7247 VGND VGND VPWR VPWR net7246 sky130_fd_sc_hd__buf_1
Xwire7257 net7258 VGND VGND VPWR VPWR net7257 sky130_fd_sc_hd__dlymetal6s2s_1
X_21568_ _01577_ _01579_ VGND VGND VPWR VPWR _01580_ sky130_fd_sc_hd__xor2_1
Xwire7268 net7269 VGND VGND VPWR VPWR net7268 sky130_fd_sc_hd__clkbuf_1
Xwire6534 net6531 VGND VGND VPWR VPWR net6534 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_185_Right_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23307_ _02968_ _03175_ _02965_ VGND VGND VPWR VPWR _03177_ sky130_fd_sc_hd__a21bo_1
X_20519_ _12304_ _12305_ VGND VGND VPWR VPWR _12306_ sky130_fd_sc_hd__nand2_1
Xwire6545 net6544 VGND VGND VPWR VPWR net6545 sky130_fd_sc_hd__buf_1
X_24287_ net4993 net4959 net4937 net4484 VGND VGND VPWR VPWR _04147_ sky130_fd_sc_hd__o31ai_1
Xwire5811 net5815 VGND VGND VPWR VPWR net5811 sky130_fd_sc_hd__buf_1
Xwire6556 net6559 VGND VGND VPWR VPWR net6556 sky130_fd_sc_hd__buf_1
Xwire5822 net5823 VGND VGND VPWR VPWR net5822 sky130_fd_sc_hd__buf_1
X_21499_ _01381_ _01382_ _01380_ VGND VGND VPWR VPWR _01512_ sky130_fd_sc_hd__o21ba_1
Xwire5833 net5834 VGND VGND VPWR VPWR net5833 sky130_fd_sc_hd__clkbuf_1
Xwire6578 net6572 VGND VGND VPWR VPWR net6578 sky130_fd_sc_hd__buf_1
X_14040_ _06298_ _06303_ VGND VGND VPWR VPWR _06304_ sky130_fd_sc_hd__xor2_1
Xwire6589 net6586 VGND VGND VPWR VPWR net6589 sky130_fd_sc_hd__clkbuf_1
Xwire5844 net5845 VGND VGND VPWR VPWR net5844 sky130_fd_sc_hd__buf_1
X_23238_ net4984 net4967 _03065_ VGND VGND VPWR VPWR _03108_ sky130_fd_sc_hd__nand3_1
Xmax_length2287 net2288 VGND VGND VPWR VPWR net2287 sky130_fd_sc_hd__clkbuf_2
Xwire5855 pid_d.mult0.b\[5\] VGND VGND VPWR VPWR net5855 sky130_fd_sc_hd__clkbuf_1
Xwire5866 net5860 VGND VGND VPWR VPWR net5866 sky130_fd_sc_hd__clkbuf_1
Xwire5877 pid_d.mult0.b\[4\] VGND VGND VPWR VPWR net5877 sky130_fd_sc_hd__clkbuf_1
Xwire5899 net5900 VGND VGND VPWR VPWR net5899 sky130_fd_sc_hd__clkbuf_1
X_23169_ net5090 net4736 VGND VGND VPWR VPWR _03039_ sky130_fd_sc_hd__and2_1
X_15991_ _08052_ net1258 VGND VGND VPWR VPWR _08059_ sky130_fd_sc_hd__xnor2_1
X_17730_ net8052 net2596 VGND VGND VPWR VPWR _09588_ sky130_fd_sc_hd__nand2_1
X_14942_ _07015_ VGND VGND VPWR VPWR _07016_ sky130_fd_sc_hd__buf_1
X_17661_ _09539_ _09540_ VGND VGND VPWR VPWR _09541_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14873_ _06954_ VGND VGND VPWR VPWR _00207_ sky130_fd_sc_hd__clkbuf_1
X_19400_ _11235_ _11232_ _11236_ _11231_ VGND VGND VPWR VPWR _11237_ sky130_fd_sc_hd__o211a_1
X_16612_ matmul0.matmul_stage_inst.mult2\[13\] net181 net3468 VGND VGND VPWR VPWR
+ _08656_ sky130_fd_sc_hd__mux2_1
X_13824_ _06051_ _06089_ _06090_ VGND VGND VPWR VPWR _06091_ sky130_fd_sc_hd__o21a_1
X_17592_ svm0.tB\[14\] net6689 VGND VGND VPWR VPWR _09473_ sky130_fd_sc_hd__and2b_1
XFILLER_0_106_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19331_ _11156_ _11160_ _11167_ VGND VGND VPWR VPWR _11168_ sky130_fd_sc_hd__a21o_1
X_16543_ _08559_ _08560_ VGND VGND VPWR VPWR _08602_ sky130_fd_sc_hd__or2b_1
X_13755_ _05979_ net727 VGND VGND VPWR VPWR _06023_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12706_ net1008 _04978_ VGND VGND VPWR VPWR _04979_ sky130_fd_sc_hd__xnor2_4
X_19262_ _11034_ net3180 _11098_ VGND VGND VPWR VPWR _11099_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16474_ _08467_ _08472_ net1507 VGND VGND VPWR VPWR _08535_ sky130_fd_sc_hd__o21ba_1
X_13686_ _05879_ _05880_ _05886_ VGND VGND VPWR VPWR _05955_ sky130_fd_sc_hd__or3_1
XFILLER_0_127_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8353 net8360 VGND VGND VPWR VPWR net8353 sky130_fd_sc_hd__buf_1
X_18213_ net6886 net6810 VGND VGND VPWR VPWR _10064_ sky130_fd_sc_hd__nand2_1
X_15425_ net1543 net2703 net1877 VGND VGND VPWR VPWR _07499_ sky130_fd_sc_hd__o21a_1
Xfanout7641 net7648 VGND VGND VPWR VPWR net7641 sky130_fd_sc_hd__buf_1
X_12637_ net7337 net3030 net2988 VGND VGND VPWR VPWR _04910_ sky130_fd_sc_hd__nand3_1
X_19193_ net3183 _11028_ _11029_ VGND VGND VPWR VPWR _11030_ sky130_fd_sc_hd__a21o_1
XFILLER_0_171_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18144_ _09901_ _09993_ _09994_ VGND VGND VPWR VPWR _09995_ sky130_fd_sc_hd__o21ba_1
Xwire8470 net8468 VGND VGND VPWR VPWR net8470 sky130_fd_sc_hd__buf_1
X_12568_ net3031 VGND VGND VPWR VPWR _04858_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15356_ _07318_ _07429_ VGND VGND VPWR VPWR _07430_ sky130_fd_sc_hd__xnor2_1
Xwire8481 net8482 VGND VGND VPWR VPWR net8481 sky130_fd_sc_hd__clkbuf_1
Xmax_length4190 net4191 VGND VGND VPWR VPWR net4190 sky130_fd_sc_hd__buf_1
Xwire160 _06462_ VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_152_Right_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6973 net6979 VGND VGND VPWR VPWR net6973 sky130_fd_sc_hd__buf_1
X_14307_ matmul0.alpha_pass\[0\] net1302 net2898 net5367 _06528_ VGND VGND VPWR VPWR
+ _06529_ sky130_fd_sc_hd__a221o_1
Xwire7780 net7781 VGND VGND VPWR VPWR net7780 sky130_fd_sc_hd__clkbuf_1
X_18075_ _09924_ _09925_ VGND VGND VPWR VPWR _09926_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire171 net172 VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15287_ net2822 net2789 VGND VGND VPWR VPWR _07361_ sky130_fd_sc_hd__nor2_1
Xwire182 net183 VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_1
Xwire193 net194 VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_1
Xhold207 cordic0.slte0.opA\[1\] VGND VGND VPWR VPWR net9160 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 pid_d.mult0.b\[9\] VGND VGND VPWR VPWR net9171 sky130_fd_sc_hd__dlygate4sd3_1
X_17026_ net6478 net6473 _06503_ net6460 VGND VGND VPWR VPWR _08986_ sky130_fd_sc_hd__a31o_1
Xhold229 pid_d.prev_error\[1\] VGND VGND VPWR VPWR net9182 sky130_fd_sc_hd__dlygate4sd3_1
X_14238_ _06477_ _06490_ _06492_ _06493_ _06494_ VGND VGND VPWR VPWR _06495_ sky130_fd_sc_hd__a311o_1
XFILLER_0_180_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14169_ _06394_ _06423_ _06424_ _06395_ _06429_ VGND VGND VPWR VPWR _06430_ sky130_fd_sc_hd__o221a_1
XFILLER_0_1_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18977_ net6313 net6340 VGND VGND VPWR VPWR _10814_ sky130_fd_sc_hd__xnor2_1
X_17928_ _09773_ VGND VGND VPWR VPWR _09779_ sky130_fd_sc_hd__inv_2
X_17859_ net3971 net3258 _09709_ VGND VGND VPWR VPWR _09710_ sky130_fd_sc_hd__or3_1
XFILLER_0_191_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20870_ net5635 net5759 _00884_ _00885_ VGND VGND VPWR VPWR _00886_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_163_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19529_ _11302_ _11301_ _11363_ VGND VGND VPWR VPWR _11366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22540_ net9114 net1701 _02532_ VGND VGND VPWR VPWR _00542_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22471_ net5713 net5721 net5746 VGND VGND VPWR VPWR _02472_ sky130_fd_sc_hd__nand3_1
XFILLER_0_174_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24210_ _04069_ _04070_ VGND VGND VPWR VPWR _04071_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21422_ net9079 net3122 net2077 _01435_ VGND VGND VPWR VPWR _00521_ sky130_fd_sc_hd__a22o_1
X_25190_ clknet_leaf_57_clk _00079_ net8711 VGND VGND VPWR VPWR matmul0.a_in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24141_ _03976_ _04002_ VGND VGND VPWR VPWR _04003_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5107 net5110 VGND VGND VPWR VPWR net5107 sky130_fd_sc_hd__clkbuf_1
X_21353_ _01278_ _01279_ _01280_ VGND VGND VPWR VPWR _01367_ sky130_fd_sc_hd__o21a_1
Xwire5118 net5119 VGND VGND VPWR VPWR net5118 sky130_fd_sc_hd__clkbuf_1
Xwire5129 net5138 VGND VGND VPWR VPWR net5129 sky130_fd_sc_hd__buf_1
XFILLER_0_31_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20304_ net4040 net6478 VGND VGND VPWR VPWR _12109_ sky130_fd_sc_hd__nor2_1
X_24072_ _03920_ _03934_ VGND VGND VPWR VPWR _03935_ sky130_fd_sc_hd__xnor2_1
Xwire4406 pid_q.out\[12\] VGND VGND VPWR VPWR net4406 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4417 pid_q.out\[11\] VGND VGND VPWR VPWR net4417 sky130_fd_sc_hd__clkbuf_1
X_21284_ _01289_ _01298_ VGND VGND VPWR VPWR _01299_ sky130_fd_sc_hd__xor2_1
Xwire4428 net4429 VGND VGND VPWR VPWR net4428 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4439 net4440 VGND VGND VPWR VPWR net4439 sky130_fd_sc_hd__clkbuf_1
X_23023_ _02891_ _02892_ VGND VGND VPWR VPWR _02893_ sky130_fd_sc_hd__xnor2_1
Xwire3705 net3706 VGND VGND VPWR VPWR net3705 sky130_fd_sc_hd__clkbuf_2
X_20235_ _12052_ net6412 net2936 VGND VGND VPWR VPWR _12053_ sky130_fd_sc_hd__mux2_1
Xwire3727 net3728 VGND VGND VPWR VPWR net3727 sky130_fd_sc_hd__buf_1
Xwire3738 _03861_ VGND VGND VPWR VPWR net3738 sky130_fd_sc_hd__buf_1
Xwire3749 _03074_ VGND VGND VPWR VPWR net3749 sky130_fd_sc_hd__clkbuf_2
X_20166_ _11927_ _11991_ _11979_ net868 VGND VGND VPWR VPWR _11992_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_196_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24974_ pid_q.kp\[6\] _04714_ net1358 VGND VGND VPWR VPWR _04742_ sky130_fd_sc_hd__mux2_1
X_20097_ net9025 net2124 net1446 _11925_ VGND VGND VPWR VPWR _00461_ sky130_fd_sc_hd__a31o_1
X_23925_ net4661 net4830 VGND VGND VPWR VPWR _03789_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23856_ _03715_ _03720_ VGND VGND VPWR VPWR _03721_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22807_ _02711_ VGND VGND VPWR VPWR _00630_ sky130_fd_sc_hd__clkbuf_1
X_23787_ _03542_ _03557_ _03556_ VGND VGND VPWR VPWR _03653_ sky130_fd_sc_hd__a21oi_1
X_20999_ _00995_ _01004_ _01014_ VGND VGND VPWR VPWR _01015_ sky130_fd_sc_hd__a21o_1
Xmax_length7799 net7791 VGND VGND VPWR VPWR net7799 sky130_fd_sc_hd__clkbuf_1
X_25526_ clknet_leaf_35_clk _00406_ net8758 VGND VGND VPWR VPWR svm0.counter\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13540_ net7710 net2331 net2326 VGND VGND VPWR VPWR _05811_ sky130_fd_sc_hd__and3_1
XFILLER_0_137_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22738_ net3718 net107 VGND VGND VPWR VPWR _02670_ sky130_fd_sc_hd__and2_1
XFILLER_0_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13471_ net7685 net1151 VGND VGND VPWR VPWR _05744_ sky130_fd_sc_hd__nand2_1
X_22669_ _02619_ net5644 net2448 VGND VGND VPWR VPWR _02621_ sky130_fd_sc_hd__mux2_1
X_25457_ clknet_leaf_100_clk _00340_ net8389 VGND VGND VPWR VPWR cordic0.vec\[1\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire7010 net7011 VGND VGND VPWR VPWR net7010 sky130_fd_sc_hd__buf_1
XFILLER_0_30_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15210_ net3586 net3579 net3594 net3592 VGND VGND VPWR VPWR _07284_ sky130_fd_sc_hd__o22a_1
XFILLER_0_164_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24408_ net376 _04192_ _04193_ _04265_ _04196_ VGND VGND VPWR VPWR _04266_ sky130_fd_sc_hd__a311o_1
Xwire7032 net7030 VGND VGND VPWR VPWR net7032 sky130_fd_sc_hd__buf_2
X_16190_ net1251 net1508 VGND VGND VPWR VPWR _08255_ sky130_fd_sc_hd__xnor2_1
Xfanout6247 net6251 VGND VGND VPWR VPWR net6247 sky130_fd_sc_hd__buf_1
X_25388_ clknet_leaf_80_clk _00271_ net8498 VGND VGND VPWR VPWR matmul0.b\[7\] sky130_fd_sc_hd__dfrtp_1
Xwire7054 net7055 VGND VGND VPWR VPWR net7054 sky130_fd_sc_hd__clkbuf_1
Xfanout6258 net6283 VGND VGND VPWR VPWR net6258 sky130_fd_sc_hd__clkbuf_2
Xfanout6269 net6281 VGND VGND VPWR VPWR net6269 sky130_fd_sc_hd__buf_1
Xwire7065 net7062 VGND VGND VPWR VPWR net7065 sky130_fd_sc_hd__buf_1
Xwire6331 net6332 VGND VGND VPWR VPWR net6331 sky130_fd_sc_hd__clkbuf_1
X_15141_ _07202_ _07203_ _07214_ VGND VGND VPWR VPWR _07215_ sky130_fd_sc_hd__o21a_1
Xwire7076 net7077 VGND VGND VPWR VPWR net7076 sky130_fd_sc_hd__buf_1
XFILLER_0_51_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24339_ _04144_ _04150_ _04143_ VGND VGND VPWR VPWR _04198_ sky130_fd_sc_hd__o21ba_1
Xwire6342 net6341 VGND VGND VPWR VPWR net6342 sky130_fd_sc_hd__buf_1
Xwire7087 net7088 VGND VGND VPWR VPWR net7087 sky130_fd_sc_hd__clkbuf_1
Xwire6364 cordic0.vec\[0\]\[0\] VGND VGND VPWR VPWR net6364 sky130_fd_sc_hd__clkbuf_1
Xfanout5568 pid_d.mult0.a\[5\] VGND VGND VPWR VPWR net5568 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15072_ _07145_ VGND VGND VPWR VPWR _07146_ sky130_fd_sc_hd__buf_1
Xwire6386 net6387 VGND VGND VPWR VPWR net6386 sky130_fd_sc_hd__buf_1
Xwire5652 net5656 VGND VGND VPWR VPWR net5652 sky130_fd_sc_hd__clkbuf_1
Xwire6397 net6398 VGND VGND VPWR VPWR net6397 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length1350 net1351 VGND VGND VPWR VPWR net1350 sky130_fd_sc_hd__clkbuf_2
Xwire5663 net5664 VGND VGND VPWR VPWR net5663 sky130_fd_sc_hd__buf_1
X_14023_ _06285_ _06286_ VGND VGND VPWR VPWR _06287_ sky130_fd_sc_hd__and2_1
X_18900_ net3922 _10597_ _10735_ _10740_ VGND VGND VPWR VPWR _10741_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_31_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19880_ _11655_ _11659_ _11656_ VGND VGND VPWR VPWR _11713_ sky130_fd_sc_hd__a21bo_1
Xwire4951 net4952 VGND VGND VPWR VPWR net4951 sky130_fd_sc_hd__buf_1
Xwire5696 net5697 VGND VGND VPWR VPWR net5696 sky130_fd_sc_hd__clkbuf_1
Xwire4973 net4974 VGND VGND VPWR VPWR net4973 sky130_fd_sc_hd__buf_1
Xwire4984 net4985 VGND VGND VPWR VPWR net4984 sky130_fd_sc_hd__buf_1
X_18831_ net6837 net3920 _10638_ _10671_ _10673_ VGND VGND VPWR VPWR _10674_ sky130_fd_sc_hd__o311a_1
Xwire4995 net4988 VGND VGND VPWR VPWR net4995 sky130_fd_sc_hd__clkbuf_1
X_18762_ _10516_ _10564_ _10606_ net421 VGND VGND VPWR VPWR _10607_ sky130_fd_sc_hd__a2bb2o_1
X_15974_ _08039_ _08041_ VGND VGND VPWR VPWR _08042_ sky130_fd_sc_hd__xor2_1
X_17713_ net9239 net1217 net1451 pid_q.curr_int\[4\] VGND VGND VPWR VPWR _00418_ sky130_fd_sc_hd__a22o_1
X_14925_ net6627 matmul0.matmul_stage_inst.d\[7\] matmul0.matmul_stage_inst.c\[7\]
+ net6535 VGND VGND VPWR VPWR _06999_ sky130_fd_sc_hd__a22o_1
X_18693_ net6829 net6809 VGND VGND VPWR VPWR _10539_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold90 pid_d.curr_error\[11\] VGND VGND VPWR VPWR net9043 sky130_fd_sc_hd__dlygate4sd3_1
X_17644_ net6684 svm0.tA\[15\] VGND VGND VPWR VPWR _09524_ sky130_fd_sc_hd__xor2_1
X_14856_ _06945_ VGND VGND VPWR VPWR _00199_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_187_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_187_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13807_ _06024_ _06074_ VGND VGND VPWR VPWR _06075_ sky130_fd_sc_hd__xnor2_1
X_17575_ _09453_ _09456_ _09452_ VGND VGND VPWR VPWR _09457_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14787_ _06904_ _06908_ _06909_ net3627 VGND VGND VPWR VPWR _06910_ sky130_fd_sc_hd__a211o_1
X_19314_ _11146_ _11150_ VGND VGND VPWR VPWR _11151_ sky130_fd_sc_hd__xnor2_2
X_16526_ _08583_ _08585_ VGND VGND VPWR VPWR _08586_ sky130_fd_sc_hd__xnor2_1
X_13738_ _05872_ _06003_ _06006_ VGND VGND VPWR VPWR _06007_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_133_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19245_ net6240 _11056_ net3178 VGND VGND VPWR VPWR _11082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16457_ net2245 _08456_ _08517_ net2628 VGND VGND VPWR VPWR _08518_ sky130_fd_sc_hd__a211o_1
XFILLER_0_183_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13669_ net7746 net1306 VGND VGND VPWR VPWR _05938_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15408_ _07360_ _07481_ VGND VGND VPWR VPWR _07482_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_171_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19176_ _11012_ _10958_ _10959_ VGND VGND VPWR VPWR _11013_ sky130_fd_sc_hd__nand3_1
X_16388_ net3415 VGND VGND VPWR VPWR _08450_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18127_ _09800_ net3265 net3339 VGND VGND VPWR VPWR _09978_ sky130_fd_sc_hd__a21o_1
X_15339_ net1878 net1275 VGND VGND VPWR VPWR _07413_ sky130_fd_sc_hd__xor2_1
XFILLER_0_182_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6792 net6797 VGND VGND VPWR VPWR net6792 sky130_fd_sc_hd__dlymetal6s2s_1
X_18058_ net6989 net7096 VGND VGND VPWR VPWR _09909_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17009_ net6500 net3335 VGND VGND VPWR VPWR _08970_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20020_ net1406 net2093 _11849_ VGND VGND VPWR VPWR _11850_ sky130_fd_sc_hd__a21oi_2
X_21971_ _01974_ _01977_ _01978_ VGND VGND VPWR VPWR _01979_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_174_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23710_ pid_q.curr_int\[3\] net3062 net2029 _03576_ VGND VGND VPWR VPWR _00668_ sky130_fd_sc_hd__a22o_1
X_20922_ _00936_ _00937_ VGND VGND VPWR VPWR _00938_ sky130_fd_sc_hd__xnor2_2
X_24690_ net3715 _04527_ VGND VGND VPWR VPWR _04528_ sky130_fd_sc_hd__or2_1
Xmax_length7029 net7027 VGND VGND VPWR VPWR net7029 sky130_fd_sc_hd__buf_1
XFILLER_0_178_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23641_ net1666 _03507_ VGND VGND VPWR VPWR _03508_ sky130_fd_sc_hd__xnor2_1
X_20853_ net5473 _00868_ VGND VGND VPWR VPWR _00869_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23572_ net2420 _03361_ _03354_ VGND VGND VPWR VPWR _03440_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20784_ _12542_ _12553_ _12554_ VGND VGND VPWR VPWR _12555_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4915 net4911 VGND VGND VPWR VPWR net4915 sky130_fd_sc_hd__buf_1
X_22523_ net4325 net3101 net8887 VGND VGND VPWR VPWR _02523_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25311_ clknet_leaf_79_clk _00194_ net8490 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.e\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire907 net908 VGND VGND VPWR VPWR net907 sky130_fd_sc_hd__buf_1
XFILLER_0_29_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length4959 net4960 VGND VGND VPWR VPWR net4959 sky130_fd_sc_hd__clkbuf_2
Xwire918 _05409_ VGND VGND VPWR VPWR net918 sky130_fd_sc_hd__buf_1
XFILLER_0_88_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire929 _04242_ VGND VGND VPWR VPWR net929 sky130_fd_sc_hd__buf_1
X_22454_ _02455_ VGND VGND VPWR VPWR _02456_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25242_ clknet_leaf_86_clk _00125_ net8531 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.a\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_161_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21405_ net860 _01418_ VGND VGND VPWR VPWR _01419_ sky130_fd_sc_hd__xnor2_1
X_25173_ clknet_leaf_54_clk _00062_ net8730 VGND VGND VPWR VPWR svm0.periodTop\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22385_ net551 net549 VGND VGND VPWR VPWR _02388_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24124_ net4579 net4866 VGND VGND VPWR VPWR _03986_ sky130_fd_sc_hd__nand2_1
X_21336_ net5654 _01349_ VGND VGND VPWR VPWR _01350_ sky130_fd_sc_hd__xor2_1
XFILLER_0_20_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4203 net4204 VGND VGND VPWR VPWR net4203 sky130_fd_sc_hd__buf_1
XFILLER_0_4_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4214 net4215 VGND VGND VPWR VPWR net4214 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4225 _06708_ VGND VGND VPWR VPWR net4225 sky130_fd_sc_hd__clkbuf_1
X_24055_ _03909_ _03917_ VGND VGND VPWR VPWR _03918_ sky130_fd_sc_hd__xnor2_2
Xwire4236 _06512_ VGND VGND VPWR VPWR net4236 sky130_fd_sc_hd__clkbuf_1
Xwire3502 net3503 VGND VGND VPWR VPWR net3502 sky130_fd_sc_hd__buf_1
X_21267_ _01278_ _01281_ VGND VGND VPWR VPWR _01282_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire4269 net4270 VGND VGND VPWR VPWR net4269 sky130_fd_sc_hd__clkbuf_1
Xwire3524 net3525 VGND VGND VPWR VPWR net3524 sky130_fd_sc_hd__clkbuf_1
X_23006_ net5086 net4613 VGND VGND VPWR VPWR _02876_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire3535 net3536 VGND VGND VPWR VPWR net3535 sky130_fd_sc_hd__buf_1
XFILLER_0_21_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20218_ _12039_ VGND VGND VPWR VPWR _00468_ sky130_fd_sc_hd__clkbuf_1
Xwire2801 _07125_ VGND VGND VPWR VPWR net2801 sky130_fd_sc_hd__buf_1
Xwire3546 net3547 VGND VGND VPWR VPWR net3546 sky130_fd_sc_hd__buf_1
X_21198_ _01144_ _01147_ _01206_ _01207_ VGND VGND VPWR VPWR _01214_ sky130_fd_sc_hd__a22o_1
Xwire3557 net3558 VGND VGND VPWR VPWR net3557 sky130_fd_sc_hd__buf_1
Xwire2823 net2826 VGND VGND VPWR VPWR net2823 sky130_fd_sc_hd__clkbuf_1
Xwire3568 _07034_ VGND VGND VPWR VPWR net3568 sky130_fd_sc_hd__buf_1
Xwire2834 net2835 VGND VGND VPWR VPWR net2834 sky130_fd_sc_hd__buf_1
Xwire3579 _07021_ VGND VGND VPWR VPWR net3579 sky130_fd_sc_hd__buf_1
XFILLER_0_21_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20149_ _11974_ _11975_ VGND VGND VPWR VPWR _11976_ sky130_fd_sc_hd__xor2_1
Xwire2867 net2868 VGND VGND VPWR VPWR net2867 sky130_fd_sc_hd__buf_1
Xwire2889 net2890 VGND VGND VPWR VPWR net2889 sky130_fd_sc_hd__buf_1
X_24957_ net8869 net136 VGND VGND VPWR VPWR _04732_ sky130_fd_sc_hd__and2b_1
X_12971_ net850 _05199_ _05168_ _05169_ VGND VGND VPWR VPWR _05244_ sky130_fd_sc_hd__and4_1
XFILLER_0_99_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14710_ net9082 net2861 net2263 net1290 VGND VGND VPWR VPWR _00146_ sky130_fd_sc_hd__a22o_1
X_23908_ _03770_ _03673_ _03771_ VGND VGND VPWR VPWR _03772_ sky130_fd_sc_hd__o21a_1
X_15690_ net3517 VGND VGND VPWR VPWR _07761_ sky130_fd_sc_hd__buf_1
X_24888_ _04683_ VGND VGND VPWR VPWR _00739_ sky130_fd_sc_hd__clkbuf_1
Xmax_length7530 net7531 VGND VGND VPWR VPWR net7530 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14641_ net8979 net2879 _06804_ VGND VGND VPWR VPWR _00125_ sky130_fd_sc_hd__a21o_1
X_23839_ net2412 _03703_ net5155 VGND VGND VPWR VPWR _03704_ sky130_fd_sc_hd__o21ba_1
Xmax_length7563 matmul0.b_in\[11\] VGND VGND VPWR VPWR net7563 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17360_ net6657 net3389 _09269_ VGND VGND VPWR VPWR _09273_ sky130_fd_sc_hd__o21ba_1
X_14572_ _06746_ _06748_ _06741_ VGND VGND VPWR VPWR _06749_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16311_ net424 _08302_ VGND VGND VPWR VPWR _08374_ sky130_fd_sc_hd__nand2_1
Xmax_length6884 net6885 VGND VGND VPWR VPWR net6884 sky130_fd_sc_hd__clkbuf_1
X_13523_ net7805 net2950 net3669 VGND VGND VPWR VPWR _05794_ sky130_fd_sc_hd__and3_1
X_25509_ clknet_leaf_36_clk _00389_ net8754 VGND VGND VPWR VPWR svm0.delta\[14\] sky130_fd_sc_hd__dfrtp_2
X_17291_ net6687 VGND VGND VPWR VPWR _09205_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19030_ _10795_ _10864_ _10817_ _10866_ VGND VGND VPWR VPWR _10867_ sky130_fd_sc_hd__a31o_1
XFILLER_0_83_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout6011 net6017 VGND VGND VPWR VPWR net6011 sky130_fd_sc_hd__buf_1
X_16242_ _08306_ VGND VGND VPWR VPWR _00224_ sky130_fd_sc_hd__clkbuf_1
X_13454_ _05699_ _05725_ _05726_ VGND VGND VPWR VPWR _05727_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6044 net6047 VGND VGND VPWR VPWR net6044 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13385_ _05553_ _05561_ VGND VGND VPWR VPWR _05658_ sky130_fd_sc_hd__xnor2_1
X_16173_ net493 net492 VGND VGND VPWR VPWR _08238_ sky130_fd_sc_hd__nand2_1
Xfanout6077 net6083 VGND VGND VPWR VPWR net6077 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout6088 net6090 VGND VGND VPWR VPWR net6088 sky130_fd_sc_hd__clkbuf_2
Xwire6150 net6146 VGND VGND VPWR VPWR net6150 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6161 net6159 VGND VGND VPWR VPWR net6161 sky130_fd_sc_hd__clkbuf_1
X_15124_ _07172_ _07173_ VGND VGND VPWR VPWR _07198_ sky130_fd_sc_hd__xnor2_1
Xwire6172 net6173 VGND VGND VPWR VPWR net6172 sky130_fd_sc_hd__buf_1
XFILLER_0_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5398 pid_d.mult0.a\[14\] VGND VGND VPWR VPWR net5398 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_10_Left_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19932_ net6007 net2498 VGND VGND VPWR VPWR _11764_ sky130_fd_sc_hd__nand2_1
X_15055_ _07128_ VGND VGND VPWR VPWR _07129_ sky130_fd_sc_hd__buf_1
Xwire5482 net5483 VGND VGND VPWR VPWR net5482 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5493 net5494 VGND VGND VPWR VPWR net5493 sky130_fd_sc_hd__clkbuf_1
X_14006_ svm0.tC\[7\] net1126 net189 net1926 VGND VGND VPWR VPWR _00024_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4770 net4761 VGND VGND VPWR VPWR net4770 sky130_fd_sc_hd__clkbuf_1
X_19863_ net2095 _11695_ VGND VGND VPWR VPWR _11696_ sky130_fd_sc_hd__xnor2_1
Xwire4781 net4782 VGND VGND VPWR VPWR net4781 sky130_fd_sc_hd__clkbuf_1
Xwire4792 net4793 VGND VGND VPWR VPWR net4792 sky130_fd_sc_hd__buf_1
XFILLER_0_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18814_ net6376 _10656_ _10623_ VGND VGND VPWR VPWR _10658_ sky130_fd_sc_hd__and3_1
X_19794_ net6008 net2100 net3138 VGND VGND VPWR VPWR _11628_ sky130_fd_sc_hd__a21oi_1
X_18745_ net6781 net2125 VGND VGND VPWR VPWR _10590_ sky130_fd_sc_hd__or2_1
X_15957_ _07963_ _07964_ _08024_ VGND VGND VPWR VPWR _08025_ sky130_fd_sc_hd__a21o_1
XFILLER_0_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14908_ net6636 matmul0.matmul_stage_inst.d\[8\] net7410 net6531 VGND VGND VPWR VPWR
+ _06982_ sky130_fd_sc_hd__a22o_1
X_18676_ _10103_ VGND VGND VPWR VPWR _10522_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15888_ net1525 net1523 VGND VGND VPWR VPWR _07957_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_188_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17627_ svm0.tB\[7\] _09477_ _09507_ VGND VGND VPWR VPWR _09508_ sky130_fd_sc_hd__o21a_1
X_14839_ _06936_ VGND VGND VPWR VPWR _00191_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17558_ net3278 svm0.tC\[10\] VGND VGND VPWR VPWR _09440_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16509_ net880 net879 VGND VGND VPWR VPWR _08569_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17489_ svm0.delta\[8\] net770 VGND VGND VPWR VPWR _09379_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19228_ net6139 _11062_ _11063_ _11064_ net3918 VGND VGND VPWR VPWR _11065_ sky130_fd_sc_hd__a311o_1
XFILLER_0_160_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19159_ net6049 VGND VGND VPWR VPWR _10996_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22170_ _02174_ _02102_ _02175_ VGND VGND VPWR VPWR _02176_ sky130_fd_sc_hd__a21o_1
XFILLER_0_83_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21121_ net5584 _01119_ _01117_ VGND VGND VPWR VPWR _01137_ sky130_fd_sc_hd__or3_1
XFILLER_0_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21052_ _01033_ _01034_ _01067_ VGND VGND VPWR VPWR _01068_ sky130_fd_sc_hd__a21o_1
Xwire2108 _11145_ VGND VGND VPWR VPWR net2108 sky130_fd_sc_hd__buf_1
Xwire2119 net2120 VGND VGND VPWR VPWR net2119 sky130_fd_sc_hd__clkbuf_1
X_20003_ _10344_ _11833_ VGND VGND VPWR VPWR _11834_ sky130_fd_sc_hd__nor2_1
X_25860_ clknet_leaf_16_clk _00733_ net8619 VGND VGND VPWR VPWR pid_q.mult0.a\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1407 _11796_ VGND VGND VPWR VPWR net1407 sky130_fd_sc_hd__clkbuf_1
Xwire1418 _11390_ VGND VGND VPWR VPWR net1418 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1429 _10586_ VGND VGND VPWR VPWR net1429 sky130_fd_sc_hd__dlymetal6s2s_1
X_24811_ net5189 _04633_ net5194 VGND VGND VPWR VPWR _04634_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25791_ clknet_leaf_60_clk _00664_ net8669 VGND VGND VPWR VPWR svm0.in_valid sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24742_ net5259 _04573_ VGND VGND VPWR VPWR _04574_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_193_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21954_ net5858 net3787 net5841 VGND VGND VPWR VPWR _01962_ sky130_fd_sc_hd__o21a_1
XFILLER_0_179_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20905_ _00918_ _00920_ VGND VGND VPWR VPWR _00921_ sky130_fd_sc_hd__and2_1
X_24673_ pid_q.curr_error\[8\] _00011_ net1374 VGND VGND VPWR VPWR _04519_ sky130_fd_sc_hd__and3_1
X_21885_ net2477 VGND VGND VPWR VPWR _01894_ sky130_fd_sc_hd__buf_1
Xmax_length6114 net6115 VGND VGND VPWR VPWR net6114 sky130_fd_sc_hd__buf_1
XFILLER_0_90_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23624_ net4664 net4899 VGND VGND VPWR VPWR _03491_ sky130_fd_sc_hd__nand2_1
X_20836_ net5741 net5597 VGND VGND VPWR VPWR _00852_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23555_ net1384 _03422_ VGND VGND VPWR VPWR _03423_ sky130_fd_sc_hd__xnor2_2
X_20767_ net5596 net5794 VGND VGND VPWR VPWR _12538_ sky130_fd_sc_hd__nand2_1
XFILLER_0_193_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire704 _01252_ VGND VGND VPWR VPWR net704 sky130_fd_sc_hd__clkbuf_1
X_22506_ _02505_ _02506_ _02417_ VGND VGND VPWR VPWR _02507_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23486_ _03241_ _03242_ _03243_ VGND VGND VPWR VPWR _03355_ sky130_fd_sc_hd__o21ai_1
Xwire715 _10152_ VGND VGND VPWR VPWR net715 sky130_fd_sc_hd__buf_1
Xwire726 _06702_ VGND VGND VPWR VPWR net726 sky130_fd_sc_hd__buf_1
X_20698_ _12466_ _12467_ _12471_ VGND VGND VPWR VPWR _12472_ sky130_fd_sc_hd__o21a_1
Xwire737 _04585_ VGND VGND VPWR VPWR net737 sky130_fd_sc_hd__buf_1
Xwire748 _03381_ VGND VGND VPWR VPWR net748 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22437_ _02358_ _02365_ _02364_ VGND VGND VPWR VPWR _02439_ sky130_fd_sc_hd__a21o_1
X_25225_ clknet_leaf_59_clk _00114_ net8694 VGND VGND VPWR VPWR svm0.vC\[13\] sky130_fd_sc_hd__dfrtp_1
Xwire759 _01250_ VGND VGND VPWR VPWR net759 sky130_fd_sc_hd__buf_1
XFILLER_0_162_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13170_ net7778 net2334 net2974 VGND VGND VPWR VPWR _05443_ sky130_fd_sc_hd__and3_1
X_25156_ clknet_leaf_44_clk _00045_ net8781 VGND VGND VPWR VPWR pid_q.target\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_22368_ _02345_ _02370_ VGND VGND VPWR VPWR _02371_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4000 _09581_ VGND VGND VPWR VPWR net4000 sky130_fd_sc_hd__buf_1
Xwire4022 net4023 VGND VGND VPWR VPWR net4022 sky130_fd_sc_hd__buf_1
X_24107_ net5059 net5028 net5075 VGND VGND VPWR VPWR _03969_ sky130_fd_sc_hd__o21ai_1
X_21319_ pid_d.prev_error\[0\] net5973 _01332_ VGND VGND VPWR VPWR _01334_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4033 net4034 VGND VGND VPWR VPWR net4033 sky130_fd_sc_hd__buf_1
X_25087_ net5172 _04831_ VGND VGND VPWR VPWR _04832_ sky130_fd_sc_hd__xnor2_1
X_22299_ net1702 _02302_ VGND VGND VPWR VPWR _02303_ sky130_fd_sc_hd__xor2_1
Xwire4044 _08966_ VGND VGND VPWR VPWR net4044 sky130_fd_sc_hd__buf_1
Xwire4055 _08896_ VGND VGND VPWR VPWR net4055 sky130_fd_sc_hd__buf_1
Xwire3310 net3311 VGND VGND VPWR VPWR net3310 sky130_fd_sc_hd__buf_1
X_24038_ net4606 net4851 VGND VGND VPWR VPWR _03901_ sky130_fd_sc_hd__nand2_1
Xwire3321 net3322 VGND VGND VPWR VPWR net3321 sky130_fd_sc_hd__clkbuf_1
Xwire4066 _08659_ VGND VGND VPWR VPWR net4066 sky130_fd_sc_hd__clkbuf_1
Xwire3332 _08971_ VGND VGND VPWR VPWR net3332 sky130_fd_sc_hd__buf_1
Xwire4077 net4078 VGND VGND VPWR VPWR net4077 sky130_fd_sc_hd__buf_1
Xwire4088 _07483_ VGND VGND VPWR VPWR net4088 sky130_fd_sc_hd__clkbuf_1
Xwire4099 net4100 VGND VGND VPWR VPWR net4099 sky130_fd_sc_hd__buf_1
X_16860_ net6471 VGND VGND VPWR VPWR _08825_ sky130_fd_sc_hd__inv_2
Xwire2631 net2632 VGND VGND VPWR VPWR net2631 sky130_fd_sc_hd__clkbuf_2
Xwire3376 _08781_ VGND VGND VPWR VPWR net3376 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2642 net2644 VGND VGND VPWR VPWR net2642 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3398 _07654_ VGND VGND VPWR VPWR net3398 sky130_fd_sc_hd__clkbuf_2
Xwire2653 _07759_ VGND VGND VPWR VPWR net2653 sky130_fd_sc_hd__clkbuf_1
Xwire2664 net2665 VGND VGND VPWR VPWR net2664 sky130_fd_sc_hd__buf_1
Xwire1930 net1931 VGND VGND VPWR VPWR net1930 sky130_fd_sc_hd__buf_1
X_15811_ _07785_ _07790_ VGND VGND VPWR VPWR _07881_ sky130_fd_sc_hd__nand2_1
Xwire2675 _07681_ VGND VGND VPWR VPWR net2675 sky130_fd_sc_hd__buf_1
Xwire1941 _05617_ VGND VGND VPWR VPWR net1941 sky130_fd_sc_hd__buf_1
Xwire2686 _07534_ VGND VGND VPWR VPWR net2686 sky130_fd_sc_hd__buf_1
X_16791_ _08785_ VGND VGND VPWR VPWR _00294_ sky130_fd_sc_hd__clkbuf_1
Xwire1952 net1953 VGND VGND VPWR VPWR net1952 sky130_fd_sc_hd__buf_1
Xwire2697 net2698 VGND VGND VPWR VPWR net2697 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1963 net1964 VGND VGND VPWR VPWR net1963 sky130_fd_sc_hd__buf_1
Xwire1974 _04924_ VGND VGND VPWR VPWR net1974 sky130_fd_sc_hd__buf_1
X_18530_ _10377_ _10378_ VGND VGND VPWR VPWR _10379_ sky130_fd_sc_hd__and2b_1
X_15742_ net2758 net1265 _07812_ VGND VGND VPWR VPWR _07813_ sky130_fd_sc_hd__o21ai_1
X_12954_ _05002_ _05226_ VGND VGND VPWR VPWR _05227_ sky130_fd_sc_hd__nand2_1
Xwire1996 net1997 VGND VGND VPWR VPWR net1996 sky130_fd_sc_hd__buf_2
XFILLER_0_88_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18461_ net3925 net3225 VGND VGND VPWR VPWR _10311_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15673_ _07691_ _07742_ _07743_ VGND VGND VPWR VPWR _07744_ sky130_fd_sc_hd__o21ai_1
X_12885_ _05156_ _05157_ VGND VGND VPWR VPWR _05158_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17412_ svm0.delta\[11\] VGND VGND VPWR VPWR _09315_ sky130_fd_sc_hd__inv_2
XFILLER_0_169_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14624_ _06512_ _06792_ _06793_ net9102 VGND VGND VPWR VPWR _00119_ sky130_fd_sc_hd__a22o_1
X_18392_ _10240_ _10242_ VGND VGND VPWR VPWR _10243_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length7382 matmul0.matmul_stage_inst.f\[11\] VGND VGND VPWR VPWR net7382 sky130_fd_sc_hd__buf_1
XFILLER_0_184_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17343_ svm0.counter\[10\] VGND VGND VPWR VPWR _09257_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14555_ _06731_ _06732_ VGND VGND VPWR VPWR _06733_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13506_ _05776_ _00411_ VGND VGND VPWR VPWR _05778_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17274_ net2982 net174 net2157 net9172 VGND VGND VPWR VPWR _00368_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14486_ _06667_ _06670_ VGND VGND VPWR VPWR _06671_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19013_ net6226 net6205 VGND VGND VPWR VPWR _10850_ sky130_fd_sc_hd__nor2b_2
X_16225_ net1254 VGND VGND VPWR VPWR _08290_ sky130_fd_sc_hd__buf_1
X_13437_ net7832 net2950 net3669 VGND VGND VPWR VPWR _05710_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16156_ _08214_ _08221_ VGND VGND VPWR VPWR _08222_ sky130_fd_sc_hd__xnor2_2
X_13368_ net5189 net2963 net2986 net7199 VGND VGND VPWR VPWR _05641_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15107_ _07177_ _07178_ _07180_ VGND VGND VPWR VPWR _07181_ sky130_fd_sc_hd__a21o_1
X_16087_ _08068_ net1257 net1521 VGND VGND VPWR VPWR _08154_ sky130_fd_sc_hd__a21o_1
X_13299_ _05501_ _05515_ net847 VGND VGND VPWR VPWR _05572_ sky130_fd_sc_hd__a21o_1
Xwire5290 net5291 VGND VGND VPWR VPWR net5290 sky130_fd_sc_hd__buf_1
X_19915_ _11745_ _11746_ _11690_ VGND VGND VPWR VPWR _11747_ sky130_fd_sc_hd__mux2_1
X_15038_ _06964_ net3521 VGND VGND VPWR VPWR _07112_ sky130_fd_sc_hd__nor2_1
X_19846_ net6128 _11445_ net6157 VGND VGND VPWR VPWR _11679_ sky130_fd_sc_hd__or3b_1
XFILLER_0_155_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16989_ net5989 _08944_ net2605 _08924_ VGND VGND VPWR VPWR _08951_ sky130_fd_sc_hd__a22o_1
X_19777_ cordic0.cos\[2\] net2942 net1782 VGND VGND VPWR VPWR _11612_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18728_ net6877 _10534_ VGND VGND VPWR VPWR _10573_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18659_ net714 _10505_ _10503_ VGND VGND VPWR VPWR _10506_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21670_ _01571_ _01573_ VGND VGND VPWR VPWR _01681_ sky130_fd_sc_hd__nand2_1
XFILLER_0_171_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20621_ _12400_ _12401_ VGND VGND VPWR VPWR _12402_ sky130_fd_sc_hd__and2b_1
XFILLER_0_188_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23340_ net5077 net4599 VGND VGND VPWR VPWR _03210_ sky130_fd_sc_hd__nand2_1
Xwire7609 net7610 VGND VGND VPWR VPWR net7609 sky130_fd_sc_hd__buf_1
X_20552_ _12333_ _12336_ VGND VGND VPWR VPWR _12337_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire6908 net6910 VGND VGND VPWR VPWR net6908 sky130_fd_sc_hd__buf_2
X_23271_ _03137_ _03135_ VGND VGND VPWR VPWR _03141_ sky130_fd_sc_hd__nor2_1
X_20483_ net2192 net2087 VGND VGND VPWR VPWR _12272_ sky130_fd_sc_hd__or2_1
X_22222_ net5800 net3786 _02226_ VGND VGND VPWR VPWR _02227_ sky130_fd_sc_hd__a21o_1
X_25010_ net7472 _04764_ _04765_ net7498 net512 VGND VGND VPWR VPWR _04766_ sky130_fd_sc_hd__a32o_1
XFILLER_0_70_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22153_ net1041 _02068_ _02067_ VGND VGND VPWR VPWR _02159_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21104_ _01117_ _01118_ _01119_ VGND VGND VPWR VPWR _01120_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22084_ _02084_ _02087_ VGND VGND VPWR VPWR _02091_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25912_ clknet_leaf_66_clk _00785_ net8659 VGND VGND VPWR VPWR pid_q.out\[8\] sky130_fd_sc_hd__dfrtp_1
X_21035_ net5641 net5775 net3836 _01049_ VGND VGND VPWR VPWR _01051_ sky130_fd_sc_hd__a211o_1
XFILLER_0_195_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1215 _09700_ VGND VGND VPWR VPWR net1215 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1226 _08991_ VGND VGND VPWR VPWR net1226 sky130_fd_sc_hd__buf_1
X_25843_ clknet_leaf_20_clk _00716_ net8747 VGND VGND VPWR VPWR pid_q.mult0.b\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1237 net1238 VGND VGND VPWR VPWR net1237 sky130_fd_sc_hd__buf_1
Xwire1248 _08391_ VGND VGND VPWR VPWR net1248 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1259 net1260 VGND VGND VPWR VPWR net1259 sky130_fd_sc_hd__clkbuf_1
X_25774_ clknet_leaf_26_clk _00647_ net8650 VGND VGND VPWR VPWR pid_d.out\[15\] sky130_fd_sc_hd__dfrtp_1
X_22986_ matmul0.beta_pass\[12\] net353 net6578 VGND VGND VPWR VPWR _02861_ sky130_fd_sc_hd__mux2_1
X_24725_ net5273 _04556_ _04557_ VGND VGND VPWR VPWR _04559_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21937_ _01943_ _01944_ VGND VGND VPWR VPWR _01945_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_195_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24656_ net1645 VGND VGND VPWR VPWR _04510_ sky130_fd_sc_hd__buf_1
X_12670_ net7813 net2338 net1968 VGND VGND VPWR VPWR _04943_ sky130_fd_sc_hd__and3_1
XFILLER_0_166_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21868_ net1171 _01876_ VGND VGND VPWR VPWR _01877_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8727 net8733 VGND VGND VPWR VPWR net8727 sky130_fd_sc_hd__buf_1
Xwire8800 net8801 VGND VGND VPWR VPWR net8800 sky130_fd_sc_hd__buf_1
X_23607_ pid_q.prev_error\[1\] net5168 VGND VGND VPWR VPWR _03475_ sky130_fd_sc_hd__nand2_1
Xwire8811 net8808 VGND VGND VPWR VPWR net8811 sky130_fd_sc_hd__buf_1
XFILLER_0_65_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20819_ _12555_ _12557_ _12552_ VGND VGND VPWR VPWR _00835_ sky130_fd_sc_hd__o21ba_1
Xwire8822 net8823 VGND VGND VPWR VPWR net8822 sky130_fd_sc_hd__buf_1
X_24587_ _04368_ _04370_ _04442_ VGND VGND VPWR VPWR _04443_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21799_ _01807_ _01808_ VGND VGND VPWR VPWR _01809_ sky130_fd_sc_hd__xnor2_1
Xwire8833 net8834 VGND VGND VPWR VPWR net8833 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4520 net4521 VGND VGND VPWR VPWR net4520 sky130_fd_sc_hd__clkbuf_1
Xwire8844 net8845 VGND VGND VPWR VPWR net8844 sky130_fd_sc_hd__clkbuf_1
X_14340_ net8233 net3643 VGND VGND VPWR VPWR _06557_ sky130_fd_sc_hd__and2_1
X_23538_ _03399_ _03404_ VGND VGND VPWR VPWR _03406_ sky130_fd_sc_hd__nand2_1
Xwire501 net502 VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire512 net513 VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8877 net8878 VGND VGND VPWR VPWR net8877 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire523 net524 VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4586 net4577 VGND VGND VPWR VPWR net4586 sky130_fd_sc_hd__clkbuf_1
Xwire534 _05762_ VGND VGND VPWR VPWR net534 sky130_fd_sc_hd__clkbuf_2
X_14271_ net64 _06511_ _06515_ net8999 VGND VGND VPWR VPWR _00044_ sky130_fd_sc_hd__a22o_1
Xwire545 net546 VGND VGND VPWR VPWR net545 sky130_fd_sc_hd__buf_1
X_23469_ net4641 net4962 VGND VGND VPWR VPWR _03338_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire556 net557 VGND VGND VPWR VPWR net556 sky130_fd_sc_hd__clkbuf_1
Xwire567 _11666_ VGND VGND VPWR VPWR net567 sky130_fd_sc_hd__buf_1
Xwire578 net579 VGND VGND VPWR VPWR net578 sky130_fd_sc_hd__buf_1
XFILLER_0_107_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16010_ _08001_ _07999_ VGND VGND VPWR VPWR _08078_ sky130_fd_sc_hd__or2b_1
X_13222_ net7650 net1972 net1969 VGND VGND VPWR VPWR _05495_ sky130_fd_sc_hd__and3_1
X_25208_ clknet_leaf_61_clk _00097_ net8671 VGND VGND VPWR VPWR matmul0.b_in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire589 _04104_ VGND VGND VPWR VPWR net589 sky130_fd_sc_hd__buf_1
XFILLER_0_27_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25139_ clknet_leaf_51_clk _00028_ net8810 VGND VGND VPWR VPWR svm0.tC\[11\] sky130_fd_sc_hd__dfrtp_1
X_13153_ _05416_ _05424_ _05425_ VGND VGND VPWR VPWR _05426_ sky130_fd_sc_hd__nand3_1
XFILLER_0_0_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13084_ _05294_ net1949 _05288_ net3688 VGND VGND VPWR VPWR _05357_ sky130_fd_sc_hd__and4_1
X_17961_ _09809_ _09811_ VGND VGND VPWR VPWR _09812_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3140 _11410_ VGND VGND VPWR VPWR net3140 sky130_fd_sc_hd__buf_1
XFILLER_0_97_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16912_ net6402 net6372 VGND VGND VPWR VPWR _08876_ sky130_fd_sc_hd__xor2_1
Xwire3151 _11382_ VGND VGND VPWR VPWR net3151 sky130_fd_sc_hd__buf_1
X_19700_ _11439_ _11535_ VGND VGND VPWR VPWR _11536_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3162 _11269_ VGND VGND VPWR VPWR net3162 sky130_fd_sc_hd__clkbuf_2
Xwire3173 _11122_ VGND VGND VPWR VPWR net3173 sky130_fd_sc_hd__buf_1
X_17892_ _09690_ _09635_ VGND VGND VPWR VPWR _09743_ sky130_fd_sc_hd__xnor2_1
Xwire3184 _10990_ VGND VGND VPWR VPWR net3184 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire2450 net2454 VGND VGND VPWR VPWR net2450 sky130_fd_sc_hd__clkbuf_1
Xwire3195 net3197 VGND VGND VPWR VPWR net3195 sky130_fd_sc_hd__buf_1
X_19631_ net3162 _11467_ VGND VGND VPWR VPWR _11468_ sky130_fd_sc_hd__xnor2_1
X_16843_ _08812_ VGND VGND VPWR VPWR _00319_ sky130_fd_sc_hd__clkbuf_1
Xwire2472 _02299_ VGND VGND VPWR VPWR net2472 sky130_fd_sc_hd__buf_1
Xwire2483 _00846_ VGND VGND VPWR VPWR net2483 sky130_fd_sc_hd__buf_1
Xwire2494 net2495 VGND VGND VPWR VPWR net2494 sky130_fd_sc_hd__buf_1
XFILLER_0_189_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19562_ _11324_ _11391_ _11395_ net6346 _11398_ VGND VGND VPWR VPWR _11399_ sky130_fd_sc_hd__a221o_1
Xwire1760 net1761 VGND VGND VPWR VPWR net1760 sky130_fd_sc_hd__buf_1
Xwire1771 net1772 VGND VGND VPWR VPWR net1771 sky130_fd_sc_hd__dlymetal6s2s_1
X_16774_ _08776_ VGND VGND VPWR VPWR _00286_ sky130_fd_sc_hd__clkbuf_1
X_13986_ _06201_ _06198_ _06250_ VGND VGND VPWR VPWR _06251_ sky130_fd_sc_hd__o21ai_1
Xwire1782 net1783 VGND VGND VPWR VPWR net1782 sky130_fd_sc_hd__clkbuf_1
Xwire1793 _09482_ VGND VGND VPWR VPWR net1793 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_189_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18513_ net3308 _10358_ _10361_ VGND VGND VPWR VPWR _10362_ sky130_fd_sc_hd__a21oi_1
X_15725_ net1851 net1537 _07795_ VGND VGND VPWR VPWR _07796_ sky130_fd_sc_hd__a21o_1
X_12937_ _05204_ _05209_ VGND VGND VPWR VPWR _05210_ sky130_fd_sc_hd__xor2_1
X_19493_ net6097 _11329_ VGND VGND VPWR VPWR _11330_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18444_ _10041_ _10292_ _10293_ VGND VGND VPWR VPWR _10294_ sky130_fd_sc_hd__o21a_1
X_15656_ _07584_ _07588_ net1272 VGND VGND VPWR VPWR _07728_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_34_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12868_ net1333 _05140_ VGND VGND VPWR VPWR _05141_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14607_ _06770_ _06771_ _06777_ VGND VGND VPWR VPWR _06780_ sky130_fd_sc_hd__mux2_1
X_18375_ net7015 net7046 VGND VGND VPWR VPWR _10226_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15587_ net1852 _07658_ VGND VGND VPWR VPWR _07659_ sky130_fd_sc_hd__xor2_1
X_12799_ _05047_ _05071_ VGND VGND VPWR VPWR _05072_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_50_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17326_ net6733 net7890 VGND VGND VPWR VPWR _09240_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_172_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14538_ net726 _06703_ VGND VGND VPWR VPWR _06717_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17257_ net2959 net155 net2162 net9129 VGND VGND VPWR VPWR _00355_ sky130_fd_sc_hd__a22o_1
X_14469_ net9072 net831 net1292 _06656_ VGND VGND VPWR VPWR _00101_ sky130_fd_sc_hd__a22o_1
XFILLER_0_181_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16208_ _08271_ _08272_ VGND VGND VPWR VPWR _08273_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_141_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17188_ net1922 _09138_ VGND VGND VPWR VPWR _09139_ sky130_fd_sc_hd__nor2_1
X_16139_ net1089 net983 VGND VGND VPWR VPWR _08205_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19829_ _11545_ _11662_ VGND VGND VPWR VPWR _11663_ sky130_fd_sc_hd__nor2_1
X_22840_ _02737_ _02738_ VGND VGND VPWR VPWR _02740_ sky130_fd_sc_hd__or2_1
XFILLER_0_190_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22771_ net4302 net8932 VGND VGND VPWR VPWR _02692_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24510_ _04272_ _04276_ _04277_ VGND VGND VPWR VPWR _04367_ sky130_fd_sc_hd__o21ba_1
X_21722_ _01730_ _01731_ VGND VGND VPWR VPWR _01733_ sky130_fd_sc_hd__or2_1
X_25490_ clknet_leaf_47_clk _00370_ net8778 VGND VGND VPWR VPWR svm0.tA\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_166_Right_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8107 net82 VGND VGND VPWR VPWR net8107 sky130_fd_sc_hd__clkbuf_1
X_24441_ net4544 net4824 VGND VGND VPWR VPWR _04299_ sky130_fd_sc_hd__nand2_1
X_21653_ _01662_ _01663_ VGND VGND VPWR VPWR _01664_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_136_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8118 net74 VGND VGND VPWR VPWR net8118 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8129 net8130 VGND VGND VPWR VPWR net8129 sky130_fd_sc_hd__clkbuf_1
X_20604_ _12367_ VGND VGND VPWR VPWR _12385_ sky130_fd_sc_hd__inv_2
Xwire7406 net7407 VGND VGND VPWR VPWR net7406 sky130_fd_sc_hd__clkbuf_1
X_24372_ net4789 _04230_ VGND VGND VPWR VPWR _04231_ sky130_fd_sc_hd__xnor2_1
X_21584_ _01472_ _01474_ _01470_ VGND VGND VPWR VPWR _01596_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_46_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7417 matmul0.matmul_stage_inst.c\[2\] VGND VGND VPWR VPWR net7417 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length3115 net3116 VGND VGND VPWR VPWR net3115 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7439 net7436 VGND VGND VPWR VPWR net7439 sky130_fd_sc_hd__buf_1
X_23323_ net4926 net4743 _03191_ _03192_ VGND VGND VPWR VPWR _03193_ sky130_fd_sc_hd__a31oi_2
Xfanout5909 net5912 VGND VGND VPWR VPWR net5909 sky130_fd_sc_hd__buf_1
X_20535_ _12305_ _12309_ _12320_ VGND VGND VPWR VPWR _12321_ sky130_fd_sc_hd__a21oi_1
Xwire6716 net6717 VGND VGND VPWR VPWR net6716 sky130_fd_sc_hd__buf_1
Xwire6727 net6729 VGND VGND VPWR VPWR net6727 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6738 svm0.counter\[1\] VGND VGND VPWR VPWR net6738 sky130_fd_sc_hd__buf_1
XFILLER_0_162_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6749 net6750 VGND VGND VPWR VPWR net6749 sky130_fd_sc_hd__buf_1
X_23254_ _03121_ _03122_ _03123_ VGND VGND VPWR VPWR _03124_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2447 net2448 VGND VGND VPWR VPWR net2447 sky130_fd_sc_hd__buf_1
X_20466_ cordic0.slte0.opA\[15\] _12249_ VGND VGND VPWR VPWR _12257_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length1724 _01539_ VGND VGND VPWR VPWR net1724 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22205_ pid_d.mult0.a\[9\] net5658 VGND VGND VPWR VPWR _02210_ sky130_fd_sc_hd__nand2b_1
X_23185_ net5065 net4757 VGND VGND VPWR VPWR _03055_ sky130_fd_sc_hd__nand2_1
X_20397_ net6467 net4037 _12175_ _12194_ _12098_ VGND VGND VPWR VPWR _12195_ sky130_fd_sc_hd__o311a_1
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22136_ _02039_ _02041_ _02040_ VGND VGND VPWR VPWR _02142_ sky130_fd_sc_hd__o21a_1
XFILLER_0_100_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22067_ net1045 net1170 _02073_ VGND VGND VPWR VPWR _02074_ sky130_fd_sc_hd__a21oi_1
Xwire1001 _05359_ VGND VGND VPWR VPWR net1001 sky130_fd_sc_hd__buf_1
Xwire1012 _04236_ VGND VGND VPWR VPWR net1012 sky130_fd_sc_hd__buf_1
X_21018_ net5541 net5930 VGND VGND VPWR VPWR _01034_ sky130_fd_sc_hd__nand2_1
Xwire1023 _03466_ VGND VGND VPWR VPWR net1023 sky130_fd_sc_hd__clkbuf_1
Xwire1034 net1035 VGND VGND VPWR VPWR net1034 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1045 _01954_ VGND VGND VPWR VPWR net1045 sky130_fd_sc_hd__buf_2
Xwire1056 _11570_ VGND VGND VPWR VPWR net1056 sky130_fd_sc_hd__clkbuf_2
X_13840_ _06057_ _06058_ _06106_ VGND VGND VPWR VPWR _06107_ sky130_fd_sc_hd__nand3_1
X_25826_ clknet_leaf_36_clk _00699_ net8750 VGND VGND VPWR VPWR pid_q.curr_error\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1067 net1068 VGND VGND VPWR VPWR net1067 sky130_fd_sc_hd__clkbuf_1
Xwire1078 net1079 VGND VGND VPWR VPWR net1078 sky130_fd_sc_hd__clkbuf_2
Xwire1089 net1090 VGND VGND VPWR VPWR net1089 sky130_fd_sc_hd__buf_1
X_13771_ _06035_ _06038_ VGND VGND VPWR VPWR _06039_ sky130_fd_sc_hd__xnor2_1
X_25757_ clknet_leaf_13_clk _00630_ net8608 VGND VGND VPWR VPWR pid_d.kp\[15\] sky130_fd_sc_hd__dfrtp_1
X_22969_ _02852_ VGND VGND VPWR VPWR _00651_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_186_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15510_ net1859 _07582_ VGND VGND VPWR VPWR _07583_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24708_ net8028 net5299 VGND VGND VPWR VPWR _04544_ sky130_fd_sc_hd__or2b_1
X_12722_ _04986_ _04987_ VGND VGND VPWR VPWR _04995_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16490_ _08521_ _08532_ _08549_ VGND VGND VPWR VPWR _08550_ sky130_fd_sc_hd__o21a_1
X_25688_ clknet_leaf_5_clk _00561_ net8567 VGND VGND VPWR VPWR pid_d.curr_error\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_133_Right_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15441_ net6616 matmul0.matmul_stage_inst.b\[13\] matmul0.matmul_stage_inst.a\[13\]
+ net6581 VGND VGND VPWR VPWR _07515_ sky130_fd_sc_hd__a22o_1
XFILLER_0_194_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24639_ _04414_ _04421_ VGND VGND VPWR VPWR _04494_ sky130_fd_sc_hd__and2b_1
X_12653_ net2341 VGND VGND VPWR VPWR _04926_ sky130_fd_sc_hd__buf_1
XFILLER_0_183_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout7812 svm0.periodTop\[5\] VGND VGND VPWR VPWR net7812 sky130_fd_sc_hd__buf_1
XFILLER_0_37_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8630 net8632 VGND VGND VPWR VPWR net8630 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_183_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18160_ _09747_ _09760_ VGND VGND VPWR VPWR _10011_ sky130_fd_sc_hd__xor2_1
Xwire8641 net8644 VGND VGND VPWR VPWR net8641 sky130_fd_sc_hd__clkbuf_1
Xmax_length5073 net5074 VGND VGND VPWR VPWR net5073 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15372_ _07443_ _07445_ VGND VGND VPWR VPWR _07446_ sky130_fd_sc_hd__or2_1
X_12584_ _04868_ VGND VGND VPWR VPWR _04869_ sky130_fd_sc_hd__buf_1
Xfanout7856 svm0.periodTop\[3\] VGND VGND VPWR VPWR net7856 sky130_fd_sc_hd__buf_1
Xmax_length5095 net5096 VGND VGND VPWR VPWR net5095 sky130_fd_sc_hd__buf_1
Xwire8663 net8661 VGND VGND VPWR VPWR net8663 sky130_fd_sc_hd__clkbuf_2
X_17111_ net3307 net1233 _09065_ _09067_ VGND VGND VPWR VPWR _00332_ sky130_fd_sc_hd__a31o_1
XFILLER_0_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire320 _06019_ VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__buf_1
Xfanout7878 net7884 VGND VGND VPWR VPWR net7878 sky130_fd_sc_hd__buf_1
Xwire8674 net8675 VGND VGND VPWR VPWR net8674 sky130_fd_sc_hd__buf_1
X_14323_ _06544_ VGND VGND VPWR VPWR _00067_ sky130_fd_sc_hd__clkbuf_1
Xwire8685 net8684 VGND VGND VPWR VPWR net8685 sky130_fd_sc_hd__buf_1
Xwire7940 net7941 VGND VGND VPWR VPWR net7940 sky130_fd_sc_hd__buf_1
Xwire331 net332 VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__clkbuf_1
X_18091_ _09930_ _09940_ _09941_ VGND VGND VPWR VPWR _09942_ sky130_fd_sc_hd__a21oi_1
Xwire7951 net7952 VGND VGND VPWR VPWR net7951 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire342 net343 VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7962 net7963 VGND VGND VPWR VPWR net7962 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7973 pid_q.target\[12\] VGND VGND VPWR VPWR net7973 sky130_fd_sc_hd__buf_1
Xwire353 _08732_ VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__clkbuf_1
X_17042_ net1831 _09001_ net8043 VGND VGND VPWR VPWR _09002_ sky130_fd_sc_hd__o21a_1
Xwire364 net365 VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7984 pid_q.target\[10\] VGND VGND VPWR VPWR net7984 sky130_fd_sc_hd__clkbuf_1
X_14254_ net1916 VGND VGND VPWR VPWR _06509_ sky130_fd_sc_hd__buf_1
XFILLER_0_20_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire386 net387 VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__buf_1
XFILLER_0_123_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire397 net398 VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__clkbuf_1
X_13205_ net919 _05476_ _05357_ VGND VGND VPWR VPWR _05478_ sky130_fd_sc_hd__o21a_1
X_14185_ _06443_ _06444_ VGND VGND VPWR VPWR _06445_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13136_ _05342_ net2303 _05407_ _05408_ VGND VGND VPWR VPWR _05409_ sky130_fd_sc_hd__o211ai_1
X_18993_ net6314 net6343 net6293 VGND VGND VPWR VPWR _10830_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_178_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13067_ net7877 _05191_ VGND VGND VPWR VPWR _05340_ sky130_fd_sc_hd__nand2_1
X_17944_ net6941 VGND VGND VPWR VPWR _09795_ sky130_fd_sc_hd__inv_2
X_17875_ _09723_ _09603_ VGND VGND VPWR VPWR _09726_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2280 net2281 VGND VGND VPWR VPWR net2280 sky130_fd_sc_hd__buf_1
XFILLER_0_75_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2291 net2292 VGND VGND VPWR VPWR net2291 sky130_fd_sc_hd__buf_1
X_19614_ net6088 net6103 VGND VGND VPWR VPWR _11451_ sky130_fd_sc_hd__nand2_1
X_16826_ net6430 matmul0.sin\[1\] net3365 VGND VGND VPWR VPWR _08804_ sky130_fd_sc_hd__mux2_1
Xwire1590 net1591 VGND VGND VPWR VPWR net1590 sky130_fd_sc_hd__buf_1
XFILLER_0_159_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19545_ net3870 VGND VGND VPWR VPWR _11382_ sky130_fd_sc_hd__buf_1
X_16757_ _08767_ VGND VGND VPWR VPWR _00278_ sky130_fd_sc_hd__clkbuf_1
X_13969_ _06224_ _06233_ VGND VGND VPWR VPWR _06234_ sky130_fd_sc_hd__xnor2_2
X_15708_ net2804 net3481 VGND VGND VPWR VPWR _07779_ sky130_fd_sc_hd__nor2_1
XFILLER_0_158_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19476_ net6299 _11265_ _10984_ VGND VGND VPWR VPWR _11313_ sky130_fd_sc_hd__a21oi_1
X_16688_ matmul0.matmul_stage_inst.mult2\[10\] matmul0.matmul_stage_inst.mult1\[10\]
+ VGND VGND VPWR VPWR _08719_ sky130_fd_sc_hd__xor2_1
XFILLER_0_152_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15639_ _07590_ _07625_ net889 VGND VGND VPWR VPWR _07711_ sky130_fd_sc_hd__a21o_1
X_18427_ net6809 _10276_ VGND VGND VPWR VPWR _10277_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18358_ _10175_ net2543 VGND VGND VPWR VPWR _10209_ sky130_fd_sc_hd__nand2_1
XFILLER_0_173_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17309_ svm0.counter\[8\] VGND VGND VPWR VPWR _09223_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18289_ net3245 net1215 net1447 VGND VGND VPWR VPWR _10140_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20320_ cordic0.slte0.opA\[2\] _12112_ VGND VGND VPWR VPWR _12124_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20251_ net15 _12061_ VGND VGND VPWR VPWR _12065_ sky130_fd_sc_hd__and2_1
Xwire3909 _10794_ VGND VGND VPWR VPWR net3909 sky130_fd_sc_hd__buf_1
X_20182_ net2580 _12007_ _11941_ VGND VGND VPWR VPWR _12008_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24990_ pid_q.kp\[14\] _04730_ net1635 VGND VGND VPWR VPWR _04750_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23941_ net5155 _03804_ _03698_ _03703_ VGND VGND VPWR VPWR _03805_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_193_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23872_ _03629_ _03635_ _03634_ VGND VGND VPWR VPWR _03737_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25611_ clknet_leaf_108_clk _00484_ net8349 VGND VGND VPWR VPWR cordic0.slte0.opA\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_193_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22823_ _02723_ _02724_ VGND VGND VPWR VPWR _02725_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25542_ clknet_leaf_29_clk _00422_ net8674 VGND VGND VPWR VPWR pid_q.prev_int\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_22754_ pid_d.ki\[9\] net3070 net1696 VGND VGND VPWR VPWR _02681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21705_ _01714_ _01715_ VGND VGND VPWR VPWR _01716_ sky130_fd_sc_hd__or2_1
X_25473_ clknet_leaf_46_clk _00353_ net8774 VGND VGND VPWR VPWR svm0.tB\[11\] sky130_fd_sc_hd__dfrtp_1
X_22685_ _02631_ net5563 net2447 VGND VGND VPWR VPWR _02632_ sky130_fd_sc_hd__mux2_1
X_24424_ net4994 _04216_ _04214_ VGND VGND VPWR VPWR _04282_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21636_ pid_d.curr_int\[5\] pid_d.prev_int\[5\] VGND VGND VPWR VPWR _01647_ sky130_fd_sc_hd__xor2_1
Xwire7203 net7204 VGND VGND VPWR VPWR net7203 sky130_fd_sc_hd__buf_1
Xwire7214 net7215 VGND VGND VPWR VPWR net7214 sky130_fd_sc_hd__clkbuf_2
Xwire7225 net7226 VGND VGND VPWR VPWR net7225 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7236 matmul0.alpha_pass\[12\] VGND VGND VPWR VPWR net7236 sky130_fd_sc_hd__buf_1
XFILLER_0_62_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24355_ net4960 net4937 net3041 VGND VGND VPWR VPWR _04214_ sky130_fd_sc_hd__o21a_1
Xwire6502 net6501 VGND VGND VPWR VPWR net6502 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout5706 net5715 VGND VGND VPWR VPWR net5706 sky130_fd_sc_hd__clkbuf_1
X_21567_ _01455_ _01457_ _01578_ VGND VGND VPWR VPWR _01579_ sky130_fd_sc_hd__a21oi_2
Xwire7258 net7249 VGND VGND VPWR VPWR net7258 sky130_fd_sc_hd__buf_1
Xwire7269 net7270 VGND VGND VPWR VPWR net7269 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23306_ _02968_ _03175_ VGND VGND VPWR VPWR _03176_ sky130_fd_sc_hd__nor2_1
Xfanout5739 net5756 VGND VGND VPWR VPWR net5739 sky130_fd_sc_hd__buf_1
XFILLER_0_144_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5801 net5798 VGND VGND VPWR VPWR net5801 sky130_fd_sc_hd__buf_1
X_20518_ net1053 _12303_ VGND VGND VPWR VPWR _12305_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6546 net6544 VGND VGND VPWR VPWR net6546 sky130_fd_sc_hd__buf_1
X_24286_ net4959 _03605_ _04145_ VGND VGND VPWR VPWR _04146_ sky130_fd_sc_hd__a21o_1
Xwire5812 net5813 VGND VGND VPWR VPWR net5812 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_16_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21498_ net5894 _01507_ _01509_ _01510_ _01508_ VGND VGND VPWR VPWR _01511_ sky130_fd_sc_hd__a32o_1
Xwire6557 net6558 VGND VGND VPWR VPWR net6557 sky130_fd_sc_hd__buf_1
Xmax_length1510 _08251_ VGND VGND VPWR VPWR net1510 sky130_fd_sc_hd__clkbuf_1
Xwire5823 net5824 VGND VGND VPWR VPWR net5823 sky130_fd_sc_hd__buf_1
Xwire6568 net6569 VGND VGND VPWR VPWR net6568 sky130_fd_sc_hd__buf_1
Xwire5834 net5835 VGND VGND VPWR VPWR net5834 sky130_fd_sc_hd__clkbuf_1
Xwire6579 matmul0.matmul_stage_inst.state\[5\] VGND VGND VPWR VPWR net6579 sky130_fd_sc_hd__clkbuf_1
Xmax_length2277 _06517_ VGND VGND VPWR VPWR net2277 sky130_fd_sc_hd__clkbuf_1
X_23237_ _03105_ _03106_ VGND VGND VPWR VPWR _03107_ sky130_fd_sc_hd__xnor2_2
X_20449_ net6370 _12232_ net6369 VGND VGND VPWR VPWR _12242_ sky130_fd_sc_hd__a21oi_1
Xwire5845 net5846 VGND VGND VPWR VPWR net5845 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5889 net5890 VGND VGND VPWR VPWR net5889 sky130_fd_sc_hd__clkbuf_1
X_23168_ _03035_ _03037_ VGND VGND VPWR VPWR _03038_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22119_ _02123_ _02124_ VGND VGND VPWR VPWR _02125_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23099_ net5037 net4693 VGND VGND VPWR VPWR _02969_ sky130_fd_sc_hd__nand2_1
X_15990_ net4068 _08055_ _08056_ _08053_ _08057_ VGND VGND VPWR VPWR _08058_ sky130_fd_sc_hd__o221a_1
X_14941_ net4153 net4148 VGND VGND VPWR VPWR _07015_ sky130_fd_sc_hd__or2_1
X_17660_ svm0.tA\[6\] net6725 VGND VGND VPWR VPWR _09540_ sky130_fd_sc_hd__and2b_1
X_14872_ net7184 matmul0.matmul_stage_inst.f\[8\] net3606 VGND VGND VPWR VPWR _06954_
+ sky130_fd_sc_hd__mux2_1
X_16611_ _08655_ VGND VGND VPWR VPWR _00244_ sky130_fd_sc_hd__clkbuf_1
X_13823_ _06050_ net840 VGND VGND VPWR VPWR _06090_ sky130_fd_sc_hd__nand2_1
X_25809_ clknet_leaf_38_clk _00682_ net8755 VGND VGND VPWR VPWR pid_q.prev_error\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_17591_ net6689 svm0.tB\[14\] VGND VGND VPWR VPWR _09472_ sky130_fd_sc_hd__and2b_1
XFILLER_0_173_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19330_ _11156_ _11160_ _11166_ VGND VGND VPWR VPWR _11167_ sky130_fd_sc_hd__o21a_1
X_16542_ net2744 net2245 VGND VGND VPWR VPWR _08601_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13754_ _05979_ net727 VGND VGND VPWR VPWR _06022_ sky130_fd_sc_hd__or2_1
X_12705_ _04945_ _04953_ VGND VGND VPWR VPWR _04978_ sky130_fd_sc_hd__xnor2_2
X_19261_ _11034_ net3180 _11038_ VGND VGND VPWR VPWR _11098_ sky130_fd_sc_hd__o21ba_1
X_16473_ _08504_ _08533_ VGND VGND VPWR VPWR _08534_ sky130_fd_sc_hd__xnor2_1
X_13685_ _05942_ _05953_ VGND VGND VPWR VPWR _05954_ sky130_fd_sc_hd__xnor2_2
Xfanout8343 net8348 VGND VGND VPWR VPWR net8343 sky130_fd_sc_hd__buf_1
XFILLER_0_122_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18212_ net3947 VGND VGND VPWR VPWR _10063_ sky130_fd_sc_hd__buf_1
X_15424_ net2229 net1866 _07497_ VGND VGND VPWR VPWR _07498_ sky130_fd_sc_hd__a21o_1
X_12636_ _04894_ VGND VGND VPWR VPWR _04909_ sky130_fd_sc_hd__clkbuf_1
X_19192_ net6312 _10843_ VGND VGND VPWR VPWR _11029_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8398 net8411 VGND VGND VPWR VPWR net8398 sky130_fd_sc_hd__clkbuf_2
X_18143_ _09901_ _09941_ _09945_ net2548 VGND VGND VPWR VPWR _09994_ sky130_fd_sc_hd__a31o_1
Xwire8460 net8461 VGND VGND VPWR VPWR net8460 sky130_fd_sc_hd__buf_1
X_15355_ _07315_ _07322_ VGND VGND VPWR VPWR _07429_ sky130_fd_sc_hd__xnor2_1
X_12567_ _04856_ VGND VGND VPWR VPWR _04857_ sky130_fd_sc_hd__buf_1
XFILLER_0_142_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8482 net8479 VGND VGND VPWR VPWR net8482 sky130_fd_sc_hd__clkbuf_1
Xfanout6952 net6960 VGND VGND VPWR VPWR net6952 sky130_fd_sc_hd__clkbuf_1
Xwire8493 net8494 VGND VGND VPWR VPWR net8493 sky130_fd_sc_hd__buf_1
X_14306_ net8312 net3645 VGND VGND VPWR VPWR _06528_ sky130_fd_sc_hd__and2_1
Xwire7770 net7769 VGND VGND VPWR VPWR net7770 sky130_fd_sc_hd__buf_1
X_18074_ _09906_ _09907_ _09849_ VGND VGND VPWR VPWR _09925_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire161 net162 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_1
Xwire7781 net7782 VGND VGND VPWR VPWR net7781 sky130_fd_sc_hd__clkbuf_1
X_15286_ net3559 net2768 VGND VGND VPWR VPWR _07360_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7792 net7793 VGND VGND VPWR VPWR net7792 sky130_fd_sc_hd__buf_1
Xfanout6985 cordic0.vec\[1\]\[7\] VGND VGND VPWR VPWR net6985 sky130_fd_sc_hd__clkbuf_1
Xwire172 net173 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_1
Xhold208 svm0.tC\[8\] VGND VGND VPWR VPWR net9161 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire183 net184 VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_1
Xhold219 svm0.tA\[10\] VGND VGND VPWR VPWR net9172 sky130_fd_sc_hd__dlygate4sd3_1
Xwire194 _04814_ VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_1
X_17025_ _08984_ VGND VGND VPWR VPWR _08985_ sky130_fd_sc_hd__buf_1
X_14237_ _06446_ _06481_ VGND VGND VPWR VPWR _06494_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14168_ _06426_ _06428_ _06369_ VGND VGND VPWR VPWR _06429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13119_ net7736 _05012_ _05250_ VGND VGND VPWR VPWR _05392_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14099_ net255 net254 VGND VGND VPWR VPWR _06362_ sky130_fd_sc_hd__nand2_1
X_18976_ net6314 net6339 VGND VGND VPWR VPWR _10813_ sky130_fd_sc_hd__and2b_1
X_17927_ _09734_ VGND VGND VPWR VPWR _09778_ sky130_fd_sc_hd__inv_2
XFILLER_0_147_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17858_ net7028 net7105 VGND VGND VPWR VPWR _09709_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_163_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16809_ net9038 matmul0.cos\[7\] net3367 VGND VGND VPWR VPWR _08795_ sky130_fd_sc_hd__mux2_1
X_17789_ net2563 _09639_ VGND VGND VPWR VPWR _09640_ sky130_fd_sc_hd__xnor2_2
X_19528_ _11307_ _11306_ VGND VGND VPWR VPWR _11365_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19459_ _10974_ net2521 VGND VGND VPWR VPWR _11296_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22470_ net2056 _02469_ _02470_ _02446_ _02441_ VGND VGND VPWR VPWR _02471_ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21421_ _04875_ net2478 _01427_ _01434_ VGND VGND VPWR VPWR _01435_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24140_ _03978_ _04001_ VGND VGND VPWR VPWR _04002_ sky130_fd_sc_hd__xnor2_1
X_21352_ _01293_ _01294_ _01365_ VGND VGND VPWR VPWR _01366_ sky130_fd_sc_hd__a21oi_2
Xwire5108 net5109 VGND VGND VPWR VPWR net5108 sky130_fd_sc_hd__buf_1
XFILLER_0_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5119 net5121 VGND VGND VPWR VPWR net5119 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20303_ net6516 net1481 _12106_ _12107_ _12092_ VGND VGND VPWR VPWR _12108_ sky130_fd_sc_hd__a32o_1
XFILLER_0_130_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24071_ _03932_ _03933_ VGND VGND VPWR VPWR _03934_ sky130_fd_sc_hd__nand2_1
X_21283_ _01292_ _01297_ VGND VGND VPWR VPWR _01298_ sky130_fd_sc_hd__xor2_1
Xwire4407 net4408 VGND VGND VPWR VPWR net4407 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4429 pid_q.out\[9\] VGND VGND VPWR VPWR net4429 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23022_ net4982 net4694 VGND VGND VPWR VPWR _02892_ sky130_fd_sc_hd__nand2_1
X_20234_ net12 _12051_ VGND VGND VPWR VPWR _12052_ sky130_fd_sc_hd__xnor2_1
Xwire3706 net3707 VGND VGND VPWR VPWR net3706 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire3717 _04867_ VGND VGND VPWR VPWR net3717 sky130_fd_sc_hd__clkbuf_1
Xwire3728 net3729 VGND VGND VPWR VPWR net3728 sky130_fd_sc_hd__clkbuf_1
Xwire3739 net3740 VGND VGND VPWR VPWR net3739 sky130_fd_sc_hd__buf_1
X_20165_ _11934_ VGND VGND VPWR VPWR _11991_ sky130_fd_sc_hd__inv_2
X_24973_ _04741_ VGND VGND VPWR VPWR _00766_ sky130_fd_sc_hd__clkbuf_1
X_20096_ _11923_ _11924_ net1438 VGND VGND VPWR VPWR _11925_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_196_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23924_ _03716_ _03718_ _03787_ VGND VGND VPWR VPWR _03788_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_58_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length7701 net7702 VGND VGND VPWR VPWR net7701 sky130_fd_sc_hd__clkbuf_1
X_23855_ _03716_ _03719_ VGND VGND VPWR VPWR _03720_ sky130_fd_sc_hd__xnor2_1
Xmax_length7712 net7713 VGND VGND VPWR VPWR net7712 sky130_fd_sc_hd__clkbuf_1
Xmax_length7723 net7722 VGND VGND VPWR VPWR net7723 sky130_fd_sc_hd__clkbuf_1
X_22806_ pid_d.kp\[15\] _02692_ net2036 VGND VGND VPWR VPWR _02711_ sky130_fd_sc_hd__mux2_1
X_23786_ net855 _03651_ VGND VGND VPWR VPWR _03652_ sky130_fd_sc_hd__xnor2_2
X_20998_ _00995_ _01004_ net1051 VGND VGND VPWR VPWR _01014_ sky130_fd_sc_hd__o21a_1
XFILLER_0_156_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25525_ clknet_leaf_35_clk _00405_ net8758 VGND VGND VPWR VPWR svm0.counter\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_22737_ _02669_ VGND VGND VPWR VPWR _00602_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13470_ net1131 _05588_ _05742_ VGND VGND VPWR VPWR _05743_ sky130_fd_sc_hd__a21oi_2
X_25456_ clknet_leaf_100_clk _00339_ net8368 VGND VGND VPWR VPWR cordic0.vec\[1\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22668_ net3098 VGND VGND VPWR VPWR _02620_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout6204 net6206 VGND VGND VPWR VPWR net6204 sky130_fd_sc_hd__buf_1
Xwire7000 net6998 VGND VGND VPWR VPWR net7000 sky130_fd_sc_hd__buf_1
XFILLER_0_180_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7011 net7008 VGND VGND VPWR VPWR net7011 sky130_fd_sc_hd__buf_1
X_24407_ net588 net587 VGND VGND VPWR VPWR _04265_ sky130_fd_sc_hd__nor2_1
Xfanout6215 net6239 VGND VGND VPWR VPWR net6215 sky130_fd_sc_hd__buf_1
XFILLER_0_36_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21619_ _01628_ net701 VGND VGND VPWR VPWR _01631_ sky130_fd_sc_hd__or2_1
XFILLER_0_180_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25387_ clknet_leaf_73_clk _00270_ net8473 VGND VGND VPWR VPWR matmul0.b\[6\] sky130_fd_sc_hd__dfrtp_1
X_22599_ net4226 _02569_ VGND VGND VPWR VPWR _02575_ sky130_fd_sc_hd__or2_1
Xwire7044 net7045 VGND VGND VPWR VPWR net7044 sky130_fd_sc_hd__clkbuf_1
Xwire7055 net7057 VGND VGND VPWR VPWR net7055 sky130_fd_sc_hd__buf_1
Xwire6310 net6306 VGND VGND VPWR VPWR net6310 sky130_fd_sc_hd__buf_1
X_15140_ net1889 _07211_ VGND VGND VPWR VPWR _07214_ sky130_fd_sc_hd__xor2_1
X_24338_ net376 _04192_ _04193_ _04196_ VGND VGND VPWR VPWR _04197_ sky130_fd_sc_hd__a31o_1
Xwire7077 net7078 VGND VGND VPWR VPWR net7077 sky130_fd_sc_hd__buf_1
XFILLER_0_23_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7088 net7086 VGND VGND VPWR VPWR net7088 sky130_fd_sc_hd__buf_1
Xwire6343 net6341 VGND VGND VPWR VPWR net6343 sky130_fd_sc_hd__buf_1
Xwire6354 net6353 VGND VGND VPWR VPWR net6354 sky130_fd_sc_hd__buf_1
Xwire7099 net7096 VGND VGND VPWR VPWR net7099 sky130_fd_sc_hd__buf_1
XFILLER_0_121_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6365 net6366 VGND VGND VPWR VPWR net6365 sky130_fd_sc_hd__clkbuf_1
Xwire5631 net5630 VGND VGND VPWR VPWR net5631 sky130_fd_sc_hd__buf_1
XFILLER_0_26_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15071_ net4098 net4096 VGND VGND VPWR VPWR _07145_ sky130_fd_sc_hd__or2_1
Xwire6376 net6375 VGND VGND VPWR VPWR net6376 sky130_fd_sc_hd__clkbuf_2
X_24269_ _04061_ _04063_ _04062_ VGND VGND VPWR VPWR _04129_ sky130_fd_sc_hd__o21ai_1
Xwire5642 net5643 VGND VGND VPWR VPWR net5642 sky130_fd_sc_hd__buf_1
Xwire6387 net6388 VGND VGND VPWR VPWR net6387 sky130_fd_sc_hd__clkbuf_1
Xwire5653 net5654 VGND VGND VPWR VPWR net5653 sky130_fd_sc_hd__buf_1
Xwire6398 cordic0.slte0.opB\[13\] VGND VGND VPWR VPWR net6398 sky130_fd_sc_hd__clkbuf_1
X_14022_ net7702 net1324 _06230_ VGND VGND VPWR VPWR _06286_ sky130_fd_sc_hd__a21o_1
Xwire5664 net5665 VGND VGND VPWR VPWR net5664 sky130_fd_sc_hd__clkbuf_1
Xwire4930 net4931 VGND VGND VPWR VPWR net4930 sky130_fd_sc_hd__clkbuf_1
Xwire5675 net5676 VGND VGND VPWR VPWR net5675 sky130_fd_sc_hd__clkbuf_1
Xfanout4879 pid_q.mult0.b\[11\] VGND VGND VPWR VPWR net4879 sky130_fd_sc_hd__buf_1
Xwire4941 net4942 VGND VGND VPWR VPWR net4941 sky130_fd_sc_hd__buf_1
Xwire5686 net5688 VGND VGND VPWR VPWR net5686 sky130_fd_sc_hd__buf_1
Xwire5697 net5698 VGND VGND VPWR VPWR net5697 sky130_fd_sc_hd__buf_1
Xwire4963 net4964 VGND VGND VPWR VPWR net4963 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4974 net4975 VGND VGND VPWR VPWR net4974 sky130_fd_sc_hd__clkbuf_1
X_18830_ net6837 _10638_ _10672_ VGND VGND VPWR VPWR _10673_ sky130_fd_sc_hd__nand3_1
Xwire4985 net4986 VGND VGND VPWR VPWR net4985 sky130_fd_sc_hd__clkbuf_1
X_15973_ net2722 net2624 VGND VGND VPWR VPWR _08041_ sky130_fd_sc_hd__nor2_1
X_18761_ _10516_ net764 _10605_ VGND VGND VPWR VPWR _10606_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17712_ net9207 net1217 net1451 pid_q.curr_int\[3\] VGND VGND VPWR VPWR _00417_ sky130_fd_sc_hd__a22o_1
X_14924_ net6545 net6585 net7392 VGND VGND VPWR VPWR _06998_ sky130_fd_sc_hd__o21a_1
XFILLER_0_101_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18692_ net6863 net2588 VGND VGND VPWR VPWR _10538_ sky130_fd_sc_hd__nand2_1
XFILLER_0_188_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold80 matmul0.matmul_stage_inst.b\[3\] VGND VGND VPWR VPWR net9033 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 matmul0.matmul_stage_inst.d\[11\] VGND VGND VPWR VPWR net9044 sky130_fd_sc_hd__dlygate4sd3_1
X_17643_ net4004 svm0.tA\[13\] VGND VGND VPWR VPWR _09523_ sky130_fd_sc_hd__nor2_1
X_14855_ matmul0.b\[0\] matmul0.matmul_stage_inst.f\[0\] net3609 VGND VGND VPWR VPWR
+ _06945_ sky130_fd_sc_hd__mux2_1
X_13806_ _06064_ _06073_ VGND VGND VPWR VPWR _06074_ sky130_fd_sc_hd__xor2_1
X_17574_ net4012 svm0.tC\[1\] svm0.tC\[0\] net4033 VGND VGND VPWR VPWR _09456_ sky130_fd_sc_hd__a211o_1
XFILLER_0_98_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14786_ net3613 _06908_ VGND VGND VPWR VPWR _06909_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19313_ net3918 net2511 VGND VGND VPWR VPWR _11150_ sky130_fd_sc_hd__xnor2_2
X_16525_ _08524_ _08530_ _08584_ VGND VGND VPWR VPWR _08585_ sky130_fd_sc_hd__o21ai_2
X_13737_ _05866_ net451 VGND VGND VPWR VPWR _06006_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_70_clk clknet_4_8__leaf_clk VGND VGND VPWR VPWR clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_16
X_19244_ _10821_ net3210 _11080_ VGND VGND VPWR VPWR _11081_ sky130_fd_sc_hd__a21oi_1
X_16456_ _08454_ _08516_ net2245 VGND VGND VPWR VPWR _08517_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_183_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13668_ _05895_ _05916_ _05917_ VGND VGND VPWR VPWR _05937_ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15407_ _07479_ _07480_ VGND VGND VPWR VPWR _07481_ sky130_fd_sc_hd__xor2_1
X_12619_ _04856_ VGND VGND VPWR VPWR _04892_ sky130_fd_sc_hd__buf_6
X_19175_ _10963_ VGND VGND VPWR VPWR _11012_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16387_ net2623 net2631 VGND VGND VPWR VPWR _08449_ sky130_fd_sc_hd__nor2_1
X_13599_ _05866_ _05868_ VGND VGND VPWR VPWR _05869_ sky130_fd_sc_hd__nor2_1
Xfanout7483 pid_q.state\[3\] VGND VGND VPWR VPWR net7483 sky130_fd_sc_hd__buf_1
Xwire8290 net8291 VGND VGND VPWR VPWR net8290 sky130_fd_sc_hd__clkbuf_1
X_18126_ net7038 _09976_ VGND VGND VPWR VPWR _09977_ sky130_fd_sc_hd__nand2_1
X_15338_ net2740 _07224_ VGND VGND VPWR VPWR _07412_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6782 net6786 VGND VGND VPWR VPWR net6782 sky130_fd_sc_hd__buf_1
XFILLER_0_13_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18057_ _09906_ _09907_ VGND VGND VPWR VPWR _09908_ sky130_fd_sc_hd__nand2_1
X_15269_ _07008_ net1286 VGND VGND VPWR VPWR _07343_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17008_ _08825_ VGND VGND VPWR VPWR _08969_ sky130_fd_sc_hd__buf_1
XFILLER_0_158_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18959_ net6248 net6231 VGND VGND VPWR VPWR _10796_ sky130_fd_sc_hd__and2b_2
X_21970_ net1047 net1171 VGND VGND VPWR VPWR _01978_ sky130_fd_sc_hd__or2_1
X_20921_ _00926_ net1186 VGND VGND VPWR VPWR _00937_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23640_ _03432_ _03437_ _03506_ VGND VGND VPWR VPWR _03507_ sky130_fd_sc_hd__a21o_1
Xmax_length6318 net6319 VGND VGND VPWR VPWR net6318 sky130_fd_sc_hd__buf_1
X_20852_ net5492 _00867_ VGND VGND VPWR VPWR _00868_ sky130_fd_sc_hd__nand2_1
XFILLER_0_178_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length5606 net5607 VGND VGND VPWR VPWR net5606 sky130_fd_sc_hd__buf_1
XFILLER_0_190_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23571_ _03430_ _03438_ VGND VGND VPWR VPWR _03439_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20783_ net5596 net5776 net5794 net5578 VGND VGND VPWR VPWR _12554_ sky130_fd_sc_hd__a22oi_1
Xclkbuf_leaf_61_clk clknet_4_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25310_ clknet_leaf_76_clk _00193_ net8462 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.e\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_22522_ net2050 VGND VGND VPWR VPWR _02522_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire908 _06123_ VGND VGND VPWR VPWR net908 sky130_fd_sc_hd__clkbuf_1
X_25241_ clknet_leaf_89_clk _00124_ net8421 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.a\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire919 _05356_ VGND VGND VPWR VPWR net919 sky130_fd_sc_hd__dlymetal6s2s_1
X_22453_ net520 net597 VGND VGND VPWR VPWR _02455_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21404_ net1050 _01313_ _01417_ VGND VGND VPWR VPWR _01418_ sky130_fd_sc_hd__o21a_2
X_25172_ clknet_leaf_55_clk _00061_ net8728 VGND VGND VPWR VPWR svm0.periodTop\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_22384_ _02386_ VGND VGND VPWR VPWR _02387_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24123_ _03893_ _03895_ _03984_ VGND VGND VPWR VPWR _03985_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_161_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21335_ net5626 net5674 VGND VGND VPWR VPWR _01349_ sky130_fd_sc_hd__nand2_4
Xwire4204 _06975_ VGND VGND VPWR VPWR net4204 sky130_fd_sc_hd__buf_1
Xwire4215 _06966_ VGND VGND VPWR VPWR net4215 sky130_fd_sc_hd__clkbuf_1
Xwire4226 net4227 VGND VGND VPWR VPWR net4226 sky130_fd_sc_hd__buf_1
X_24054_ _03915_ _03916_ VGND VGND VPWR VPWR _03917_ sky130_fd_sc_hd__nor2_1
X_21266_ _01279_ _01280_ VGND VGND VPWR VPWR _01281_ sky130_fd_sc_hd__xnor2_1
Xwire4248 net4249 VGND VGND VPWR VPWR net4248 sky130_fd_sc_hd__buf_1
Xwire4259 net4261 VGND VGND VPWR VPWR net4259 sky130_fd_sc_hd__buf_1
XFILLER_0_12_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3514 net3518 VGND VGND VPWR VPWR net3514 sky130_fd_sc_hd__clkbuf_1
X_23005_ _02871_ _02874_ VGND VGND VPWR VPWR _02875_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_25_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3525 _07063_ VGND VGND VPWR VPWR net3525 sky130_fd_sc_hd__buf_1
X_20217_ _12038_ cordic0.slte0.opB\[3\] net2937 VGND VGND VPWR VPWR _12039_ sky130_fd_sc_hd__mux2_1
Xwire3536 _07061_ VGND VGND VPWR VPWR net3536 sky130_fd_sc_hd__buf_1
X_21197_ _01166_ _01202_ _01206_ _01207_ _01212_ VGND VGND VPWR VPWR _01213_ sky130_fd_sc_hd__o221a_1
Xwire3547 net3548 VGND VGND VPWR VPWR net3547 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3558 _07039_ VGND VGND VPWR VPWR net3558 sky130_fd_sc_hd__buf_1
Xwire2813 net2814 VGND VGND VPWR VPWR net2813 sky130_fd_sc_hd__buf_1
Xwire2824 net2825 VGND VGND VPWR VPWR net2824 sky130_fd_sc_hd__buf_1
Xwire3569 net3570 VGND VGND VPWR VPWR net3569 sky130_fd_sc_hd__buf_1
X_20148_ _11947_ _11946_ _11941_ VGND VGND VPWR VPWR _11975_ sky130_fd_sc_hd__mux2_1
Xwire2835 _07041_ VGND VGND VPWR VPWR net2835 sky130_fd_sc_hd__clkbuf_1
Xwire2846 net2847 VGND VGND VPWR VPWR net2846 sky130_fd_sc_hd__clkbuf_2
Xwire2857 net2859 VGND VGND VPWR VPWR net2857 sky130_fd_sc_hd__buf_1
Xwire2868 net2870 VGND VGND VPWR VPWR net2868 sky130_fd_sc_hd__dlymetal6s2s_1
X_24956_ _04731_ VGND VGND VPWR VPWR _00759_ sky130_fd_sc_hd__clkbuf_1
X_12970_ _05168_ _05169_ net850 _05242_ VGND VGND VPWR VPWR _05243_ sky130_fd_sc_hd__a211oi_1
X_20079_ _11906_ _11907_ VGND VGND VPWR VPWR _11908_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_188_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23907_ pid_q.curr_int\[5\] VGND VGND VPWR VPWR _03771_ sky130_fd_sc_hd__inv_2
X_24887_ _04682_ net4570 net1997 VGND VGND VPWR VPWR _04683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14640_ net7437 net7182 net2878 VGND VGND VPWR VPWR _06804_ sky130_fd_sc_hd__and3_1
X_23838_ net5121 net5095 VGND VGND VPWR VPWR _03703_ sky130_fd_sc_hd__nor2_1
Xmax_length6830 net6828 VGND VGND VPWR VPWR net6830 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_71_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14571_ _06733_ _06747_ VGND VGND VPWR VPWR _06748_ sky130_fd_sc_hd__nor2_1
X_23769_ net1661 _03633_ VGND VGND VPWR VPWR _03635_ sky130_fd_sc_hd__or2_1
XFILLER_0_196_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_52_clk clknet_4_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_16
X_16310_ _08297_ _08299_ _08372_ VGND VGND VPWR VPWR _08373_ sky130_fd_sc_hd__o21a_1
X_13522_ net7866 net2946 net1938 VGND VGND VPWR VPWR _05793_ sky130_fd_sc_hd__and3_1
X_25508_ clknet_leaf_39_clk _00388_ net8754 VGND VGND VPWR VPWR svm0.delta\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17290_ net9199 net1924 net1462 VGND VGND VPWR VPWR _00374_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16241_ matmul0.matmul_stage_inst.mult1\[9\] net305 net2681 VGND VGND VPWR VPWR _08306_
+ sky130_fd_sc_hd__mux2_1
X_13453_ _05590_ net844 net845 VGND VGND VPWR VPWR _05726_ sky130_fd_sc_hd__a21o_1
X_25439_ clknet_leaf_91_clk _00322_ net8426 VGND VGND VPWR VPWR matmul0.sin\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_153_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16172_ _08237_ VGND VGND VPWR VPWR _00223_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_149_Left_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13384_ _05486_ _05558_ VGND VGND VPWR VPWR _05657_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6140 net6145 VGND VGND VPWR VPWR net6140 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15123_ _07191_ _07193_ _07196_ VGND VGND VPWR VPWR _07197_ sky130_fd_sc_hd__o21a_1
Xwire6162 net6163 VGND VGND VPWR VPWR net6162 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6173 net6169 VGND VGND VPWR VPWR net6173 sky130_fd_sc_hd__buf_1
Xfanout5388 net5392 VGND VGND VPWR VPWR net5388 sky130_fd_sc_hd__buf_1
XFILLER_0_121_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6184 net6182 VGND VGND VPWR VPWR net6184 sky130_fd_sc_hd__buf_1
Xwire5450 net5451 VGND VGND VPWR VPWR net5450 sky130_fd_sc_hd__clkbuf_1
Xwire6195 net6196 VGND VGND VPWR VPWR net6195 sky130_fd_sc_hd__buf_1
Xwire5461 net5462 VGND VGND VPWR VPWR net5461 sky130_fd_sc_hd__buf_1
X_19931_ _11761_ _11506_ net3856 net6049 _11762_ VGND VGND VPWR VPWR _11763_ sky130_fd_sc_hd__a221o_1
X_15054_ _07126_ _07127_ VGND VGND VPWR VPWR _07128_ sky130_fd_sc_hd__or2_1
Xwire5472 net5473 VGND VGND VPWR VPWR net5472 sky130_fd_sc_hd__buf_1
Xwire5483 net5484 VGND VGND VPWR VPWR net5483 sky130_fd_sc_hd__buf_1
X_14005_ _06217_ _06269_ VGND VGND VPWR VPWR _06270_ sky130_fd_sc_hd__xnor2_1
Xwire5494 net5495 VGND VGND VPWR VPWR net5494 sky130_fd_sc_hd__buf_1
Xwire4760 net4759 VGND VGND VPWR VPWR net4760 sky130_fd_sc_hd__buf_1
X_19862_ net6041 net6010 net6031 VGND VGND VPWR VPWR _11695_ sky130_fd_sc_hd__o21ai_1
Xwire4782 net4783 VGND VGND VPWR VPWR net4782 sky130_fd_sc_hd__clkbuf_1
X_18813_ net6376 _10623_ _10656_ VGND VGND VPWR VPWR _10657_ sky130_fd_sc_hd__a21oi_1
X_19793_ net6032 _11624_ _11626_ net6067 VGND VGND VPWR VPWR _11627_ sky130_fd_sc_hd__o211a_1
X_18744_ net6781 net2125 VGND VGND VPWR VPWR _10589_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_158_Left_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15956_ _07963_ _07964_ _07965_ VGND VGND VPWR VPWR _08024_ sky130_fd_sc_hd__o21a_1
X_14907_ net4206 net4202 net4210 net4208 VGND VGND VPWR VPWR _06981_ sky130_fd_sc_hd__o22a_1
X_15887_ _07951_ _07955_ VGND VGND VPWR VPWR _07956_ sky130_fd_sc_hd__xor2_1
X_18675_ net6893 net2131 net3231 VGND VGND VPWR VPWR _10521_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17626_ svm0.tB\[7\] _09477_ net4006 VGND VGND VPWR VPWR _09507_ sky130_fd_sc_hd__a21o_1
XFILLER_0_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14838_ matmul0.a\[8\] matmul0.matmul_stage_inst.e\[8\] _06928_ VGND VGND VPWR VPWR
+ _06936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_187_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17557_ net3278 svm0.tC\[10\] VGND VGND VPWR VPWR _09439_ sky130_fd_sc_hd__and2_1
X_14769_ net7448 _06895_ _06896_ net7459 net3621 VGND VGND VPWR VPWR _06897_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_43_clk clknet_4_15__leaf_clk VGND VGND VPWR VPWR clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16508_ net2638 _08565_ _08566_ _08563_ VGND VGND VPWR VPWR _08568_ sky130_fd_sc_hd__a31oi_1
X_17488_ _09299_ _09372_ _09377_ VGND VGND VPWR VPWR _09378_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19227_ net6139 net3175 VGND VGND VPWR VPWR _11064_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_167_Left_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16439_ _08466_ _08474_ _08440_ VGND VGND VPWR VPWR _08500_ sky130_fd_sc_hd__a21o_1
XFILLER_0_171_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19158_ net6069 VGND VGND VPWR VPWR _10995_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18109_ _09951_ _09959_ VGND VGND VPWR VPWR _09960_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_169_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19089_ net3896 net3192 net3202 VGND VGND VPWR VPWR _10926_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21120_ net5603 _01054_ _01134_ _01135_ VGND VGND VPWR VPWR _01136_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21051_ _01033_ _01034_ _01032_ VGND VGND VPWR VPWR _01067_ sky130_fd_sc_hd__o21a_1
Xwire2109 _10956_ VGND VGND VPWR VPWR net2109 sky130_fd_sc_hd__buf_1
X_20002_ _11824_ _11832_ VGND VGND VPWR VPWR _11833_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_176_Left_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1408 _11770_ VGND VGND VPWR VPWR net1408 sky130_fd_sc_hd__buf_1
Xwire1419 _11340_ VGND VGND VPWR VPWR net1419 sky130_fd_sc_hd__buf_1
X_24810_ net7955 _04628_ VGND VGND VPWR VPWR _04633_ sky130_fd_sc_hd__or2_1
XFILLER_0_185_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25790_ clknet_leaf_64_clk _00663_ net8668 VGND VGND VPWR VPWR matmul0.beta_pass\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24741_ _04570_ _04571_ _04572_ VGND VGND VPWR VPWR _04573_ sky130_fd_sc_hd__o21a_1
XFILLER_0_154_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21953_ net2474 _01854_ _01960_ VGND VGND VPWR VPWR _01961_ sky130_fd_sc_hd__o21ai_1
X_20904_ net5906 _00896_ _00919_ VGND VGND VPWR VPWR _00920_ sky130_fd_sc_hd__a21o_1
X_24672_ net9123 net1376 _04518_ VGND VGND VPWR VPWR _00688_ sky130_fd_sc_hd__a21o_1
X_21884_ _01892_ VGND VGND VPWR VPWR _01893_ sky130_fd_sc_hd__inv_2
X_23623_ net4636 net4922 VGND VGND VPWR VPWR _03490_ sky130_fd_sc_hd__nand2_1
XFILLER_0_166_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20835_ net5687 net5637 VGND VGND VPWR VPWR _00851_ sky130_fd_sc_hd__nand2_1
XFILLER_0_194_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23554_ _03410_ _03421_ VGND VGND VPWR VPWR _03422_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_185_Left_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length4713 net4714 VGND VGND VPWR VPWR net4713 sky130_fd_sc_hd__clkbuf_1
X_20766_ net5612 net5776 VGND VGND VPWR VPWR _12537_ sky130_fd_sc_hd__nand2_1
X_22505_ _02447_ _02504_ _02500_ VGND VGND VPWR VPWR _02506_ sky130_fd_sc_hd__a21o_1
Xwire705 net706 VGND VGND VPWR VPWR net705 sky130_fd_sc_hd__clkbuf_1
X_23485_ _03350_ _03353_ VGND VGND VPWR VPWR _03354_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire716 net717 VGND VGND VPWR VPWR net716 sky130_fd_sc_hd__buf_1
Xwire727 _05982_ VGND VGND VPWR VPWR net727 sky130_fd_sc_hd__buf_1
X_20697_ _12466_ _12467_ net3132 VGND VGND VPWR VPWR _12471_ sky130_fd_sc_hd__a21o_1
Xwire738 _04576_ VGND VGND VPWR VPWR net738 sky130_fd_sc_hd__buf_1
X_25224_ clknet_leaf_59_clk _00113_ net8693 VGND VGND VPWR VPWR svm0.vC\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire749 net750 VGND VGND VPWR VPWR net749 sky130_fd_sc_hd__buf_1
X_22436_ _02429_ _02437_ VGND VGND VPWR VPWR _02438_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25155_ clknet_leaf_44_clk _00044_ net8781 VGND VGND VPWR VPWR pid_q.target\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_161_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22367_ _02367_ _02369_ VGND VGND VPWR VPWR _02370_ sky130_fd_sc_hd__xor2_1
XFILLER_0_33_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24106_ _03964_ _03967_ VGND VGND VPWR VPWR _03968_ sky130_fd_sc_hd__xnor2_2
Xwire4012 net4013 VGND VGND VPWR VPWR net4012 sky130_fd_sc_hd__buf_1
XFILLER_0_103_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21318_ pid_d.prev_error\[0\] net5973 _01332_ VGND VGND VPWR VPWR _01333_ sky130_fd_sc_hd__and3_1
Xwire4023 _09230_ VGND VGND VPWR VPWR net4023 sky130_fd_sc_hd__buf_1
X_25086_ net5174 _04824_ _04830_ VGND VGND VPWR VPWR _04831_ sky130_fd_sc_hd__o21a_1
Xwire4034 _09196_ VGND VGND VPWR VPWR net4034 sky130_fd_sc_hd__clkbuf_1
X_22298_ _02299_ net2471 VGND VGND VPWR VPWR _02302_ sky130_fd_sc_hd__xnor2_2
Xwire3300 net3301 VGND VGND VPWR VPWR net3300 sky130_fd_sc_hd__clkbuf_1
Xwire4056 _08848_ VGND VGND VPWR VPWR net4056 sky130_fd_sc_hd__clkbuf_1
X_24037_ net4626 net4834 VGND VGND VPWR VPWR _03900_ sky130_fd_sc_hd__nand2_1
Xwire3322 net3323 VGND VGND VPWR VPWR net3322 sky130_fd_sc_hd__buf_1
Xwire4067 _08644_ VGND VGND VPWR VPWR net4067 sky130_fd_sc_hd__buf_1
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21249_ net5962 net5399 VGND VGND VPWR VPWR _01264_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_194_Left_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4078 _07573_ VGND VGND VPWR VPWR net4078 sky130_fd_sc_hd__clkbuf_1
Xwire3344 _08927_ VGND VGND VPWR VPWR net3344 sky130_fd_sc_hd__clkbuf_1
Xwire4089 net4090 VGND VGND VPWR VPWR net4089 sky130_fd_sc_hd__buf_1
Xwire3355 net3356 VGND VGND VPWR VPWR net3355 sky130_fd_sc_hd__buf_1
Xwire2621 net2622 VGND VGND VPWR VPWR net2621 sky130_fd_sc_hd__clkbuf_2
Xwire2632 net2633 VGND VGND VPWR VPWR net2632 sky130_fd_sc_hd__buf_1
Xwire3388 _08647_ VGND VGND VPWR VPWR net3388 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2654 net2655 VGND VGND VPWR VPWR net2654 sky130_fd_sc_hd__buf_1
Xwire3399 net3400 VGND VGND VPWR VPWR net3399 sky130_fd_sc_hd__buf_1
X_15810_ _07768_ net1530 net1535 VGND VGND VPWR VPWR _07880_ sky130_fd_sc_hd__o21ai_1
Xwire1920 net1921 VGND VGND VPWR VPWR net1920 sky130_fd_sc_hd__clkbuf_1
Xwire2665 _07715_ VGND VGND VPWR VPWR net2665 sky130_fd_sc_hd__buf_1
Xwire1931 net1932 VGND VGND VPWR VPWR net1931 sky130_fd_sc_hd__buf_1
Xwire2676 _07670_ VGND VGND VPWR VPWR net2676 sky130_fd_sc_hd__buf_1
X_16790_ net7581 matmul0.a\[14\] net3373 VGND VGND VPWR VPWR _08785_ sky130_fd_sc_hd__mux2_1
Xwire1942 net1943 VGND VGND VPWR VPWR net1942 sky130_fd_sc_hd__buf_1
Xwire2687 net2688 VGND VGND VPWR VPWR net2687 sky130_fd_sc_hd__clkbuf_1
Xwire1953 net1954 VGND VGND VPWR VPWR net1953 sky130_fd_sc_hd__buf_1
X_15741_ net1529 net1850 VGND VGND VPWR VPWR _07812_ sky130_fd_sc_hd__xnor2_1
X_24939_ net8867 net145 VGND VGND VPWR VPWR _04720_ sky130_fd_sc_hd__and2b_1
XFILLER_0_172_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1975 net1976 VGND VGND VPWR VPWR net1975 sky130_fd_sc_hd__buf_1
X_12953_ net789 _05031_ VGND VGND VPWR VPWR _05226_ sky130_fd_sc_hd__xnor2_1
Xwire1986 _04905_ VGND VGND VPWR VPWR net1986 sky130_fd_sc_hd__buf_1
Xmax_length8040 pid_q.target\[0\] VGND VGND VPWR VPWR net8040 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18460_ net3925 net3225 VGND VGND VPWR VPWR _10310_ sky130_fd_sc_hd__nor2_1
X_15672_ _07696_ _07701_ VGND VGND VPWR VPWR _07743_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12884_ net7823 _04962_ net2971 VGND VGND VPWR VPWR _05157_ sky130_fd_sc_hd__and3_1
Xmax_length8073 net8074 VGND VGND VPWR VPWR net8073 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17411_ _09311_ net615 _09312_ _09314_ VGND VGND VPWR VPWR _00385_ sky130_fd_sc_hd__a31o_1
Xmax_length7361 net7362 VGND VGND VPWR VPWR net7361 sky130_fd_sc_hd__buf_1
X_14623_ net6456 _06785_ VGND VGND VPWR VPWR _06793_ sky130_fd_sc_hd__nand2_1
X_18391_ _10041_ _10241_ VGND VGND VPWR VPWR _10242_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length7383 matmul0.matmul_stage_inst.f\[10\] VGND VGND VPWR VPWR net7383 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_25_clk clknet_4_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_28_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17342_ net6691 _09214_ _09218_ _09220_ _09255_ VGND VGND VPWR VPWR _09256_ sky130_fd_sc_hd__a311o_1
Xmax_length6671 net6663 VGND VGND VPWR VPWR net6671 sky130_fd_sc_hd__clkbuf_1
X_14554_ net7257 net5223 VGND VGND VPWR VPWR _06732_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length6693 net6690 VGND VGND VPWR VPWR net6693 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13505_ _05777_ VGND VGND VPWR VPWR _00411_ sky130_fd_sc_hd__clkbuf_1
X_17273_ _09191_ net187 net1798 net8971 VGND VGND VPWR VPWR _00367_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14485_ _06668_ _06669_ VGND VGND VPWR VPWR _06670_ sky130_fd_sc_hd__xnor2_1
Xmax_length5992 net5993 VGND VGND VPWR VPWR net5992 sky130_fd_sc_hd__buf_1
XFILLER_0_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19012_ net6114 net6155 VGND VGND VPWR VPWR _10849_ sky130_fd_sc_hd__xnor2_1
X_16224_ net979 _08288_ VGND VGND VPWR VPWR _08289_ sky130_fd_sc_hd__xnor2_1
X_13436_ net4255 VGND VGND VPWR VPWR _05709_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16155_ net1088 net1511 VGND VGND VPWR VPWR _08221_ sky130_fd_sc_hd__xor2_1
X_13367_ _05528_ _05534_ _05639_ VGND VGND VPWR VPWR _05640_ sky130_fd_sc_hd__o21a_1
XFILLER_0_134_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15106_ _07177_ _07178_ _07129_ net3464 VGND VGND VPWR VPWR _07180_ sky130_fd_sc_hd__o211a_1
X_16086_ _08064_ _08151_ _08152_ VGND VGND VPWR VPWR _08153_ sky130_fd_sc_hd__a21o_1
X_13298_ _05570_ VGND VGND VPWR VPWR _05571_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5280 net5281 VGND VGND VPWR VPWR net5280 sky130_fd_sc_hd__clkbuf_1
Xwire5291 net5292 VGND VGND VPWR VPWR net5291 sky130_fd_sc_hd__clkbuf_1
X_19914_ _11329_ VGND VGND VPWR VPWR _11746_ sky130_fd_sc_hd__inv_2
X_15037_ _07109_ _07110_ VGND VGND VPWR VPWR _07111_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_43_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4590 net4591 VGND VGND VPWR VPWR net4590 sky130_fd_sc_hd__dlymetal6s2s_1
X_19845_ net2506 net6130 net6157 VGND VGND VPWR VPWR _11678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19776_ _11609_ _11555_ _11558_ VGND VGND VPWR VPWR _11611_ sky130_fd_sc_hd__nand3_1
X_16988_ _08946_ _08947_ _08948_ net4049 _08825_ net4059 VGND VGND VPWR VPWR _08950_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_147_Right_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18727_ _10570_ net1430 _10571_ VGND VGND VPWR VPWR _10572_ sky130_fd_sc_hd__o21a_1
X_15939_ _08003_ _08006_ VGND VGND VPWR VPWR _08008_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18658_ _10504_ VGND VGND VPWR VPWR _10505_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_189_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17609_ net6747 VGND VGND VPWR VPWR _09490_ sky130_fd_sc_hd__inv_2
XFILLER_0_149_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18589_ net6792 _10436_ _10372_ VGND VGND VPWR VPWR _10437_ sky130_fd_sc_hd__o21a_1
XFILLER_0_188_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_16_clk clknet_4_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20620_ _12399_ _12391_ net707 VGND VGND VPWR VPWR _12401_ sky130_fd_sc_hd__or3_1
XFILLER_0_80_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20551_ _12334_ _12335_ net1053 _12320_ VGND VGND VPWR VPWR _12336_ sky130_fd_sc_hd__o211ai_2
Xmax_length3308 net3309 VGND VGND VPWR VPWR net3308 sky130_fd_sc_hd__buf_1
XFILLER_0_11_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6909 net6910 VGND VGND VPWR VPWR net6909 sky130_fd_sc_hd__buf_1
X_23270_ _03130_ _03139_ VGND VGND VPWR VPWR _03140_ sky130_fd_sc_hd__nand2_1
X_20482_ _12268_ _12270_ net6461 VGND VGND VPWR VPWR _12271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22221_ net5800 net3786 net5780 VGND VGND VPWR VPWR _02226_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22152_ net1168 _02157_ VGND VGND VPWR VPWR _02158_ sky130_fd_sc_hd__xnor2_1
X_21103_ net5607 net5911 VGND VGND VPWR VPWR _01119_ sky130_fd_sc_hd__nand2_2
XFILLER_0_121_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22083_ _02084_ _02089_ VGND VGND VPWR VPWR _02090_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25911_ clknet_leaf_29_clk _00784_ net8654 VGND VGND VPWR VPWR pid_q.out\[7\] sky130_fd_sc_hd__dfrtp_1
X_21034_ _01049_ net3836 net5775 net5635 VGND VGND VPWR VPWR _01050_ sky130_fd_sc_hd__o211a_1
Xwire1205 net1206 VGND VGND VPWR VPWR net1205 sky130_fd_sc_hd__buf_1
Xwire1216 net1219 VGND VGND VPWR VPWR net1216 sky130_fd_sc_hd__buf_1
X_25842_ clknet_leaf_20_clk _00715_ net8743 VGND VGND VPWR VPWR pid_q.mult0.b\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1238 net1239 VGND VGND VPWR VPWR net1238 sky130_fd_sc_hd__clkbuf_1
Xwire1249 _08331_ VGND VGND VPWR VPWR net1249 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_114_Right_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25773_ clknet_leaf_24_clk _00646_ net8583 VGND VGND VPWR VPWR pid_d.out\[14\] sky130_fd_sc_hd__dfrtp_2
X_22985_ _02860_ VGND VGND VPWR VPWR _00659_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24724_ _04556_ _04557_ net5273 VGND VGND VPWR VPWR _04558_ sky130_fd_sc_hd__a21oi_1
X_21936_ net5763 net5432 VGND VGND VPWR VPWR _01944_ sky130_fd_sc_hd__nand2_1
XFILLER_0_167_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24655_ net7477 net8874 net2146 VGND VGND VPWR VPWR _04509_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_167_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21867_ _01860_ _01875_ VGND VGND VPWR VPWR _01876_ sky130_fd_sc_hd__xnor2_2
Xfanout8717 net8722 VGND VGND VPWR VPWR net8717 sky130_fd_sc_hd__buf_1
XFILLER_0_37_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23606_ net696 _03473_ VGND VGND VPWR VPWR _03474_ sky130_fd_sc_hd__xor2_1
Xmax_length5222 net5223 VGND VGND VPWR VPWR net5222 sky130_fd_sc_hd__buf_1
Xwire8801 net8802 VGND VGND VPWR VPWR net8801 sky130_fd_sc_hd__buf_1
XFILLER_0_167_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20818_ _12513_ _12518_ _00833_ VGND VGND VPWR VPWR _00834_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_182_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24586_ _04368_ _04370_ _04366_ VGND VGND VPWR VPWR _04442_ sky130_fd_sc_hd__o21ba_1
Xwire8812 net8813 VGND VGND VPWR VPWR net8812 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21798_ _01649_ _01725_ _01724_ VGND VGND VPWR VPWR _01808_ sky130_fd_sc_hd__a21oi_1
Xwire8823 net8824 VGND VGND VPWR VPWR net8823 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8834 net8835 VGND VGND VPWR VPWR net8834 sky130_fd_sc_hd__buf_1
XFILLER_0_166_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23537_ _03399_ _03404_ VGND VGND VPWR VPWR _03405_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length5277 net5278 VGND VGND VPWR VPWR net5277 sky130_fd_sc_hd__clkbuf_1
Xwire8845 net8846 VGND VGND VPWR VPWR net8845 sky130_fd_sc_hd__clkbuf_1
Xwire8856 net8857 VGND VGND VPWR VPWR net8856 sky130_fd_sc_hd__buf_1
XFILLER_0_181_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20749_ _12508_ _12519_ VGND VGND VPWR VPWR _12520_ sky130_fd_sc_hd__xnor2_2
Xwire502 _07559_ VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8867 net8868 VGND VGND VPWR VPWR net8867 sky130_fd_sc_hd__buf_1
Xwire513 net514 VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__clkbuf_1
Xwire8878 net8879 VGND VGND VPWR VPWR net8878 sky130_fd_sc_hd__clkbuf_1
Xwire524 net525 VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__buf_1
X_14270_ net63 net2931 net2278 net9103 VGND VGND VPWR VPWR _00043_ sky130_fd_sc_hd__a22o_1
Xwire8889 net8887 VGND VGND VPWR VPWR net8889 sky130_fd_sc_hd__buf_1
Xwire535 _05240_ VGND VGND VPWR VPWR net535 sky130_fd_sc_hd__clkbuf_1
X_23468_ net4662 net4944 VGND VGND VPWR VPWR _03337_ sky130_fd_sc_hd__nand2_2
Xwire546 net547 VGND VGND VPWR VPWR net546 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire557 net558 VGND VGND VPWR VPWR net557 sky130_fd_sc_hd__clkbuf_1
X_13221_ _05459_ _05492_ _05493_ VGND VGND VPWR VPWR _05494_ sky130_fd_sc_hd__a21o_1
X_25207_ clknet_leaf_62_clk _00096_ net8666 VGND VGND VPWR VPWR matmul0.b_in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire568 net569 VGND VGND VPWR VPWR net568 sky130_fd_sc_hd__buf_1
Xwire579 net580 VGND VGND VPWR VPWR net579 sky130_fd_sc_hd__clkbuf_1
X_22419_ net5691 net5390 VGND VGND VPWR VPWR _02421_ sky130_fd_sc_hd__nand2_1
X_23399_ _03265_ _03268_ VGND VGND VPWR VPWR _03269_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25138_ clknet_4_14__leaf_clk _00027_ net8832 VGND VGND VPWR VPWR svm0.tC\[10\] sky130_fd_sc_hd__dfrtp_1
X_13152_ _05417_ _05418_ _05423_ VGND VGND VPWR VPWR _05425_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13083_ _05342_ _05355_ VGND VGND VPWR VPWR _05356_ sky130_fd_sc_hd__xnor2_1
X_25069_ net3734 _04811_ net4424 VGND VGND VPWR VPWR _04816_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_27_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17960_ net7141 _09810_ VGND VGND VPWR VPWR _09811_ sky130_fd_sc_hd__xnor2_1
Xwire3141 net3142 VGND VGND VPWR VPWR net3141 sky130_fd_sc_hd__buf_1
X_16911_ net6404 cordic0.slte0.opA\[9\] VGND VGND VPWR VPWR _08875_ sky130_fd_sc_hd__xor2_1
Xwire3152 net3153 VGND VGND VPWR VPWR net3152 sky130_fd_sc_hd__buf_1
XFILLER_0_109_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3163 net3164 VGND VGND VPWR VPWR net3163 sky130_fd_sc_hd__clkbuf_1
X_17891_ net7027 net3970 _09740_ _09741_ _09682_ VGND VGND VPWR VPWR _09742_ sky130_fd_sc_hd__a221o_1
Xwire3174 net3175 VGND VGND VPWR VPWR net3174 sky130_fd_sc_hd__buf_1
Xwire2440 net2441 VGND VGND VPWR VPWR net2440 sky130_fd_sc_hd__buf_1
Xwire3185 net3186 VGND VGND VPWR VPWR net3185 sky130_fd_sc_hd__clkbuf_2
Xwire2451 net2452 VGND VGND VPWR VPWR net2451 sky130_fd_sc_hd__buf_1
X_19630_ _11465_ _11466_ VGND VGND VPWR VPWR _11467_ sky130_fd_sc_hd__xnor2_1
Xwire2462 _02520_ VGND VGND VPWR VPWR net2462 sky130_fd_sc_hd__clkbuf_1
X_16842_ cordic0.sin\[9\] matmul0.sin\[9\] net3366 VGND VGND VPWR VPWR _08812_ sky130_fd_sc_hd__mux2_1
Xwire2473 _02225_ VGND VGND VPWR VPWR net2473 sky130_fd_sc_hd__buf_1
XFILLER_0_18_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2484 _00809_ VGND VGND VPWR VPWR net2484 sky130_fd_sc_hd__buf_1
XFILLER_0_176_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1750 _11464_ VGND VGND VPWR VPWR net1750 sky130_fd_sc_hd__clkbuf_1
Xwire2495 net2496 VGND VGND VPWR VPWR net2495 sky130_fd_sc_hd__clkbuf_1
X_19561_ net6252 _11393_ _11396_ _11397_ VGND VGND VPWR VPWR _11398_ sky130_fd_sc_hd__and4_1
Xwire1761 _10540_ VGND VGND VPWR VPWR net1761 sky130_fd_sc_hd__clkbuf_1
X_13985_ _06201_ _06198_ net906 VGND VGND VPWR VPWR _06250_ sky130_fd_sc_hd__a21bo_1
X_16773_ matmul0.a_in\[6\] matmul0.a\[6\] _08770_ VGND VGND VPWR VPWR _08776_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1783 _09597_ VGND VGND VPWR VPWR net1783 sky130_fd_sc_hd__clkbuf_1
Xwire1794 _09438_ VGND VGND VPWR VPWR net1794 sky130_fd_sc_hd__clkbuf_1
X_18512_ net7076 _10304_ _10359_ _10360_ net6970 VGND VGND VPWR VPWR _10361_ sky130_fd_sc_hd__o2111a_1
X_12936_ net790 _05208_ VGND VGND VPWR VPWR _05209_ sky130_fd_sc_hd__xnor2_1
X_15724_ net1851 net1537 _07674_ VGND VGND VPWR VPWR _07795_ sky130_fd_sc_hd__o21a_1
X_19492_ net6128 net6116 VGND VGND VPWR VPWR _11329_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_87_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18443_ _10041_ _10292_ _10241_ VGND VGND VPWR VPWR _10293_ sky130_fd_sc_hd__a21o_1
X_12867_ net1007 net1594 _05139_ VGND VGND VPWR VPWR _05140_ sky130_fd_sc_hd__o21ai_1
X_15655_ net2776 net2666 _07718_ _07719_ _07726_ VGND VGND VPWR VPWR _07727_ sky130_fd_sc_hd__a32o_1
Xmax_length7180 matmul0.cos\[4\] VGND VGND VPWR VPWR net7180 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length7191 matmul0.b\[1\] VGND VGND VPWR VPWR net7191 sky130_fd_sc_hd__clkbuf_1
X_14606_ _06778_ VGND VGND VPWR VPWR _06779_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15586_ net3398 _07657_ VGND VGND VPWR VPWR _07658_ sky130_fd_sc_hd__xnor2_2
X_18374_ _10223_ _10224_ VGND VGND VPWR VPWR _10225_ sky130_fd_sc_hd__xor2_1
X_12798_ _05067_ _05070_ VGND VGND VPWR VPWR _05071_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17325_ _09236_ _09237_ _09238_ net4032 VGND VGND VPWR VPWR _09239_ sky130_fd_sc_hd__a22o_1
X_14537_ net5247 _06710_ _06715_ VGND VGND VPWR VPWR _06716_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17256_ net2959 net158 net2162 net9141 VGND VGND VPWR VPWR _00354_ sky130_fd_sc_hd__a22o_1
X_14468_ net7364 net5311 VGND VGND VPWR VPWR _06656_ sky130_fd_sc_hd__xor2_1
XFILLER_0_154_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13419_ net7921 net1317 _05690_ _05691_ VGND VGND VPWR VPWR _05692_ sky130_fd_sc_hd__a31o_1
X_16207_ net2746 net3435 VGND VGND VPWR VPWR _08272_ sky130_fd_sc_hd__nor2_1
XFILLER_0_180_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17187_ net617 _09137_ VGND VGND VPWR VPWR _09138_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_144_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14399_ _06602_ VGND VGND VPWR VPWR _00085_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16138_ _08120_ _08125_ _08203_ VGND VGND VPWR VPWR _08204_ sky130_fd_sc_hd__o21a_1
X_16069_ _08050_ net1258 _08132_ _08133_ _08135_ VGND VGND VPWR VPWR _08136_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_5_clk clknet_4_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_166_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19828_ _11606_ _11608_ VGND VGND VPWR VPWR _11662_ sky130_fd_sc_hd__and2b_1
XFILLER_0_166_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19759_ _11580_ _11593_ VGND VGND VPWR VPWR _11594_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_190_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22770_ _02691_ VGND VGND VPWR VPWR _00613_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21721_ _01730_ _01731_ VGND VGND VPWR VPWR _01732_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24440_ net4515 _04289_ _04295_ _04297_ VGND VGND VPWR VPWR _04298_ sky130_fd_sc_hd__o211a_1
X_21652_ net5593 net5680 VGND VGND VPWR VPWR _01663_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8108 net8109 VGND VGND VPWR VPWR net8108 sky130_fd_sc_hd__buf_1
XFILLER_0_93_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8119 net7 VGND VGND VPWR VPWR net8119 sky130_fd_sc_hd__buf_1
XFILLER_0_75_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20603_ net3163 _12375_ _12383_ VGND VGND VPWR VPWR _12384_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24371_ net4554 net4581 net3053 VGND VGND VPWR VPWR _04230_ sky130_fd_sc_hd__and3_1
XFILLER_0_163_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21583_ _01589_ _01594_ VGND VGND VPWR VPWR _01595_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3105 _02519_ VGND VGND VPWR VPWR net3105 sky130_fd_sc_hd__buf_1
Xwire7418 net7419 VGND VGND VPWR VPWR net7418 sky130_fd_sc_hd__clkbuf_1
Xwire7429 net7430 VGND VGND VPWR VPWR net7429 sky130_fd_sc_hd__clkbuf_1
X_23322_ net4887 net4880 net4760 net4771 VGND VGND VPWR VPWR _03192_ sky130_fd_sc_hd__and4_1
XFILLER_0_145_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6706 net6707 VGND VGND VPWR VPWR net6706 sky130_fd_sc_hd__buf_1
X_20534_ _12311_ _12319_ VGND VGND VPWR VPWR _12320_ sky130_fd_sc_hd__xnor2_1
Xmax_length3149 net3150 VGND VGND VPWR VPWR net3149 sky130_fd_sc_hd__buf_1
XFILLER_0_7_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6728 svm0.counter\[5\] VGND VGND VPWR VPWR net6728 sky130_fd_sc_hd__buf_1
Xwire6739 net6740 VGND VGND VPWR VPWR net6739 sky130_fd_sc_hd__buf_1
X_23253_ _03116_ _03119_ VGND VGND VPWR VPWR _03123_ sky130_fd_sc_hd__xor2_2
X_20465_ cordic0.slte0.opA\[15\] _12249_ VGND VGND VPWR VPWR _12256_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22204_ _02122_ _02124_ _02208_ VGND VGND VPWR VPWR _02209_ sky130_fd_sc_hd__a21oi_1
X_23184_ net5040 net4777 VGND VGND VPWR VPWR _03054_ sky130_fd_sc_hd__nand2_1
X_20396_ _12192_ _12193_ net3313 VGND VGND VPWR VPWR _12194_ sky130_fd_sc_hd__a21o_1
X_22135_ _02031_ _02032_ _02140_ VGND VGND VPWR VPWR _02141_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_11_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22066_ net1045 net1170 _02071_ _02072_ VGND VGND VPWR VPWR _02073_ sky130_fd_sc_hd__o211a_1
Xwire1002 _05230_ VGND VGND VPWR VPWR net1002 sky130_fd_sc_hd__clkbuf_1
X_21017_ net5528 net5950 VGND VGND VPWR VPWR _01033_ sky130_fd_sc_hd__nand2_1
Xwire1013 net1014 VGND VGND VPWR VPWR net1013 sky130_fd_sc_hd__clkbuf_2
Xwire1024 net1025 VGND VGND VPWR VPWR net1024 sky130_fd_sc_hd__buf_1
Xwire1035 _02235_ VGND VGND VPWR VPWR net1035 sky130_fd_sc_hd__clkbuf_1
Xwire1046 _01890_ VGND VGND VPWR VPWR net1046 sky130_fd_sc_hd__buf_1
X_25825_ clknet_leaf_37_clk _00698_ net8744 VGND VGND VPWR VPWR pid_q.curr_error\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1057 _11540_ VGND VGND VPWR VPWR net1057 sky130_fd_sc_hd__buf_1
XFILLER_0_96_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1068 _10529_ VGND VGND VPWR VPWR net1068 sky130_fd_sc_hd__clkbuf_1
Xwire1079 net1080 VGND VGND VPWR VPWR net1079 sky130_fd_sc_hd__clkbuf_2
X_13770_ _06036_ _06037_ VGND VGND VPWR VPWR _06038_ sky130_fd_sc_hd__xnor2_1
X_25756_ clknet_leaf_13_clk _00629_ net8606 VGND VGND VPWR VPWR pid_d.kp\[14\] sky130_fd_sc_hd__dfrtp_1
X_22968_ matmul0.beta_pass\[3\] net2202 net6567 VGND VGND VPWR VPWR _02852_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12721_ _04984_ _04989_ _04993_ VGND VGND VPWR VPWR _04994_ sky130_fd_sc_hd__a21oi_4
X_24707_ net1642 VGND VGND VPWR VPWR _04543_ sky130_fd_sc_hd__buf_1
X_21919_ _01832_ _01834_ _01926_ VGND VGND VPWR VPWR _01927_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_139_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25687_ clknet_leaf_2_clk _00560_ net8572 VGND VGND VPWR VPWR pid_d.curr_error\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_179_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22899_ _02792_ VGND VGND VPWR VPWR _00641_ sky130_fd_sc_hd__clkbuf_1
X_15440_ net6631 matmul0.matmul_stage_inst.d\[13\] matmul0.matmul_stage_inst.c\[13\]
+ net6533 VGND VGND VPWR VPWR _07514_ sky130_fd_sc_hd__a22o_1
X_24638_ _04421_ _04414_ VGND VGND VPWR VPWR _04493_ sky130_fd_sc_hd__or2b_1
X_12652_ net5304 _04892_ net3694 net2990 svm0.vC\[1\] VGND VGND VPWR VPWR _04925_
+ sky130_fd_sc_hd__a32oi_1
XFILLER_0_183_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout8569 net8575 VGND VGND VPWR VPWR net8569 sky130_fd_sc_hd__dlymetal6s2s_1
X_15371_ net2704 _07444_ _07224_ net3445 VGND VGND VPWR VPWR _07445_ sky130_fd_sc_hd__o211a_1
Xwire8631 net8632 VGND VGND VPWR VPWR net8631 sky130_fd_sc_hd__buf_1
X_24569_ net4514 net4807 VGND VGND VPWR VPWR _04425_ sky130_fd_sc_hd__nand2_1
X_12583_ net8863 net7496 VGND VGND VPWR VPWR _04868_ sky130_fd_sc_hd__and2_1
Xfanout7835 svm0.periodTop\[4\] VGND VGND VPWR VPWR net7835 sky130_fd_sc_hd__buf_1
Xwire8642 net8643 VGND VGND VPWR VPWR net8642 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17110_ net3307 _09066_ VGND VGND VPWR VPWR _09067_ sky130_fd_sc_hd__nor2_1
Xwire310 _08305_ VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__clkbuf_1
X_14322_ _06529_ matmul0.a_in\[0\] net904 VGND VGND VPWR VPWR _06544_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8675 net8673 VGND VGND VPWR VPWR net8675 sky130_fd_sc_hd__dlymetal6s2s_1
X_18090_ _09914_ _09923_ _09929_ VGND VGND VPWR VPWR _09941_ sky130_fd_sc_hd__a21oi_1
Xwire321 _06016_ VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__buf_1
XFILLER_0_163_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7941 net7934 VGND VGND VPWR VPWR net7941 sky130_fd_sc_hd__buf_1
XFILLER_0_37_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8686 net8684 VGND VGND VPWR VPWR net8686 sky130_fd_sc_hd__buf_1
Xwire332 net333 VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__clkbuf_1
Xwire7952 net7953 VGND VGND VPWR VPWR net7952 sky130_fd_sc_hd__clkbuf_1
Xwire8697 net8701 VGND VGND VPWR VPWR net8697 sky130_fd_sc_hd__clkbuf_1
Xwire343 net344 VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__buf_1
Xwire7963 net7964 VGND VGND VPWR VPWR net7963 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17041_ net2171 _09000_ VGND VGND VPWR VPWR _09001_ sky130_fd_sc_hd__xor2_1
XFILLER_0_20_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire354 net355 VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__buf_1
Xwire7974 net7975 VGND VGND VPWR VPWR net7974 sky130_fd_sc_hd__buf_1
XFILLER_0_29_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire365 _08086_ VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__clkbuf_1
X_14253_ net2284 VGND VGND VPWR VPWR _06508_ sky130_fd_sc_hd__buf_1
XFILLER_0_162_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7985 net7986 VGND VGND VPWR VPWR net7985 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire376 net377 VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__clkbuf_2
Xwire7996 net7997 VGND VGND VPWR VPWR net7996 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_150_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire387 net388 VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__clkbuf_1
X_13204_ net919 _05476_ VGND VGND VPWR VPWR _05477_ sky130_fd_sc_hd__and2_1
Xwire398 net399 VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14184_ net7602 net1121 VGND VGND VPWR VPWR _06444_ sky130_fd_sc_hd__nand2_1
Xmax_length2971 net2972 VGND VGND VPWR VPWR net2971 sky130_fd_sc_hd__buf_1
XFILLER_0_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2982 net2983 VGND VGND VPWR VPWR net2982 sky130_fd_sc_hd__buf_1
X_13135_ _05290_ _05296_ _05342_ net7936 VGND VGND VPWR VPWR _05408_ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18992_ _10828_ VGND VGND VPWR VPWR _10829_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_29_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13066_ net7908 net1948 VGND VGND VPWR VPWR _05339_ sky130_fd_sc_hd__nand2_1
X_17943_ net3240 _09793_ VGND VGND VPWR VPWR _09794_ sky130_fd_sc_hd__xnor2_1
X_17874_ _09723_ _09603_ _09724_ VGND VGND VPWR VPWR _09725_ sky130_fd_sc_hd__a21oi_1
Xwire2270 net2271 VGND VGND VPWR VPWR net2270 sky130_fd_sc_hd__clkbuf_1
Xwire2281 net2282 VGND VGND VPWR VPWR net2281 sky130_fd_sc_hd__buf_1
X_19613_ net2505 _11449_ VGND VGND VPWR VPWR _11450_ sky130_fd_sc_hd__xnor2_2
X_16825_ net4287 VGND VGND VPWR VPWR _08803_ sky130_fd_sc_hd__buf_1
Xwire2292 net2293 VGND VGND VPWR VPWR net2292 sky130_fd_sc_hd__buf_1
XFILLER_0_136_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire1591 _05293_ VGND VGND VPWR VPWR net1591 sky130_fd_sc_hd__buf_1
X_19544_ net6116 net6105 _11328_ VGND VGND VPWR VPWR _11381_ sky130_fd_sc_hd__a21o_1
Xmax_cap1 net9247 VGND VGND VPWR VPWR net9246 sky130_fd_sc_hd__clkbuf_1
X_16756_ net7556 matmul0.b\[14\] net3381 VGND VGND VPWR VPWR _08767_ sky130_fd_sc_hd__mux2_1
X_13968_ _06227_ _06232_ VGND VGND VPWR VPWR _06233_ sky130_fd_sc_hd__xnor2_1
X_15707_ net3458 net2766 VGND VGND VPWR VPWR _07778_ sky130_fd_sc_hd__nor2_1
X_12919_ net7933 net1949 VGND VGND VPWR VPWR _05192_ sky130_fd_sc_hd__nand2_1
X_19475_ _10984_ _11265_ _11311_ _11122_ VGND VGND VPWR VPWR _11312_ sky130_fd_sc_hd__a22o_1
X_13899_ _06128_ _06163_ _06164_ VGND VGND VPWR VPWR _06165_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_61_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16687_ _08716_ _08712_ _08717_ VGND VGND VPWR VPWR _08718_ sky130_fd_sc_hd__a21o_1
XFILLER_0_159_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18426_ _10275_ VGND VGND VPWR VPWR _10276_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_174_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15638_ _07667_ _07709_ VGND VGND VPWR VPWR _07710_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18357_ _10175_ net2543 VGND VGND VPWR VPWR _10208_ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15569_ _07641_ VGND VGND VPWR VPWR _00216_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_185_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17308_ net7765 net1795 net7742 VGND VGND VPWR VPWR _09222_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18288_ net963 _09834_ VGND VGND VPWR VPWR _10139_ sky130_fd_sc_hd__nand2_1
X_17239_ svm0.state\[1\] VGND VGND VPWR VPWR _09186_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20250_ _12064_ VGND VGND VPWR VPWR _00475_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20181_ _11974_ _11944_ VGND VGND VPWR VPWR _12007_ sky130_fd_sc_hd__or2b_1
XFILLER_0_177_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23940_ _03701_ _03698_ VGND VGND VPWR VPWR _03804_ sky130_fd_sc_hd__nand2_1
XFILLER_0_193_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23871_ net1164 _03637_ _03735_ VGND VGND VPWR VPWR _03736_ sky130_fd_sc_hd__a21o_1
XFILLER_0_193_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25610_ clknet_leaf_108_clk _00483_ net8350 VGND VGND VPWR VPWR cordic0.slte0.opA\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_22822_ net5366 net5984 VGND VGND VPWR VPWR _02724_ sky130_fd_sc_hd__xor2_1
Xmax_length7916 net7917 VGND VGND VPWR VPWR net7916 sky130_fd_sc_hd__buf_1
XFILLER_0_196_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25541_ clknet_leaf_33_clk _00421_ net8674 VGND VGND VPWR VPWR pid_q.prev_int\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_22753_ net4303 net8924 VGND VGND VPWR VPWR _02680_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21704_ net2069 _01713_ VGND VGND VPWR VPWR _01715_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25472_ clknet_leaf_48_clk _00352_ net8761 VGND VGND VPWR VPWR svm0.tB\[10\] sky130_fd_sc_hd__dfrtp_1
X_22684_ pid_d.ki\[5\] net2439 net2993 pid_d.kp\[5\] VGND VGND VPWR VPWR _02631_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24423_ net2020 net2404 _04280_ VGND VGND VPWR VPWR _04281_ sky130_fd_sc_hd__o21ai_1
X_21635_ _01644_ _01542_ _01645_ VGND VGND VPWR VPWR _01646_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire7204 net7205 VGND VGND VPWR VPWR net7204 sky130_fd_sc_hd__clkbuf_1
Xwire7215 net7216 VGND VGND VPWR VPWR net7215 sky130_fd_sc_hd__buf_1
XFILLER_0_35_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24354_ _04204_ _04212_ VGND VGND VPWR VPWR _04213_ sky130_fd_sc_hd__xnor2_2
Xwire7226 matmul0.alpha_pass\[12\] VGND VGND VPWR VPWR net7226 sky130_fd_sc_hd__clkbuf_1
X_21566_ _01455_ _01457_ _01456_ VGND VGND VPWR VPWR _01578_ sky130_fd_sc_hd__o21a_1
Xwire7237 net7238 VGND VGND VPWR VPWR net7237 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_35_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7248 matmul0.alpha_pass\[11\] VGND VGND VPWR VPWR net7248 sky130_fd_sc_hd__buf_1
XFILLER_0_151_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5718 net5734 VGND VGND VPWR VPWR net5718 sky130_fd_sc_hd__buf_1
XFILLER_0_16_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2201 _08818_ VGND VGND VPWR VPWR net2201 sky130_fd_sc_hd__clkbuf_1
X_23305_ net1031 VGND VGND VPWR VPWR _03175_ sky130_fd_sc_hd__inv_2
Xwire6525 net6526 VGND VGND VPWR VPWR net6525 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_63_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_112_Left_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20517_ net1053 _12303_ VGND VGND VPWR VPWR _12304_ sky130_fd_sc_hd__or2_1
Xmax_length2223 net2224 VGND VGND VPWR VPWR net2223 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24285_ net4960 _03605_ net4994 VGND VGND VPWR VPWR _04145_ sky130_fd_sc_hd__o21a_1
X_21497_ net5416 net5894 VGND VGND VPWR VPWR _01510_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5813 net5814 VGND VGND VPWR VPWR net5813 sky130_fd_sc_hd__buf_1
Xwire6558 net6559 VGND VGND VPWR VPWR net6558 sky130_fd_sc_hd__buf_1
XFILLER_0_127_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire6569 net6567 VGND VGND VPWR VPWR net6569 sky130_fd_sc_hd__buf_1
Xwire5824 net5825 VGND VGND VPWR VPWR net5824 sky130_fd_sc_hd__clkbuf_1
X_23236_ _02974_ _02975_ VGND VGND VPWR VPWR _03106_ sky130_fd_sc_hd__xnor2_1
Xwire5835 net5837 VGND VGND VPWR VPWR net5835 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20448_ net6511 _12133_ _12145_ _12233_ VGND VGND VPWR VPWR _12241_ sky130_fd_sc_hd__a22o_1
Xwire5846 net5840 VGND VGND VPWR VPWR net5846 sky130_fd_sc_hd__clkbuf_1
Xwire5857 net5858 VGND VGND VPWR VPWR net5857 sky130_fd_sc_hd__buf_1
XFILLER_0_132_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5868 net5869 VGND VGND VPWR VPWR net5868 sky130_fd_sc_hd__buf_1
Xwire5879 net5880 VGND VGND VPWR VPWR net5879 sky130_fd_sc_hd__buf_1
X_23167_ _03030_ _03036_ VGND VGND VPWR VPWR _03037_ sky130_fd_sc_hd__xnor2_1
X_20379_ net4055 _12159_ _12168_ VGND VGND VPWR VPWR _12178_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22118_ net5497 net5672 VGND VGND VPWR VPWR _02124_ sky130_fd_sc_hd__nand2_1
X_23098_ _02966_ _02967_ VGND VGND VPWR VPWR _02968_ sky130_fd_sc_hd__xor2_2
XFILLER_0_100_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22049_ net2067 _01965_ _02054_ _02055_ VGND VGND VPWR VPWR _02056_ sky130_fd_sc_hd__a31o_1
X_14940_ net6536 net6588 matmul0.matmul_stage_inst.e\[6\] VGND VGND VPWR VPWR _07014_
+ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_121_Left_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14871_ _06953_ VGND VGND VPWR VPWR _00206_ sky130_fd_sc_hd__clkbuf_1
X_16610_ matmul0.matmul_stage_inst.mult2\[12\] net209 net3468 VGND VGND VPWR VPWR
+ _08655_ sky130_fd_sc_hd__mux2_1
X_13822_ _06050_ net840 VGND VGND VPWR VPWR _06089_ sky130_fd_sc_hd__nor2_1
X_25808_ clknet_leaf_38_clk _00681_ net8755 VGND VGND VPWR VPWR pid_q.prev_error\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_17590_ svm0.calc_ready net2568 net769 net9000 net3384 VGND VGND VPWR VPWR _00407_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_35_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13753_ _05992_ net503 _06000_ VGND VGND VPWR VPWR _06021_ sky130_fd_sc_hd__o21ai_1
X_16541_ net1084 net976 net879 _08595_ _08599_ VGND VGND VPWR VPWR _08600_ sky130_fd_sc_hd__a311o_1
X_25739_ clknet_leaf_13_clk _00612_ net8608 VGND VGND VPWR VPWR pid_d.ki\[13\] sky130_fd_sc_hd__dfrtp_1
X_12704_ net4260 net1960 VGND VGND VPWR VPWR _04977_ sky130_fd_sc_hd__nor2_1
X_19260_ _11045_ _11094_ _11096_ VGND VGND VPWR VPWR _11097_ sky130_fd_sc_hd__or3b_1
X_13684_ _05945_ _05952_ VGND VGND VPWR VPWR _05953_ sky130_fd_sc_hd__xnor2_1
X_16472_ _08521_ _08532_ VGND VGND VPWR VPWR _08533_ sky130_fd_sc_hd__xor2_1
XFILLER_0_167_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18211_ net2552 _10060_ _10061_ VGND VGND VPWR VPWR _10062_ sky130_fd_sc_hd__a21o_1
X_12635_ net7852 net1985 net2363 VGND VGND VPWR VPWR _04908_ sky130_fd_sc_hd__and3_1
X_15423_ net2229 net1866 net1868 VGND VGND VPWR VPWR _07497_ sky130_fd_sc_hd__o21a_1
X_19191_ _10955_ _10880_ VGND VGND VPWR VPWR _11028_ sky130_fd_sc_hd__xor2_2
XFILLER_0_127_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout8388 net8415 VGND VGND VPWR VPWR net8388 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_130_Left_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18142_ _09987_ _09944_ _09989_ _09939_ VGND VGND VPWR VPWR _09993_ sky130_fd_sc_hd__o22a_1
X_15354_ _07418_ _07423_ _07427_ VGND VGND VPWR VPWR _07428_ sky130_fd_sc_hd__a21o_1
Xfanout7665 net7675 VGND VGND VPWR VPWR net7665 sky130_fd_sc_hd__buf_1
X_12566_ _04855_ VGND VGND VPWR VPWR _04856_ sky130_fd_sc_hd__buf_2
XFILLER_0_53_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8472 net8471 VGND VGND VPWR VPWR net8472 sky130_fd_sc_hd__buf_1
XFILLER_0_14_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8483 net8485 VGND VGND VPWR VPWR net8483 sky130_fd_sc_hd__buf_1
XFILLER_0_182_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8494 net8492 VGND VGND VPWR VPWR net8494 sky130_fd_sc_hd__buf_1
Xwire7760 net7761 VGND VGND VPWR VPWR net7760 sky130_fd_sc_hd__buf_1
X_14305_ _06526_ VGND VGND VPWR VPWR _06527_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15285_ net1901 _07357_ _07358_ VGND VGND VPWR VPWR _07359_ sky130_fd_sc_hd__a21o_1
X_18073_ _09849_ _09906_ _09907_ VGND VGND VPWR VPWR _09924_ sky130_fd_sc_hd__and3_1
Xwire162 net163 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_1
Xwire173 _08592_ VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_1
Xwire7793 net7794 VGND VGND VPWR VPWR net7793 sky130_fd_sc_hd__buf_1
XFILLER_0_34_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length3480 _07151_ VGND VGND VPWR VPWR net3480 sky130_fd_sc_hd__clkbuf_1
Xwire184 net185 VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_1
Xhold209 svm0.delta\[13\] VGND VGND VPWR VPWR net9162 sky130_fd_sc_hd__dlygate4sd3_1
X_14236_ net1304 _06492_ VGND VGND VPWR VPWR _06493_ sky130_fd_sc_hd__and2_1
X_17024_ net7029 VGND VGND VPWR VPWR _08984_ sky130_fd_sc_hd__inv_2
Xwire195 _04505_ VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14167_ _06427_ _06394_ _06425_ _06366_ VGND VGND VPWR VPWR _06428_ sky130_fd_sc_hd__o22a_1
X_13118_ net7736 _05011_ _05250_ net1619 net7783 VGND VGND VPWR VPWR _05391_ sky130_fd_sc_hd__a32oi_2
X_14098_ net282 net319 _06359_ VGND VGND VPWR VPWR _06361_ sky130_fd_sc_hd__a21o_1
X_18975_ net6270 net6290 VGND VGND VPWR VPWR _10812_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13049_ net789 _05004_ VGND VGND VPWR VPWR _05322_ sky130_fd_sc_hd__nand2_1
X_17926_ _09761_ _09771_ VGND VGND VPWR VPWR _09777_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17857_ _08984_ net7105 _09707_ VGND VGND VPWR VPWR _09708_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16808_ _08794_ VGND VGND VPWR VPWR _00302_ sky130_fd_sc_hd__clkbuf_1
X_17788_ net3260 net3259 VGND VGND VPWR VPWR _09639_ sky130_fd_sc_hd__xnor2_1
X_19527_ _11306_ _11307_ _11363_ VGND VGND VPWR VPWR _11364_ sky130_fd_sc_hd__mux2_1
X_16739_ net7568 matmul0.b\[6\] net3702 VGND VGND VPWR VPWR _08758_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19458_ _10974_ net2521 VGND VGND VPWR VPWR _11295_ sky130_fd_sc_hd__nor2_1
X_18409_ _10203_ _10259_ VGND VGND VPWR VPWR _10260_ sky130_fd_sc_hd__xor2_1
X_19389_ net6358 _11225_ VGND VGND VPWR VPWR _11226_ sky130_fd_sc_hd__nor2_1
XFILLER_0_189_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21420_ net4298 _01432_ _01433_ VGND VGND VPWR VPWR _01434_ sky130_fd_sc_hd__or3_1
XFILLER_0_86_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21351_ _01293_ _01294_ _01295_ VGND VGND VPWR VPWR _01365_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5109 net5110 VGND VGND VPWR VPWR net5109 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20302_ net6516 net2600 VGND VGND VPWR VPWR _12107_ sky130_fd_sc_hd__nand2_1
X_24070_ _03922_ _03931_ VGND VGND VPWR VPWR _03933_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21282_ _01293_ _01296_ VGND VGND VPWR VPWR _01297_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_188_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4408 net4409 VGND VGND VPWR VPWR net4408 sky130_fd_sc_hd__clkbuf_1
Xwire4419 net4420 VGND VGND VPWR VPWR net4419 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23021_ net4969 net4715 VGND VGND VPWR VPWR _02891_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20233_ net8122 _12050_ VGND VGND VPWR VPWR _12051_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3707 net3708 VGND VGND VPWR VPWR net3707 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3718 net3719 VGND VGND VPWR VPWR net3718 sky130_fd_sc_hd__buf_1
Xwire3729 _04531_ VGND VGND VPWR VPWR net3729 sky130_fd_sc_hd__clkbuf_1
X_20164_ net9006 net2122 net1444 _11990_ VGND VGND VPWR VPWR _00463_ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24972_ pid_q.kp\[5\] _04712_ net1357 VGND VGND VPWR VPWR _04741_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20095_ _11913_ _11922_ VGND VGND VPWR VPWR _11924_ sky130_fd_sc_hd__nand2_1
X_23923_ _03716_ _03718_ _03717_ VGND VGND VPWR VPWR _03787_ sky130_fd_sc_hd__o21ai_1
Xmax_length8425 net8423 VGND VGND VPWR VPWR net8425 sky130_fd_sc_hd__clkbuf_2
X_23854_ _03717_ _03718_ VGND VGND VPWR VPWR _03719_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22805_ _02710_ VGND VGND VPWR VPWR _00629_ sky130_fd_sc_hd__clkbuf_1
X_23785_ _03641_ _03650_ VGND VGND VPWR VPWR _03651_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20997_ _01011_ _01012_ VGND VGND VPWR VPWR _01013_ sky130_fd_sc_hd__nand2_1
Xmax_length7768 net7763 VGND VGND VPWR VPWR net7768 sky130_fd_sc_hd__buf_1
X_25524_ clknet_leaf_48_clk _00404_ net8759 VGND VGND VPWR VPWR svm0.counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_22736_ pid_d.ki\[3\] _02668_ net1688 VGND VGND VPWR VPWR _02669_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25455_ clknet_4_1__leaf_clk _00338_ net8362 VGND VGND VPWR VPWR cordic0.vec\[1\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_22667_ pid_d.ki\[0\] net3010 net2994 pid_d.kp\[0\] VGND VGND VPWR VPWR _02619_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24406_ net588 net587 VGND VGND VPWR VPWR _04264_ sky130_fd_sc_hd__nand2_1
Xwire7001 net7002 VGND VGND VPWR VPWR net7001 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21618_ _01447_ _01519_ _01629_ VGND VGND VPWR VPWR _01630_ sky130_fd_sc_hd__o21a_1
Xwire7023 net7018 VGND VGND VPWR VPWR net7023 sky130_fd_sc_hd__buf_1
X_25386_ clknet_leaf_74_clk _00269_ net8466 VGND VGND VPWR VPWR matmul0.b\[5\] sky130_fd_sc_hd__dfrtp_1
X_22598_ net4226 _02569_ VGND VGND VPWR VPWR _02574_ sky130_fd_sc_hd__nand2_1
Xclkbuf_4_7__f_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_4_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xwire6300 net6297 VGND VGND VPWR VPWR net6300 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_30_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7045 net7043 VGND VGND VPWR VPWR net7045 sky130_fd_sc_hd__buf_1
X_24337_ net634 net633 _04195_ VGND VGND VPWR VPWR _04196_ sky130_fd_sc_hd__o21ai_1
Xwire7056 net7057 VGND VGND VPWR VPWR net7056 sky130_fd_sc_hd__buf_1
X_21549_ _01557_ _01560_ VGND VGND VPWR VPWR _01561_ sky130_fd_sc_hd__xnor2_1
Xwire7078 net7079 VGND VGND VPWR VPWR net7078 sky130_fd_sc_hd__buf_1
Xfanout5548 pid_d.mult0.a\[6\] VGND VGND VPWR VPWR net5548 sky130_fd_sc_hd__buf_1
Xwire6355 net6357 VGND VGND VPWR VPWR net6355 sky130_fd_sc_hd__buf_1
Xfanout4814 pid_q.mult0.b\[14\] VGND VGND VPWR VPWR net4814 sky130_fd_sc_hd__buf_1
X_15070_ net6546 net6594 net7386 VGND VGND VPWR VPWR _07144_ sky130_fd_sc_hd__o21a_1
X_24268_ _04126_ _04127_ VGND VGND VPWR VPWR _04128_ sky130_fd_sc_hd__xor2_2
Xwire5621 net5622 VGND VGND VPWR VPWR net5621 sky130_fd_sc_hd__buf_1
Xwire6366 net6367 VGND VGND VPWR VPWR net6366 sky130_fd_sc_hd__clkbuf_1
Xwire5632 net5633 VGND VGND VPWR VPWR net5632 sky130_fd_sc_hd__clkbuf_1
Xwire5643 net5639 VGND VGND VPWR VPWR net5643 sky130_fd_sc_hd__buf_1
Xwire6388 net6389 VGND VGND VPWR VPWR net6388 sky130_fd_sc_hd__clkbuf_1
X_14021_ net7702 net1324 _06230_ net1316 net7718 VGND VGND VPWR VPWR _06285_ sky130_fd_sc_hd__a32o_1
Xmax_length1341 net1342 VGND VGND VPWR VPWR net1341 sky130_fd_sc_hd__clkbuf_1
Xwire5654 net5655 VGND VGND VPWR VPWR net5654 sky130_fd_sc_hd__clkbuf_2
Xwire6399 net6400 VGND VGND VPWR VPWR net6399 sky130_fd_sc_hd__buf_1
X_23219_ _03085_ _03087_ _03088_ _03084_ _03083_ VGND VGND VPWR VPWR _03089_ sky130_fd_sc_hd__a32o_1
Xwire5665 net5666 VGND VGND VPWR VPWR net5665 sky130_fd_sc_hd__clkbuf_1
Xwire4931 net4932 VGND VGND VPWR VPWR net4931 sky130_fd_sc_hd__clkbuf_1
X_24199_ _03986_ _03988_ _04059_ VGND VGND VPWR VPWR _04060_ sky130_fd_sc_hd__a21bo_1
Xwire5676 net5677 VGND VGND VPWR VPWR net5676 sky130_fd_sc_hd__buf_1
Xwire4942 net4943 VGND VGND VPWR VPWR net4942 sky130_fd_sc_hd__buf_1
Xwire5687 net5685 VGND VGND VPWR VPWR net5687 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4953 net4954 VGND VGND VPWR VPWR net4953 sky130_fd_sc_hd__buf_1
Xwire5698 net5699 VGND VGND VPWR VPWR net5698 sky130_fd_sc_hd__clkbuf_1
Xwire4964 net4962 VGND VGND VPWR VPWR net4964 sky130_fd_sc_hd__buf_1
Xwire4975 net4976 VGND VGND VPWR VPWR net4975 sky130_fd_sc_hd__clkbuf_1
Xwire4986 net4987 VGND VGND VPWR VPWR net4986 sky130_fd_sc_hd__buf_1
Xwire4997 net4998 VGND VGND VPWR VPWR net4997 sky130_fd_sc_hd__buf_1
X_18760_ _10516_ net764 _10561_ VGND VGND VPWR VPWR _10605_ sky130_fd_sc_hd__a21o_1
X_15972_ net3436 VGND VGND VPWR VPWR _08040_ sky130_fd_sc_hd__buf_1
X_17711_ pid_q.prev_int\[2\] net1218 net1452 net5180 VGND VGND VPWR VPWR _00416_ sky130_fd_sc_hd__a22o_1
X_14923_ net6613 net6638 matmul0.matmul_stage_inst.f\[4\] VGND VGND VPWR VPWR _06997_
+ sky130_fd_sc_hd__o21a_1
X_18691_ _10533_ _10536_ VGND VGND VPWR VPWR _10537_ sky130_fd_sc_hd__xnor2_1
Xhold70 pid_q.target\[2\] VGND VGND VPWR VPWR net9023 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 matmul0.matmul_stage_inst.c\[8\] VGND VGND VPWR VPWR net9034 sky130_fd_sc_hd__dlygate4sd3_1
X_17642_ _09520_ _09521_ VGND VGND VPWR VPWR _09522_ sky130_fd_sc_hd__or2_1
Xhold92 matmul0.matmul_stage_inst.d\[8\] VGND VGND VPWR VPWR net9045 sky130_fd_sc_hd__dlygate4sd3_1
X_14854_ _06944_ VGND VGND VPWR VPWR _00198_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13805_ _06067_ _06072_ VGND VGND VPWR VPWR _06073_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_188_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17573_ _09444_ _09445_ _09450_ _09454_ VGND VGND VPWR VPWR _09455_ sky130_fd_sc_hd__and4b_1
X_14785_ _06818_ net7148 VGND VGND VPWR VPWR _06908_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19312_ _11049_ _10838_ _11148_ net6354 VGND VGND VPWR VPWR _11149_ sky130_fd_sc_hd__a22o_1
X_16524_ _08524_ _08530_ _08471_ VGND VGND VPWR VPWR _08584_ sky130_fd_sc_hd__a21bo_1
X_13736_ _05872_ _06003_ _06004_ VGND VGND VPWR VPWR _06005_ sky130_fd_sc_hd__o21a_1
XFILLER_0_168_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19243_ net3877 _11079_ VGND VGND VPWR VPWR _11080_ sky130_fd_sc_hd__xor2_1
X_16455_ net2744 net2204 net2750 VGND VGND VPWR VPWR _08516_ sky130_fd_sc_hd__a21o_1
X_13667_ net9149 net1127 net284 net1927 VGND VGND VPWR VPWR _00019_ sky130_fd_sc_hd__a22o_1
X_15406_ net3573 net3569 net4105 net4101 VGND VGND VPWR VPWR _07480_ sky130_fd_sc_hd__o22a_1
Xfanout7440 net7443 VGND VGND VPWR VPWR net7440 sky130_fd_sc_hd__buf_1
X_12618_ net2992 VGND VGND VPWR VPWR _04891_ sky130_fd_sc_hd__clkbuf_1
X_19174_ _10994_ _11010_ VGND VGND VPWR VPWR _11011_ sky130_fd_sc_hd__xnor2_1
X_13598_ _05867_ VGND VGND VPWR VPWR _05868_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16386_ net2625 net2218 VGND VGND VPWR VPWR _08448_ sky130_fd_sc_hd__nor2_1
Xfanout7462 net7469 VGND VGND VPWR VPWR net7462 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8280 net8281 VGND VGND VPWR VPWR net8280 sky130_fd_sc_hd__clkbuf_1
X_18125_ net3255 _09748_ _09973_ net7061 _09975_ VGND VGND VPWR VPWR _09976_ sky130_fd_sc_hd__a221o_1
XFILLER_0_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8291 net8292 VGND VGND VPWR VPWR net8291 sky130_fd_sc_hd__clkbuf_1
X_15337_ _07405_ _07410_ VGND VGND VPWR VPWR _07411_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout6772 net6787 VGND VGND VPWR VPWR net6772 sky130_fd_sc_hd__buf_1
XFILLER_0_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1 clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18056_ _08913_ net3257 net3969 net7062 VGND VGND VPWR VPWR _09907_ sky130_fd_sc_hd__a211o_1
Xwire7590 net7591 VGND VGND VPWR VPWR net7590 sky130_fd_sc_hd__clkbuf_1
X_15268_ net991 _07213_ net830 _07217_ VGND VGND VPWR VPWR _07342_ sky130_fd_sc_hd__o22ai_2
X_17007_ net6480 net3364 VGND VGND VPWR VPWR _08968_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14219_ _06476_ _06477_ VGND VGND VPWR VPWR _06478_ sky130_fd_sc_hd__and2b_1
X_15199_ net4190 net4184 net4121 net4116 VGND VGND VPWR VPWR _07273_ sky130_fd_sc_hd__o22a_1
XFILLER_0_158_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18958_ net6298 _10794_ VGND VGND VPWR VPWR _10795_ sky130_fd_sc_hd__or2_2
XFILLER_0_174_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17909_ _09756_ _09758_ _09759_ VGND VGND VPWR VPWR _09760_ sky130_fd_sc_hd__o21a_1
X_18889_ net302 _10730_ VGND VGND VPWR VPWR _10731_ sky130_fd_sc_hd__xor2_1
X_20920_ net1392 net1187 VGND VGND VPWR VPWR _00936_ sky130_fd_sc_hd__nand2_1
XFILLER_0_174_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20851_ net5906 _00865_ _00866_ VGND VGND VPWR VPWR _00867_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23570_ _03432_ _03437_ VGND VGND VPWR VPWR _03438_ sky130_fd_sc_hd__xnor2_1
X_20782_ net5596 net5578 net5776 net5794 VGND VGND VPWR VPWR _12553_ sky130_fd_sc_hd__nand4_1
XFILLER_0_49_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22521_ net4325 net2462 net8887 VGND VGND VPWR VPWR _02521_ sky130_fd_sc_hd__o21a_1
Xmax_length4928 net4929 VGND VGND VPWR VPWR net4928 sky130_fd_sc_hd__buf_1
XFILLER_0_146_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4939 net4933 VGND VGND VPWR VPWR net4939 sky130_fd_sc_hd__clkbuf_1
X_25240_ clknet_leaf_69_clk _00123_ net8468 VGND VGND VPWR VPWR matmul0.op\[1\] sky130_fd_sc_hd__dfrtp_1
Xwire909 net910 VGND VGND VPWR VPWR net909 sky130_fd_sc_hd__buf_1
X_22452_ _02450_ _02453_ VGND VGND VPWR VPWR _02454_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21403_ _00838_ net1393 net1050 _01313_ _01255_ VGND VGND VPWR VPWR _01417_ sky130_fd_sc_hd__a221o_1
X_25171_ clknet_leaf_54_clk _00060_ net8729 VGND VGND VPWR VPWR svm0.periodTop\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_22383_ net551 net549 VGND VGND VPWR VPWR _02386_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24122_ _03893_ _03895_ _03894_ VGND VGND VPWR VPWR _03984_ sky130_fd_sc_hd__o21ai_1
X_21334_ net5687 net5616 VGND VGND VPWR VPWR _01348_ sky130_fd_sc_hd__and2_1
XFILLER_0_163_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24053_ _03911_ _03913_ VGND VGND VPWR VPWR _03916_ sky130_fd_sc_hd__nor2_1
Xwire4216 net4217 VGND VGND VPWR VPWR net4216 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_163_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4227 net4228 VGND VGND VPWR VPWR net4227 sky130_fd_sc_hd__clkbuf_1
X_21265_ net5761 net5570 VGND VGND VPWR VPWR _01280_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4249 net4250 VGND VGND VPWR VPWR net4249 sky130_fd_sc_hd__buf_1
Xwire3504 net3505 VGND VGND VPWR VPWR net3504 sky130_fd_sc_hd__clkbuf_1
X_23004_ _02872_ _02873_ VGND VGND VPWR VPWR _02874_ sky130_fd_sc_hd__xor2_1
Xwire3515 net3517 VGND VGND VPWR VPWR net3515 sky130_fd_sc_hd__clkbuf_1
X_20216_ net8 _12037_ VGND VGND VPWR VPWR _12038_ sky130_fd_sc_hd__xnor2_1
Xwire3526 net3527 VGND VGND VPWR VPWR net3526 sky130_fd_sc_hd__buf_1
X_21196_ _01166_ _01202_ _01210_ net5881 _01211_ VGND VGND VPWR VPWR _01212_ sky130_fd_sc_hd__a221o_1
Xwire3537 net3538 VGND VGND VPWR VPWR net3537 sky130_fd_sc_hd__buf_1
Xwire2803 net2804 VGND VGND VPWR VPWR net2803 sky130_fd_sc_hd__buf_1
Xwire3548 net3549 VGND VGND VPWR VPWR net3548 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_4_15__f_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_4_15__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_159_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3559 net3560 VGND VGND VPWR VPWR net3559 sky130_fd_sc_hd__buf_1
Xwire2814 _07100_ VGND VGND VPWR VPWR net2814 sky130_fd_sc_hd__buf_1
Xwire2825 _07087_ VGND VGND VPWR VPWR net2825 sky130_fd_sc_hd__clkbuf_1
X_20147_ _11938_ _11973_ VGND VGND VPWR VPWR _11974_ sky130_fd_sc_hd__xnor2_1
Xwire2836 net2837 VGND VGND VPWR VPWR net2836 sky130_fd_sc_hd__buf_1
Xwire2847 net2848 VGND VGND VPWR VPWR net2847 sky130_fd_sc_hd__clkbuf_1
Xwire2858 net2859 VGND VGND VPWR VPWR net2858 sky130_fd_sc_hd__buf_1
Xwire2869 _06820_ VGND VGND VPWR VPWR net2869 sky130_fd_sc_hd__buf_1
X_24955_ pid_q.ki\[14\] _04730_ net1637 VGND VGND VPWR VPWR _04731_ sky130_fd_sc_hd__mux2_1
X_20078_ net2581 net2092 VGND VGND VPWR VPWR _11907_ sky130_fd_sc_hd__nor2_1
X_23906_ pid_q.prev_int\[5\] VGND VGND VPWR VPWR _03770_ sky130_fd_sc_hd__inv_2
X_24886_ pid_q.ki\[10\] net2398 net3700 pid_q.kp\[10\] VGND VGND VPWR VPWR _04682_
+ sky130_fd_sc_hd__a22o_1
Xmax_length7510 net7511 VGND VGND VPWR VPWR net7510 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_196_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23837_ net5096 net3744 _03519_ VGND VGND VPWR VPWR _03702_ sky130_fd_sc_hd__and3_1
Xmax_length6820 net6821 VGND VGND VPWR VPWR net6820 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14570_ _06730_ _06731_ _06739_ VGND VGND VPWR VPWR _06747_ sky130_fd_sc_hd__o21a_1
Xmax_length7576 matmul0.b_in\[0\] VGND VGND VPWR VPWR net7576 sky130_fd_sc_hd__clkbuf_1
X_23768_ net1661 _03633_ VGND VGND VPWR VPWR _03634_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13521_ net7838 net1577 VGND VGND VPWR VPWR _05792_ sky130_fd_sc_hd__nand2_1
X_25507_ clknet_leaf_39_clk _00387_ net8754 VGND VGND VPWR VPWR svm0.delta\[12\] sky130_fd_sc_hd__dfrtp_1
X_22719_ net8096 net8098 net8106 net86 VGND VGND VPWR VPWR _02655_ sky130_fd_sc_hd__or4_1
XFILLER_0_95_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23699_ _03486_ _03565_ VGND VGND VPWR VPWR _03566_ sky130_fd_sc_hd__xnor2_1
X_13452_ net916 _05724_ VGND VGND VPWR VPWR _05725_ sky130_fd_sc_hd__xnor2_1
X_16240_ _08241_ _08304_ VGND VGND VPWR VPWR _08305_ sky130_fd_sc_hd__xnor2_1
X_25438_ clknet_leaf_94_clk _00321_ net8426 VGND VGND VPWR VPWR matmul0.sin\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_165_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6024 net6036 VGND VGND VPWR VPWR net6024 sky130_fd_sc_hd__buf_1
Xfanout6035 cordic0.vec\[0\]\[16\] VGND VGND VPWR VPWR net6035 sky130_fd_sc_hd__buf_1
X_13383_ _05553_ _05561_ VGND VGND VPWR VPWR _05656_ sky130_fd_sc_hd__nand2_1
X_25369_ clknet_leaf_81_clk _00252_ net8500 VGND VGND VPWR VPWR matmul0.alpha_pass\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_16171_ matmul0.matmul_stage_inst.mult1\[8\] net311 net2681 VGND VGND VPWR VPWR _08237_
+ sky130_fd_sc_hd__mux2_1
Xfanout6068 net6075 VGND VGND VPWR VPWR net6068 sky130_fd_sc_hd__buf_1
XFILLER_0_63_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6130 net6127 VGND VGND VPWR VPWR net6130 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_51_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6141 net6142 VGND VGND VPWR VPWR net6141 sky130_fd_sc_hd__clkbuf_1
X_15122_ net3503 net3453 _07064_ _07195_ VGND VGND VPWR VPWR _07196_ sky130_fd_sc_hd__a22o_1
Xwire6152 net6151 VGND VGND VPWR VPWR net6152 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_181_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6163 net6159 VGND VGND VPWR VPWR net6163 sky130_fd_sc_hd__buf_1
Xwire6174 net6169 VGND VGND VPWR VPWR net6174 sky130_fd_sc_hd__buf_1
XFILLER_0_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5440 net5441 VGND VGND VPWR VPWR net5440 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19930_ net6065 net6049 VGND VGND VPWR VPWR _11762_ sky130_fd_sc_hd__nor2_1
X_15053_ net6610 net6534 matmul0.matmul_stage_inst.b\[0\] VGND VGND VPWR VPWR _07127_
+ sky130_fd_sc_hd__o21a_1
Xwire5451 net5452 VGND VGND VPWR VPWR net5451 sky130_fd_sc_hd__clkbuf_1
Xwire6196 net6197 VGND VGND VPWR VPWR net6196 sky130_fd_sc_hd__buf_1
XFILLER_0_32_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5462 net5466 VGND VGND VPWR VPWR net5462 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_128_Right_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5473 net5474 VGND VGND VPWR VPWR net5473 sky130_fd_sc_hd__clkbuf_2
X_14004_ _06265_ _06268_ VGND VGND VPWR VPWR _06269_ sky130_fd_sc_hd__xor2_1
Xwire5484 net5485 VGND VGND VPWR VPWR net5484 sky130_fd_sc_hd__buf_1
Xwire4750 net4751 VGND VGND VPWR VPWR net4750 sky130_fd_sc_hd__clkbuf_1
Xwire5495 net5490 VGND VGND VPWR VPWR net5495 sky130_fd_sc_hd__buf_1
X_19861_ _11503_ net3867 _11560_ _11693_ VGND VGND VPWR VPWR _11694_ sky130_fd_sc_hd__a22o_1
Xwire4772 net4771 VGND VGND VPWR VPWR net4772 sky130_fd_sc_hd__clkbuf_2
Xwire4783 net4779 VGND VGND VPWR VPWR net4783 sky130_fd_sc_hd__clkbuf_1
X_18812_ _10625_ _10655_ VGND VGND VPWR VPWR _10656_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19792_ net3862 _11625_ VGND VGND VPWR VPWR _11626_ sky130_fd_sc_hd__or2b_1
XFILLER_0_37_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18743_ _10530_ _10486_ _10531_ net6796 _10587_ VGND VGND VPWR VPWR _10588_ sky130_fd_sc_hd__a221o_1
X_15955_ _08019_ _08022_ VGND VGND VPWR VPWR _08023_ sky130_fd_sc_hd__xnor2_1
X_14906_ _06968_ _06979_ VGND VGND VPWR VPWR _06980_ sky130_fd_sc_hd__xnor2_1
X_18674_ net1431 _10483_ _10519_ VGND VGND VPWR VPWR _10520_ sky130_fd_sc_hd__a21o_1
X_15886_ net4071 _07952_ _07953_ net2718 _07954_ VGND VGND VPWR VPWR _07955_ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17625_ net4018 svm0.tB\[3\] svm0.tB\[2\] _09451_ _09505_ VGND VGND VPWR VPWR _09506_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_187_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14837_ _06935_ VGND VGND VPWR VPWR _00190_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17556_ _09434_ _09436_ _09437_ VGND VGND VPWR VPWR _09438_ sky130_fd_sc_hd__and3b_1
XFILLER_0_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14768_ net7448 net7149 VGND VGND VPWR VPWR _06896_ sky130_fd_sc_hd__nand2_1
X_16507_ net2638 _08563_ _08565_ _08566_ VGND VGND VPWR VPWR _08567_ sky130_fd_sc_hd__and4_1
X_13719_ net7831 net1929 VGND VGND VPWR VPWR _05988_ sky130_fd_sc_hd__nand2_1
X_17487_ _09299_ _09372_ net4005 VGND VGND VPWR VPWR _09377_ sky130_fd_sc_hd__o21a_1
X_14699_ net9094 net2862 net2262 net1910 VGND VGND VPWR VPWR _00143_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19226_ net3178 _11056_ _11048_ VGND VGND VPWR VPWR _11063_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16438_ _08476_ _08497_ _08498_ VGND VGND VPWR VPWR _08499_ sky130_fd_sc_hd__o21a_1
XFILLER_0_183_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19157_ _10982_ _10993_ VGND VGND VPWR VPWR _10994_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_15_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16369_ net303 _08431_ VGND VGND VPWR VPWR _08432_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_169_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18108_ _09954_ _09958_ VGND VGND VPWR VPWR _09959_ sky130_fd_sc_hd__xnor2_1
Xfanout6580 net6585 VGND VGND VPWR VPWR net6580 sky130_fd_sc_hd__buf_1
X_19088_ net3191 _10924_ _10911_ VGND VGND VPWR VPWR _10925_ sky130_fd_sc_hd__a21o_1
Xfanout6591 matmul0.matmul_stage_inst.state\[4\] VGND VGND VPWR VPWR net6591 sky130_fd_sc_hd__buf_1
X_18039_ _09889_ _09026_ net2555 VGND VGND VPWR VPWR _09890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21050_ net5567 VGND VGND VPWR VPWR _01066_ sky130_fd_sc_hd__inv_2
X_20001_ net351 net487 _11825_ _11828_ _11831_ VGND VGND VPWR VPWR _11832_ sky130_fd_sc_hd__a32o_1
XFILLER_0_185_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1409 _11760_ VGND VGND VPWR VPWR net1409 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_185_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24740_ net8007 _04567_ VGND VGND VPWR VPWR _04572_ sky130_fd_sc_hd__or2_1
X_21952_ net2474 _01854_ _01850_ VGND VGND VPWR VPWR _01960_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_55_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20903_ net5906 _00896_ _00898_ VGND VGND VPWR VPWR _00919_ sky130_fd_sc_hd__o21a_1
X_24671_ pid_q.curr_error\[7\] net2384 net1373 VGND VGND VPWR VPWR _04518_ sky130_fd_sc_hd__and3_1
X_21883_ _01885_ _01891_ VGND VGND VPWR VPWR _01892_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23622_ net4677 net4875 VGND VGND VPWR VPWR _03489_ sky130_fd_sc_hd__nand2_2
XFILLER_0_89_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20834_ _00844_ _00849_ VGND VGND VPWR VPWR _00850_ sky130_fd_sc_hd__xnor2_1
Xmax_length5404 net5405 VGND VGND VPWR VPWR net5404 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23553_ _03415_ _03420_ VGND VGND VPWR VPWR _03421_ sky130_fd_sc_hd__xnor2_2
Xmax_length5437 net5438 VGND VGND VPWR VPWR net5437 sky130_fd_sc_hd__clkbuf_1
X_20765_ _12520_ _12535_ VGND VGND VPWR VPWR _12536_ sky130_fd_sc_hd__xor2_2
XFILLER_0_92_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22504_ _02447_ _02504_ _02502_ VGND VGND VPWR VPWR _02505_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23484_ _03351_ _03352_ VGND VGND VPWR VPWR _03353_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20696_ net3132 _12469_ _12470_ VGND VGND VPWR VPWR _00515_ sky130_fd_sc_hd__a21oi_1
Xwire706 _01251_ VGND VGND VPWR VPWR net706 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire717 net718 VGND VGND VPWR VPWR net717 sky130_fd_sc_hd__clkbuf_1
Xwire728 net729 VGND VGND VPWR VPWR net728 sky130_fd_sc_hd__buf_1
X_25223_ clknet_leaf_60_clk _00112_ net8690 VGND VGND VPWR VPWR svm0.vC\[11\] sky130_fd_sc_hd__dfrtp_1
Xwire739 net740 VGND VGND VPWR VPWR net739 sky130_fd_sc_hd__buf_1
X_22435_ _02431_ _02436_ VGND VGND VPWR VPWR _02437_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25154_ clknet_leaf_41_clk _00043_ net8767 VGND VGND VPWR VPWR pid_q.target\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_22366_ _02283_ _02302_ _02368_ VGND VGND VPWR VPWR _02369_ sky130_fd_sc_hd__o21a_1
XFILLER_0_131_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24105_ _03965_ _03966_ VGND VGND VPWR VPWR _03967_ sky130_fd_sc_hd__xnor2_1
Xwire4002 net4003 VGND VGND VPWR VPWR net4002 sky130_fd_sc_hd__buf_1
XFILLER_0_14_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21317_ pid_d.prev_error\[1\] net5972 VGND VGND VPWR VPWR _01332_ sky130_fd_sc_hd__xnor2_1
Xwire4013 _09339_ VGND VGND VPWR VPWR net4013 sky130_fd_sc_hd__buf_1
X_25085_ net5174 _04824_ net4406 VGND VGND VPWR VPWR _04830_ sky130_fd_sc_hd__a21o_1
Xwire4024 net4025 VGND VGND VPWR VPWR net4024 sky130_fd_sc_hd__clkbuf_1
X_22297_ net3778 _02229_ _02300_ VGND VGND VPWR VPWR _02301_ sky130_fd_sc_hd__or3_1
XFILLER_0_131_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24036_ _03782_ _03784_ _03898_ VGND VGND VPWR VPWR _03899_ sky130_fd_sc_hd__a21bo_1
Xwire4046 _08954_ VGND VGND VPWR VPWR net4046 sky130_fd_sc_hd__clkbuf_2
Xwire3301 net3302 VGND VGND VPWR VPWR net3301 sky130_fd_sc_hd__buf_1
Xwire4057 net4058 VGND VGND VPWR VPWR net4057 sky130_fd_sc_hd__buf_1
Xwire3312 _09051_ VGND VGND VPWR VPWR net3312 sky130_fd_sc_hd__buf_1
X_21248_ _00826_ _00827_ _01262_ VGND VGND VPWR VPWR _01263_ sky130_fd_sc_hd__a21bo_1
Xwire3323 net3324 VGND VGND VPWR VPWR net3323 sky130_fd_sc_hd__buf_1
Xwire3334 net3335 VGND VGND VPWR VPWR net3334 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire4079 net4080 VGND VGND VPWR VPWR net4079 sky130_fd_sc_hd__buf_1
Xwire2600 net2601 VGND VGND VPWR VPWR net2600 sky130_fd_sc_hd__buf_1
Xwire2611 _08882_ VGND VGND VPWR VPWR net2611 sky130_fd_sc_hd__clkbuf_1
Xwire3356 _08909_ VGND VGND VPWR VPWR net3356 sky130_fd_sc_hd__clkbuf_1
X_21179_ _01194_ VGND VGND VPWR VPWR _01195_ sky130_fd_sc_hd__inv_2
Xwire3367 _08792_ VGND VGND VPWR VPWR net3367 sky130_fd_sc_hd__clkbuf_2
Xwire2622 _08450_ VGND VGND VPWR VPWR net2622 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2633 _07866_ VGND VGND VPWR VPWR net2633 sky130_fd_sc_hd__buf_1
Xwire3378 _08770_ VGND VGND VPWR VPWR net3378 sky130_fd_sc_hd__clkbuf_2
Xwire3389 _08645_ VGND VGND VPWR VPWR net3389 sky130_fd_sc_hd__buf_1
Xwire2655 net2657 VGND VGND VPWR VPWR net2655 sky130_fd_sc_hd__buf_1
Xwire1910 _06844_ VGND VGND VPWR VPWR net1910 sky130_fd_sc_hd__clkbuf_1
Xwire1921 net1922 VGND VGND VPWR VPWR net1921 sky130_fd_sc_hd__buf_1
XFILLER_0_99_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2666 net2667 VGND VGND VPWR VPWR net2666 sky130_fd_sc_hd__buf_1
XFILLER_0_99_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1932 net1933 VGND VGND VPWR VPWR net1932 sky130_fd_sc_hd__clkbuf_1
Xwire2677 _07579_ VGND VGND VPWR VPWR net2677 sky130_fd_sc_hd__buf_1
Xwire1943 net1944 VGND VGND VPWR VPWR net1943 sky130_fd_sc_hd__buf_1
Xwire2688 net2689 VGND VGND VPWR VPWR net2688 sky130_fd_sc_hd__clkbuf_1
Xwire1954 net1955 VGND VGND VPWR VPWR net1954 sky130_fd_sc_hd__buf_1
Xwire2699 _07438_ VGND VGND VPWR VPWR net2699 sky130_fd_sc_hd__buf_1
Xwire1965 net1966 VGND VGND VPWR VPWR net1965 sky130_fd_sc_hd__clkbuf_2
X_15740_ net2780 net2221 VGND VGND VPWR VPWR _07811_ sky130_fd_sc_hd__nor2_1
X_24938_ _04719_ VGND VGND VPWR VPWR _00753_ sky130_fd_sc_hd__clkbuf_1
Xwire1976 net1977 VGND VGND VPWR VPWR net1976 sky130_fd_sc_hd__buf_1
X_12952_ _05221_ _05222_ _05224_ VGND VGND VPWR VPWR _05225_ sky130_fd_sc_hd__a21oi_1
Xwire1987 net1989 VGND VGND VPWR VPWR net1987 sky130_fd_sc_hd__buf_1
Xwire1998 _04668_ VGND VGND VPWR VPWR net1998 sky130_fd_sc_hd__buf_1
XFILLER_0_169_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15671_ _07696_ _07701_ VGND VGND VPWR VPWR _07742_ sky130_fd_sc_hd__nor2_1
X_24869_ _04670_ net4707 net1996 VGND VGND VPWR VPWR _04671_ sky130_fd_sc_hd__mux2_1
X_12883_ net7848 _04956_ net2975 VGND VGND VPWR VPWR _05156_ sky130_fd_sc_hd__and3_1
X_17410_ net611 _09313_ _09311_ VGND VGND VPWR VPWR _09314_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14622_ net6446 cordic0.in_valid _06497_ VGND VGND VPWR VPWR _06792_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_185_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18390_ net6979 net7071 VGND VGND VPWR VPWR _10241_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_96_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length7395 matmul0.matmul_stage_inst.e\[4\] VGND VGND VPWR VPWR net7395 sky130_fd_sc_hd__clkbuf_1
X_17341_ _09228_ net1220 _09253_ _09254_ VGND VGND VPWR VPWR _09255_ sky130_fd_sc_hd__or4_1
X_14553_ net7264 net5238 VGND VGND VPWR VPWR _06731_ sky130_fd_sc_hd__or2_2
XFILLER_0_184_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6694 net6690 VGND VGND VPWR VPWR net6694 sky130_fd_sc_hd__clkbuf_2
X_13504_ net2961 net2984 VGND VGND VPWR VPWR _05777_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17272_ _09191_ net218 net1798 net9100 VGND VGND VPWR VPWR _00366_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14484_ net7336 net5287 VGND VGND VPWR VPWR _06669_ sky130_fd_sc_hd__xor2_2
XFILLER_0_99_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19011_ net6319 _10841_ _10844_ net6303 _10847_ VGND VGND VPWR VPWR _10848_ sky130_fd_sc_hd__a221o_1
X_16223_ _08286_ _08287_ VGND VGND VPWR VPWR _08288_ sky130_fd_sc_hd__or2b_1
X_13435_ net7901 net2946 net1938 VGND VGND VPWR VPWR _05708_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13366_ net7926 net1582 _05534_ _05533_ VGND VGND VPWR VPWR _05639_ sky130_fd_sc_hd__a31o_1
X_16154_ net3459 net2733 net3409 net1849 VGND VGND VPWR VPWR _08220_ sky130_fd_sc_hd__and4_1
XFILLER_0_2_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15105_ net4143 net4140 VGND VGND VPWR VPWR _07179_ sky130_fd_sc_hd__or2_1
X_13297_ _05567_ _05568_ _05569_ VGND VGND VPWR VPWR _05570_ sky130_fd_sc_hd__o21ai_2
X_16085_ _08066_ _08073_ VGND VGND VPWR VPWR _08152_ sky130_fd_sc_hd__nor2_1
Xwire5270 net5271 VGND VGND VPWR VPWR net5270 sky130_fd_sc_hd__buf_1
X_19913_ net6117 _11686_ net3869 VGND VGND VPWR VPWR _11745_ sky130_fd_sc_hd__mux2_1
X_15036_ _07097_ _07098_ VGND VGND VPWR VPWR _07110_ sky130_fd_sc_hd__xnor2_1
Xwire5281 net5282 VGND VGND VPWR VPWR net5281 sky130_fd_sc_hd__clkbuf_1
Xwire5292 net5293 VGND VGND VPWR VPWR net5292 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4580 net4581 VGND VGND VPWR VPWR net4580 sky130_fd_sc_hd__buf_1
X_19844_ net1188 _11675_ _11676_ VGND VGND VPWR VPWR _11677_ sky130_fd_sc_hd__a21oi_1
Xwire4591 net4592 VGND VGND VPWR VPWR net4591 sky130_fd_sc_hd__buf_1
XFILLER_0_43_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3890 _10879_ VGND VGND VPWR VPWR net3890 sky130_fd_sc_hd__buf_1
X_19775_ _11555_ _11558_ _11609_ VGND VGND VPWR VPWR _11610_ sky130_fd_sc_hd__a21o_1
X_16987_ net6309 net6254 net6277 net6216 net6498 net6518 VGND VGND VPWR VPWR _08949_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_64_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18726_ _10570_ net1430 _10543_ VGND VGND VPWR VPWR _10571_ sky130_fd_sc_hd__a21o_1
XFILLER_0_155_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15938_ _08003_ _08006_ VGND VGND VPWR VPWR _08007_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18657_ net605 _10456_ VGND VGND VPWR VPWR _10504_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15869_ net2650 net2657 VGND VGND VPWR VPWR _07938_ sky130_fd_sc_hd__nor2_1
X_17608_ svm0.tB\[8\] net4025 net6706 _09486_ VGND VGND VPWR VPWR _09489_ sky130_fd_sc_hd__o2bb2a_1
X_18588_ net6833 net6817 VGND VGND VPWR VPWR _10436_ sky130_fd_sc_hd__nand2_1
XFILLER_0_175_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17539_ svm0.tC\[13\] VGND VGND VPWR VPWR _09421_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20550_ net6326 _12301_ _12302_ VGND VGND VPWR VPWR _12335_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length3309 net3310 VGND VGND VPWR VPWR net3309 sky130_fd_sc_hd__buf_1
XFILLER_0_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19209_ net6152 VGND VGND VPWR VPWR _11046_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20481_ net6758 net3849 _08836_ VGND VGND VPWR VPWR _12270_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22220_ _02130_ _02131_ _02224_ VGND VGND VPWR VPWR _02225_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_113_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22151_ net1036 _02156_ VGND VGND VPWR VPWR _02157_ sky130_fd_sc_hd__xnor2_1
X_21102_ net5581 net5929 VGND VGND VPWR VPWR _01118_ sky130_fd_sc_hd__nand2_1
X_22082_ net2059 net1044 _02088_ VGND VGND VPWR VPWR _02089_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_196_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25910_ clknet_leaf_28_clk _00783_ net8656 VGND VGND VPWR VPWR pid_q.out\[6\] sky130_fd_sc_hd__dfrtp_1
X_21033_ net5629 VGND VGND VPWR VPWR _01049_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1206 _10325_ VGND VGND VPWR VPWR net1206 sky130_fd_sc_hd__clkbuf_1
X_25841_ clknet_leaf_20_clk _00714_ net8610 VGND VGND VPWR VPWR pid_q.mult0.b\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1228 net1229 VGND VGND VPWR VPWR net1228 sky130_fd_sc_hd__clkbuf_1
Xwire1239 _08917_ VGND VGND VPWR VPWR net1239 sky130_fd_sc_hd__buf_1
X_25772_ clknet_leaf_27_clk _00645_ net8650 VGND VGND VPWR VPWR pid_d.out\[13\] sky130_fd_sc_hd__dfrtp_1
X_22984_ net5218 net423 net6568 VGND VGND VPWR VPWR _02860_ sky130_fd_sc_hd__mux2_1
X_24723_ _04550_ _04551_ net8017 net4232 VGND VGND VPWR VPWR _04557_ sky130_fd_sc_hd__a211o_1
X_21935_ net5784 net5408 VGND VGND VPWR VPWR _01943_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24654_ net1647 VGND VGND VPWR VPWR _04508_ sky130_fd_sc_hd__buf_1
X_21866_ _01862_ net1718 VGND VGND VPWR VPWR _01875_ sky130_fd_sc_hd__xor2_1
Xmax_length5212 matmul0.beta_pass\[12\] VGND VGND VPWR VPWR net5212 sky130_fd_sc_hd__clkbuf_1
X_23605_ _03470_ _03472_ VGND VGND VPWR VPWR _03473_ sky130_fd_sc_hd__and2_1
X_20817_ _12513_ _12518_ _12508_ VGND VGND VPWR VPWR _00833_ sky130_fd_sc_hd__o21ba_1
Xwire8802 net8792 VGND VGND VPWR VPWR net8802 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24585_ _04410_ _04440_ VGND VGND VPWR VPWR _04441_ sky130_fd_sc_hd__xnor2_2
X_21797_ _01804_ _01806_ VGND VGND VPWR VPWR _01807_ sky130_fd_sc_hd__xor2_1
Xwire8824 net8825 VGND VGND VPWR VPWR net8824 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8835 net8836 VGND VGND VPWR VPWR net8835 sky130_fd_sc_hd__clkbuf_1
X_23536_ _03400_ _03403_ VGND VGND VPWR VPWR _03404_ sky130_fd_sc_hd__xnor2_1
X_20748_ _12513_ _12518_ VGND VGND VPWR VPWR _12519_ sky130_fd_sc_hd__xor2_1
Xwire8846 net8847 VGND VGND VPWR VPWR net8846 sky130_fd_sc_hd__clkbuf_1
Xmax_length5278 net5279 VGND VGND VPWR VPWR net5278 sky130_fd_sc_hd__buf_1
Xwire8857 net8858 VGND VGND VPWR VPWR net8857 sky130_fd_sc_hd__clkbuf_1
Xwire503 _05998_ VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__buf_1
Xmax_length4544 net4545 VGND VGND VPWR VPWR net4544 sky130_fd_sc_hd__clkbuf_1
Xwire8868 net8866 VGND VGND VPWR VPWR net8868 sky130_fd_sc_hd__buf_1
Xwire514 net515 VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__buf_1
Xwire8879 net8880 VGND VGND VPWR VPWR net8879 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23467_ _03269_ _03278_ _03277_ VGND VGND VPWR VPWR _03336_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_64_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire525 _01727_ VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_190_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire536 net537 VGND VGND VPWR VPWR net536 sky130_fd_sc_hd__clkbuf_1
X_20679_ net6091 _12445_ VGND VGND VPWR VPWR _12455_ sky130_fd_sc_hd__and2_1
Xwire547 net548 VGND VGND VPWR VPWR net547 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13220_ net7672 _05216_ _05458_ VGND VGND VPWR VPWR _05493_ sky130_fd_sc_hd__and3_1
Xwire558 net559 VGND VGND VPWR VPWR net558 sky130_fd_sc_hd__clkbuf_1
X_22418_ net5434 net5646 VGND VGND VPWR VPWR _02420_ sky130_fd_sc_hd__and2b_1
Xmax_length3865 _11436_ VGND VGND VPWR VPWR net3865 sky130_fd_sc_hd__clkbuf_1
Xwire569 net570 VGND VGND VPWR VPWR net569 sky130_fd_sc_hd__dlymetal6s2s_1
X_25206_ clknet_leaf_82_clk _00095_ net8709 VGND VGND VPWR VPWR matmul0.b_in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23398_ _03266_ _03267_ VGND VGND VPWR VPWR _03268_ sky130_fd_sc_hd__xor2_1
Xmax_length3887 net3888 VGND VGND VPWR VPWR net3887 sky130_fd_sc_hd__buf_1
XFILLER_0_100_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13151_ _05417_ _05418_ _05423_ VGND VGND VPWR VPWR _05424_ sky130_fd_sc_hd__nand3_1
X_25137_ clknet_leaf_51_clk _00026_ net8809 VGND VGND VPWR VPWR svm0.tC\[9\] sky130_fd_sc_hd__dfrtp_1
X_22349_ _01405_ net5647 VGND VGND VPWR VPWR _02352_ sky130_fd_sc_hd__nand2_2
X_13082_ net7933 _05353_ _05349_ _05354_ VGND VGND VPWR VPWR _05355_ sky130_fd_sc_hd__o2bb2a_1
X_25068_ net4424 _04813_ net193 net1629 _04815_ VGND VGND VPWR VPWR _00787_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3120 _00872_ VGND VGND VPWR VPWR net3120 sky130_fd_sc_hd__clkbuf_1
X_24019_ _03880_ _03881_ VGND VGND VPWR VPWR _03882_ sky130_fd_sc_hd__xnor2_1
X_16910_ net6407 cordic0.slte0.opA\[8\] VGND VGND VPWR VPWR _08874_ sky130_fd_sc_hd__xor2_1
Xwire3131 _11489_ VGND VGND VPWR VPWR net3131 sky130_fd_sc_hd__buf_1
Xwire3142 _11410_ VGND VGND VPWR VPWR net3142 sky130_fd_sc_hd__buf_1
Xwire3153 net3154 VGND VGND VPWR VPWR net3153 sky130_fd_sc_hd__clkbuf_2
X_17890_ net7027 net7091 VGND VGND VPWR VPWR _09741_ sky130_fd_sc_hd__or2b_1
Xwire3164 net3165 VGND VGND VPWR VPWR net3164 sky130_fd_sc_hd__buf_1
Xwire2430 _03102_ VGND VGND VPWR VPWR net2430 sky130_fd_sc_hd__buf_1
Xwire3175 _11061_ VGND VGND VPWR VPWR net3175 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire2441 net2442 VGND VGND VPWR VPWR net2441 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3186 _10973_ VGND VGND VPWR VPWR net3186 sky130_fd_sc_hd__clkbuf_2
X_16841_ _08811_ VGND VGND VPWR VPWR _00318_ sky130_fd_sc_hd__clkbuf_1
Xwire2452 net2453 VGND VGND VPWR VPWR net2452 sky130_fd_sc_hd__clkbuf_1
Xwire3197 net3198 VGND VGND VPWR VPWR net3197 sky130_fd_sc_hd__buf_1
Xwire2474 _01852_ VGND VGND VPWR VPWR net2474 sky130_fd_sc_hd__buf_1
Xwire1740 net1741 VGND VGND VPWR VPWR net1740 sky130_fd_sc_hd__clkbuf_2
Xwire2485 _12532_ VGND VGND VPWR VPWR net2485 sky130_fd_sc_hd__buf_1
X_19560_ net2513 _10938_ VGND VGND VPWR VPWR _11397_ sky130_fd_sc_hd__nand2_1
Xwire1751 _11322_ VGND VGND VPWR VPWR net1751 sky130_fd_sc_hd__buf_1
Xwire2496 _11865_ VGND VGND VPWR VPWR net2496 sky130_fd_sc_hd__clkbuf_1
X_16772_ _08775_ VGND VGND VPWR VPWR _00285_ sky130_fd_sc_hd__clkbuf_1
X_13984_ net836 _06203_ VGND VGND VPWR VPWR _06249_ sky130_fd_sc_hd__and2_1
Xwire1762 net1763 VGND VGND VPWR VPWR net1762 sky130_fd_sc_hd__buf_1
Xwire1773 _10238_ VGND VGND VPWR VPWR net1773 sky130_fd_sc_hd__buf_1
XFILLER_0_189_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18511_ net6982 net7070 net3229 VGND VGND VPWR VPWR _10360_ sky130_fd_sc_hd__or3b_1
Xwire1784 net1785 VGND VGND VPWR VPWR net1784 sky130_fd_sc_hd__buf_1
Xwire1795 _09210_ VGND VGND VPWR VPWR net1795 sky130_fd_sc_hd__buf_1
X_15723_ net1852 _07658_ _07793_ VGND VGND VPWR VPWR _07794_ sky130_fd_sc_hd__a21o_1
X_12935_ _05206_ net736 _05207_ VGND VGND VPWR VPWR _05208_ sky130_fd_sc_hd__a21o_1
X_19491_ net6085 net6048 VGND VGND VPWR VPWR _11328_ sky130_fd_sc_hd__xnor2_2
X_18442_ net7014 net7099 VGND VGND VPWR VPWR _10292_ sky130_fd_sc_hd__nand2_1
X_15654_ net2661 _07722_ _07725_ net2755 VGND VGND VPWR VPWR _07726_ sky130_fd_sc_hd__a211o_1
XFILLER_0_157_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12866_ _05137_ _05138_ net1594 net1007 VGND VGND VPWR VPWR _05139_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_158_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14605_ _06771_ _06770_ _06777_ VGND VGND VPWR VPWR _06778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18373_ net6807 net6774 VGND VGND VPWR VPWR _10224_ sky130_fd_sc_hd__xnor2_2
X_15585_ _07655_ _07656_ VGND VGND VPWR VPWR _07657_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12797_ _05068_ _05069_ VGND VGND VPWR VPWR _05070_ sky130_fd_sc_hd__nand2_1
X_17324_ _04973_ _09236_ VGND VGND VPWR VPWR _09238_ sky130_fd_sc_hd__nor2_1
XFILLER_0_173_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14536_ net5247 _06710_ net7278 VGND VGND VPWR VPWR _06715_ sky130_fd_sc_hd__o21a_1
XFILLER_0_154_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17255_ net2958 net157 net2161 net9176 VGND VGND VPWR VPWR _00353_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14467_ _06654_ VGND VGND VPWR VPWR _06655_ sky130_fd_sc_hd__buf_1
XFILLER_0_181_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16206_ net3431 net2786 VGND VGND VPWR VPWR _08271_ sky130_fd_sc_hd__nand2_1
X_13418_ _05688_ net2944 VGND VGND VPWR VPWR _05691_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17186_ net618 _09129_ _09136_ VGND VGND VPWR VPWR _09137_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_183_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14398_ _06601_ matmul0.b_in\[2\] net901 VGND VGND VPWR VPWR _06602_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_180_Right_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16137_ _08120_ _08125_ _08118_ VGND VGND VPWR VPWR _08203_ sky130_fd_sc_hd__a21o_1
X_13349_ _05618_ _05620_ net7893 _05527_ VGND VGND VPWR VPWR _05622_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_11_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16068_ _08050_ _08134_ _08049_ VGND VGND VPWR VPWR _08135_ sky130_fd_sc_hd__o21a_1
XFILLER_0_110_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15019_ net2826 _07092_ _07090_ VGND VGND VPWR VPWR _07093_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_16_Left_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19827_ _11655_ _11660_ VGND VGND VPWR VPWR _11661_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_75_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19758_ _11584_ _11592_ VGND VGND VPWR VPWR _11593_ sky130_fd_sc_hd__xor2_1
XFILLER_0_182_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18709_ _10485_ _10491_ VGND VGND VPWR VPWR _10555_ sky130_fd_sc_hd__nor2_1
X_19689_ _11517_ _11524_ VGND VGND VPWR VPWR _11525_ sky130_fd_sc_hd__xor2_1
XFILLER_0_151_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21720_ pid_d.prev_error\[5\] net5969 VGND VGND VPWR VPWR _01731_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_182_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21651_ net5688 net5566 VGND VGND VPWR VPWR _01662_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8109 net8110 VGND VGND VPWR VPWR net8109 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20602_ net3914 net1822 net1740 VGND VGND VPWR VPWR _12383_ sky130_fd_sc_hd__mux2_1
X_24370_ net1655 net1654 _04228_ VGND VGND VPWR VPWR _04229_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_25_Left_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21582_ _01591_ _01593_ VGND VGND VPWR VPWR _01594_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7408 net7409 VGND VGND VPWR VPWR net7408 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7419 matmul0.matmul_stage_inst.c\[1\] VGND VGND VPWR VPWR net7419 sky130_fd_sc_hd__clkbuf_1
X_23321_ net4887 net4760 net4771 net4864 VGND VGND VPWR VPWR _03191_ sky130_fd_sc_hd__a22o_1
X_20533_ net3193 net2079 VGND VGND VPWR VPWR _12319_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3128 net3129 VGND VGND VPWR VPWR net3128 sky130_fd_sc_hd__clkbuf_1
Xwire6707 net6708 VGND VGND VPWR VPWR net6707 sky130_fd_sc_hd__buf_1
XFILLER_0_172_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23252_ _03014_ _03024_ VGND VGND VPWR VPWR _03122_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20464_ net8044 cordic0.slte0.opA\[15\] _12249_ _12253_ _12255_ VGND VGND VPWR VPWR
+ _00498_ sky130_fd_sc_hd__o221a_1
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22203_ _02122_ _02124_ _02123_ VGND VGND VPWR VPWR _02208_ sky130_fd_sc_hd__o21a_1
Xmax_length1715 net1716 VGND VGND VPWR VPWR net1715 sky130_fd_sc_hd__buf_1
XFILLER_0_162_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23183_ net5145 net4723 _03051_ _03052_ VGND VGND VPWR VPWR _03053_ sky130_fd_sc_hd__a31o_1
X_20395_ _08835_ net1223 VGND VGND VPWR VPWR _12193_ sky130_fd_sc_hd__nand2_1
X_22134_ _02031_ _02032_ _02030_ VGND VGND VPWR VPWR _02140_ sky130_fd_sc_hd__o21ai_1
X_22065_ net1715 _01969_ VGND VGND VPWR VPWR _02072_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_34_Left_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21016_ net5556 net5910 VGND VGND VPWR VPWR _01032_ sky130_fd_sc_hd__nand2_1
Xwire1003 _05220_ VGND VGND VPWR VPWR net1003 sky130_fd_sc_hd__buf_1
Xwire1014 _04089_ VGND VGND VPWR VPWR net1014 sky130_fd_sc_hd__clkbuf_1
Xwire1025 net1026 VGND VGND VPWR VPWR net1025 sky130_fd_sc_hd__clkbuf_1
Xwire1036 net1037 VGND VGND VPWR VPWR net1036 sky130_fd_sc_hd__buf_1
X_25824_ clknet_leaf_38_clk _00697_ net8746 VGND VGND VPWR VPWR pid_q.curr_error\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xwire1047 _01829_ VGND VGND VPWR VPWR net1047 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1058 net1059 VGND VGND VPWR VPWR net1058 sky130_fd_sc_hd__buf_1
Xwire1069 _10450_ VGND VGND VPWR VPWR net1069 sky130_fd_sc_hd__buf_1
X_25755_ clknet_leaf_13_clk _00628_ net8608 VGND VGND VPWR VPWR pid_d.kp\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22967_ _02851_ VGND VGND VPWR VPWR _00650_ sky130_fd_sc_hd__clkbuf_1
X_24706_ net9055 _04530_ net1011 net1642 VGND VGND VPWR VPWR _00698_ sky130_fd_sc_hd__a22o_1
X_12720_ _04984_ _04989_ _04992_ VGND VGND VPWR VPWR _04993_ sky130_fd_sc_hd__o21a_1
X_21918_ _01832_ _01834_ _01833_ VGND VGND VPWR VPWR _01926_ sky130_fd_sc_hd__o21a_1
XFILLER_0_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25686_ clknet_leaf_3_clk _00559_ net8572 VGND VGND VPWR VPWR pid_d.curr_error\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_168_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22898_ net8899 _02791_ VGND VGND VPWR VPWR _02792_ sky130_fd_sc_hd__and2_1
X_24637_ _04474_ _04491_ VGND VGND VPWR VPWR _04492_ sky130_fd_sc_hd__xnor2_1
X_12651_ net2344 VGND VGND VPWR VPWR _04924_ sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_43_Left_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length5020 net5011 VGND VGND VPWR VPWR net5020 sky130_fd_sc_hd__buf_1
X_21849_ net1719 _01857_ VGND VGND VPWR VPWR _01858_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8537 net8844 VGND VGND VPWR VPWR net8537 sky130_fd_sc_hd__buf_1
XFILLER_0_127_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8610 net8611 VGND VGND VPWR VPWR net8610 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8621 net8620 VGND VGND VPWR VPWR net8621 sky130_fd_sc_hd__buf_2
X_12582_ net4311 pid_d.state\[0\] net4327 _04867_ VGND VGND VPWR VPWR _00015_ sky130_fd_sc_hd__a211o_1
XFILLER_0_26_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15370_ _07438_ net2824 VGND VGND VPWR VPWR _07444_ sky130_fd_sc_hd__nor2_1
Xwire8632 net8629 VGND VGND VPWR VPWR net8632 sky130_fd_sc_hd__dlymetal6s2s_1
X_24568_ net4823 net4506 VGND VGND VPWR VPWR _04424_ sky130_fd_sc_hd__nand2_1
Xwire8643 net8633 VGND VGND VPWR VPWR net8643 sky130_fd_sc_hd__buf_1
XFILLER_0_154_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length5086 net5087 VGND VGND VPWR VPWR net5086 sky130_fd_sc_hd__clkbuf_1
Xwire300 net301 VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__clkbuf_1
X_14321_ _06542_ VGND VGND VPWR VPWR _06543_ sky130_fd_sc_hd__buf_1
XFILLER_0_80_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7920 net7921 VGND VGND VPWR VPWR net7920 sky130_fd_sc_hd__clkbuf_1
X_23519_ _03386_ _03387_ net7511 VGND VGND VPWR VPWR _03388_ sky130_fd_sc_hd__o21a_1
Xwire311 net312 VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__buf_1
Xwire322 _05862_ VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__buf_1
Xwire7931 net7932 VGND VGND VPWR VPWR net7931 sky130_fd_sc_hd__buf_1
Xmax_length4363 net4365 VGND VGND VPWR VPWR net4363 sky130_fd_sc_hd__buf_1
Xwire333 net334 VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__buf_1
X_24499_ _04286_ _04305_ net1650 VGND VGND VPWR VPWR _04356_ sky130_fd_sc_hd__o21a_1
XFILLER_0_135_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7953 net7954 VGND VGND VPWR VPWR net7953 sky130_fd_sc_hd__clkbuf_1
Xwire8698 net8700 VGND VGND VPWR VPWR net8698 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire7964 net7965 VGND VGND VPWR VPWR net7964 sky130_fd_sc_hd__clkbuf_1
Xwire344 net345 VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__clkbuf_1
X_17040_ net7057 net967 _08994_ _08996_ _08999_ VGND VGND VPWR VPWR _09000_ sky130_fd_sc_hd__o311a_1
XFILLER_0_68_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14252_ net8047 net2932 VGND VGND VPWR VPWR _06507_ sky130_fd_sc_hd__nand2_1
Xwire355 net356 VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__clkbuf_1
Xwire366 _06319_ VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__buf_1
Xwire7975 net7976 VGND VGND VPWR VPWR net7975 sky130_fd_sc_hd__clkbuf_1
Xwire7986 net7987 VGND VGND VPWR VPWR net7986 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire377 net378 VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__clkbuf_1
Xwire7997 net7998 VGND VGND VPWR VPWR net7997 sky130_fd_sc_hd__clkbuf_1
Xwire388 _08090_ VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__clkbuf_1
X_13203_ net1001 VGND VGND VPWR VPWR _05476_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire399 net400 VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__buf_1
X_14183_ net7626 net1120 VGND VGND VPWR VPWR _06443_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13134_ _05342_ net2303 _05406_ VGND VGND VPWR VPWR _05407_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18991_ net6343 net6357 VGND VGND VPWR VPWR _10828_ sky130_fd_sc_hd__or2b_1
X_13065_ net7846 net2966 net2305 VGND VGND VPWR VPWR _05338_ sky130_fd_sc_hd__and3_1
X_17942_ net6912 net6851 VGND VGND VPWR VPWR _09793_ sky130_fd_sc_hd__xor2_2
XFILLER_0_178_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17873_ _09605_ _09610_ VGND VGND VPWR VPWR _09724_ sky130_fd_sc_hd__nor2_1
Xwire2260 _06841_ VGND VGND VPWR VPWR net2260 sky130_fd_sc_hd__clkbuf_1
Xwire2271 net2272 VGND VGND VPWR VPWR net2271 sky130_fd_sc_hd__clkbuf_1
X_19612_ net3136 _11448_ VGND VGND VPWR VPWR _11449_ sky130_fd_sc_hd__nor2_2
X_16824_ _08802_ VGND VGND VPWR VPWR _00310_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2282 net2283 VGND VGND VPWR VPWR net2282 sky130_fd_sc_hd__clkbuf_1
Xwire2293 _05609_ VGND VGND VPWR VPWR net2293 sky130_fd_sc_hd__buf_1
XFILLER_0_45_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1570 _05764_ VGND VGND VPWR VPWR net1570 sky130_fd_sc_hd__buf_1
X_19543_ net2106 _11379_ VGND VGND VPWR VPWR _11380_ sky130_fd_sc_hd__xnor2_2
Xwire1581 net1582 VGND VGND VPWR VPWR net1581 sky130_fd_sc_hd__clkbuf_1
X_16755_ _08766_ VGND VGND VPWR VPWR _00277_ sky130_fd_sc_hd__clkbuf_1
X_13967_ _06228_ _06231_ VGND VGND VPWR VPWR _06232_ sky130_fd_sc_hd__xnor2_2
X_15706_ _07680_ net1266 _07776_ VGND VGND VPWR VPWR _07777_ sky130_fd_sc_hd__o21ai_1
X_12918_ net2304 net2964 VGND VGND VPWR VPWR _05191_ sky130_fd_sc_hd__and2_1
X_19474_ _11266_ _11310_ VGND VGND VPWR VPWR _11311_ sky130_fd_sc_hd__nand2_1
X_16686_ _08716_ _08712_ matmul0.matmul_stage_inst.mult2\[9\] VGND VGND VPWR VPWR
+ _08717_ sky130_fd_sc_hd__o21ba_1
X_13898_ net7788 net1568 _06132_ VGND VGND VPWR VPWR _06164_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18425_ net6826 net3983 VGND VGND VPWR VPWR _10275_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15637_ net888 _07708_ VGND VGND VPWR VPWR _07709_ sky130_fd_sc_hd__xor2_1
XFILLER_0_185_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12849_ _05118_ _05121_ VGND VGND VPWR VPWR _05122_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_152_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18356_ _10171_ VGND VGND VPWR VPWR _10207_ sky130_fd_sc_hd__inv_2
X_15568_ matmul0.matmul_stage_inst.mult1\[1\] net440 net2678 VGND VGND VPWR VPWR _07641_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_185_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17307_ net7765 net7742 net1795 VGND VGND VPWR VPWR _09221_ sky130_fd_sc_hd__nor3_1
XFILLER_0_44_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14519_ net9068 net832 _06699_ net2886 VGND VGND VPWR VPWR _00108_ sky130_fd_sc_hd__a22o_1
X_18287_ _10074_ _10075_ _10137_ VGND VGND VPWR VPWR _10138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15499_ net6622 net6643 net7380 VGND VGND VPWR VPWR _07572_ sky130_fd_sc_hd__o21a_1
XFILLER_0_182_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17238_ net2957 VGND VGND VPWR VPWR _09185_ sky130_fd_sc_hd__buf_1
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17169_ _09120_ _09121_ VGND VGND VPWR VPWR _00336_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20180_ _11944_ _11974_ VGND VGND VPWR VPWR _12006_ sky130_fd_sc_hd__or2b_1
XFILLER_0_12_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23870_ net1164 _03637_ _03614_ VGND VGND VPWR VPWR _03735_ sky130_fd_sc_hd__o21a_1
Xmax_length8607 net8605 VGND VGND VPWR VPWR net8607 sky130_fd_sc_hd__buf_1
XFILLER_0_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length8618 net8619 VGND VGND VPWR VPWR net8618 sky130_fd_sc_hd__buf_1
X_22821_ pid_d.out\[0\] net5986 VGND VGND VPWR VPWR _02723_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25540_ clknet_leaf_32_clk _00420_ net8683 VGND VGND VPWR VPWR pid_q.prev_int\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_22752_ _02679_ VGND VGND VPWR VPWR _00607_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21703_ net2069 _01713_ VGND VGND VPWR VPWR _01714_ sky130_fd_sc_hd__nor2_1
X_25471_ clknet_leaf_46_clk _00351_ net8811 VGND VGND VPWR VPWR svm0.tB\[9\] sky130_fd_sc_hd__dfrtp_1
X_22683_ _02630_ VGND VGND VPWR VPWR _00587_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24422_ net2409 net2404 VGND VGND VPWR VPWR _04280_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21634_ _01644_ _01542_ pid_d.curr_int\[4\] VGND VGND VPWR VPWR _01645_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_81_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7205 net7206 VGND VGND VPWR VPWR net7205 sky130_fd_sc_hd__clkbuf_1
Xwire7216 net7217 VGND VGND VPWR VPWR net7216 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24353_ _04206_ _04211_ VGND VGND VPWR VPWR _04212_ sky130_fd_sc_hd__xor2_1
Xwire7227 net7228 VGND VGND VPWR VPWR net7227 sky130_fd_sc_hd__buf_1
X_21565_ _01466_ _01468_ _01576_ VGND VGND VPWR VPWR _01577_ sky130_fd_sc_hd__a21oi_2
Xwire7238 net7239 VGND VGND VPWR VPWR net7238 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6504 net6503 VGND VGND VPWR VPWR net6504 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_118_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23304_ _03009_ _03171_ _03172_ _03173_ VGND VGND VPWR VPWR _03174_ sky130_fd_sc_hd__a22o_1
X_20516_ _12301_ _12302_ VGND VGND VPWR VPWR _12303_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24284_ net2020 net1657 net2409 VGND VGND VPWR VPWR _04144_ sky130_fd_sc_hd__a21o_1
Xwire6526 net6527 VGND VGND VPWR VPWR net6526 sky130_fd_sc_hd__buf_1
XFILLER_0_144_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire6537 net6535 VGND VGND VPWR VPWR net6537 sky130_fd_sc_hd__buf_1
X_21496_ net5427 _01508_ _01506_ net5416 VGND VGND VPWR VPWR _01509_ sky130_fd_sc_hd__o211ai_1
Xwire6548 net6549 VGND VGND VPWR VPWR net6548 sky130_fd_sc_hd__buf_1
Xmax_length2235 _07377_ VGND VGND VPWR VPWR net2235 sky130_fd_sc_hd__buf_1
Xwire5803 net5807 VGND VGND VPWR VPWR net5803 sky130_fd_sc_hd__buf_1
XFILLER_0_133_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5814 net5815 VGND VGND VPWR VPWR net5814 sky130_fd_sc_hd__buf_1
X_23235_ net5000 net4739 VGND VGND VPWR VPWR _03105_ sky130_fd_sc_hd__nand2_1
Xwire6559 net6560 VGND VGND VPWR VPWR net6559 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_166_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5825 net5826 VGND VGND VPWR VPWR net5825 sky130_fd_sc_hd__clkbuf_1
X_20447_ _08857_ _12226_ VGND VGND VPWR VPWR _12240_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5847 net5853 VGND VGND VPWR VPWR net5847 sky130_fd_sc_hd__clkbuf_1
Xwire5858 net5859 VGND VGND VPWR VPWR net5858 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire5869 net5873 VGND VGND VPWR VPWR net5869 sky130_fd_sc_hd__buf_1
X_23166_ _03028_ _03029_ VGND VGND VPWR VPWR _03036_ sky130_fd_sc_hd__xnor2_1
X_20378_ _12174_ _12176_ net6495 VGND VGND VPWR VPWR _12177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22117_ net5692 net5481 VGND VGND VPWR VPWR _02123_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23097_ net4912 net4758 VGND VGND VPWR VPWR _02967_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22048_ net5817 net5841 net5858 VGND VGND VPWR VPWR _02055_ sky130_fd_sc_hd__and3_1
X_14870_ net7185 matmul0.matmul_stage_inst.f\[7\] net3606 VGND VGND VPWR VPWR _06953_
+ sky130_fd_sc_hd__mux2_1
X_13821_ _06064_ _06073_ _06087_ VGND VGND VPWR VPWR _06088_ sky130_fd_sc_hd__o21ai_1
X_25807_ clknet_leaf_30_clk _00680_ net8673 VGND VGND VPWR VPWR pid_q.curr_int\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23999_ _03860_ _03773_ _03861_ VGND VGND VPWR VPWR _03862_ sky130_fd_sc_hd__o21a_1
XFILLER_0_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16540_ _08597_ _08598_ net1078 VGND VGND VPWR VPWR _08599_ sky130_fd_sc_hd__mux2_1
X_13752_ _05862_ net321 net320 VGND VGND VPWR VPWR _06020_ sky130_fd_sc_hd__o21ai_1
X_25738_ clknet_leaf_13_clk _00611_ net8614 VGND VGND VPWR VPWR pid_d.ki\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12703_ net2323 net2319 VGND VGND VPWR VPWR _04976_ sky130_fd_sc_hd__nand2_1
X_16471_ _08524_ _08531_ VGND VGND VPWR VPWR _08532_ sky130_fd_sc_hd__xnor2_2
X_13683_ _05950_ _05951_ VGND VGND VPWR VPWR _05952_ sky130_fd_sc_hd__and2_1
X_25669_ clknet_leaf_5_clk _00542_ net8565 VGND VGND VPWR VPWR pid_d.prev_error\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout8334 net8339 VGND VGND VPWR VPWR net8334 sky130_fd_sc_hd__buf_1
X_18210_ net3239 net3238 _10058_ _10059_ VGND VGND VPWR VPWR _10061_ sky130_fd_sc_hd__and4_1
X_15422_ _07478_ _07495_ VGND VGND VPWR VPWR _07496_ sky130_fd_sc_hd__xor2_2
X_12634_ net2989 VGND VGND VPWR VPWR _04907_ sky130_fd_sc_hd__clkbuf_1
X_19190_ net6259 net3900 _11024_ net3877 _11026_ VGND VGND VPWR VPWR _11027_ sky130_fd_sc_hd__a221o_1
Xfanout7611 net7620 VGND VGND VPWR VPWR net7611 sky130_fd_sc_hd__buf_1
Xfanout7633 net7635 VGND VGND VPWR VPWR net7633 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_53_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18141_ _09939_ _09988_ _09989_ _09991_ net2548 VGND VGND VPWR VPWR _09992_ sky130_fd_sc_hd__o221a_1
Xwire8440 net8438 VGND VGND VPWR VPWR net8440 sky130_fd_sc_hd__buf_1
X_15353_ _07418_ _07423_ _07426_ VGND VGND VPWR VPWR _07427_ sky130_fd_sc_hd__o21ba_1
Xwire8451 net8450 VGND VGND VPWR VPWR net8451 sky130_fd_sc_hd__buf_1
X_12565_ net6748 net6598 VGND VGND VPWR VPWR _04855_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6932 net6936 VGND VGND VPWR VPWR net6932 sky130_fd_sc_hd__clkbuf_2
Xwire8473 net8474 VGND VGND VPWR VPWR net8473 sky130_fd_sc_hd__dlymetal6s2s_1
X_14304_ net6448 net6454 net6444 VGND VGND VPWR VPWR _06526_ sky130_fd_sc_hd__nor3_1
Xmax_length4171 net4172 VGND VGND VPWR VPWR net4171 sky130_fd_sc_hd__buf_1
Xwire7750 net7751 VGND VGND VPWR VPWR net7750 sky130_fd_sc_hd__clkbuf_1
X_18072_ _09917_ _09921_ _09922_ VGND VGND VPWR VPWR _09923_ sky130_fd_sc_hd__o21ai_1
Xwire7761 net7762 VGND VGND VPWR VPWR net7761 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15284_ net2839 _07045_ _07050_ _07051_ VGND VGND VPWR VPWR _07358_ sky130_fd_sc_hd__o22a_1
Xmax_length4193 net4194 VGND VGND VPWR VPWR net4193 sky130_fd_sc_hd__buf_1
Xwire7772 net7773 VGND VGND VPWR VPWR net7772 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire7783 net7785 VGND VGND VPWR VPWR net7783 sky130_fd_sc_hd__buf_1
Xwire163 net164 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_1
Xwire174 _06399_ VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__buf_1
X_17023_ net3336 _08982_ _08983_ _08981_ VGND VGND VPWR VPWR _00328_ sky130_fd_sc_hd__a2bb2o_1
Xwire7794 net7795 VGND VGND VPWR VPWR net7794 sky130_fd_sc_hd__clkbuf_1
X_14235_ net1119 _06472_ _06491_ _06470_ VGND VGND VPWR VPWR _06492_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout6998 net7002 VGND VGND VPWR VPWR net6998 sky130_fd_sc_hd__clkbuf_2
Xwire185 net186 VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_1
Xwire196 net197 VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2780 net2781 VGND VGND VPWR VPWR net2780 sky130_fd_sc_hd__buf_1
XFILLER_0_141_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14166_ _06368_ VGND VGND VPWR VPWR _06427_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13117_ _05388_ _05389_ VGND VGND VPWR VPWR _05390_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14097_ net282 net319 _06359_ _06280_ VGND VGND VPWR VPWR _06360_ sky130_fd_sc_hd__a31o_1
X_18974_ _10810_ VGND VGND VPWR VPWR _10811_ sky130_fd_sc_hd__clkbuf_2
X_13048_ net789 _05004_ VGND VGND VPWR VPWR _05321_ sky130_fd_sc_hd__nor2_1
X_17925_ _09734_ _09774_ _09775_ VGND VGND VPWR VPWR _09776_ sky130_fd_sc_hd__o21ai_1
X_17856_ net7029 net7124 net7140 VGND VGND VPWR VPWR _09707_ sky130_fd_sc_hd__or3b_1
XFILLER_0_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2090 _12204_ VGND VGND VPWR VPWR net2090 sky130_fd_sc_hd__clkbuf_1
X_16807_ net8975 matmul0.cos\[6\] net3368 VGND VGND VPWR VPWR _08794_ sky130_fd_sc_hd__mux2_1
X_17787_ net4043 net3993 _09635_ net3992 _09637_ VGND VGND VPWR VPWR _09638_ sky130_fd_sc_hd__a221o_1
XFILLER_0_191_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14999_ _07072_ VGND VGND VPWR VPWR _07073_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19526_ _11353_ _11362_ VGND VGND VPWR VPWR _11363_ sky130_fd_sc_hd__xnor2_2
X_16738_ _08757_ VGND VGND VPWR VPWR _00269_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19457_ _11291_ net3158 VGND VGND VPWR VPWR _11294_ sky130_fd_sc_hd__xor2_1
X_16669_ matmul0.alpha_pass\[7\] net823 net6563 VGND VGND VPWR VPWR _08703_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18408_ _10257_ _10258_ VGND VGND VPWR VPWR _10259_ sky130_fd_sc_hd__and2b_1
X_19388_ _11025_ _11180_ VGND VGND VPWR VPWR _11225_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18339_ net1074 _10128_ _10127_ VGND VGND VPWR VPWR _10190_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_84_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout8890 net8900 VGND VGND VPWR VPWR net8890 sky130_fd_sc_hd__buf_1
XFILLER_0_16_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21350_ _01360_ _01363_ VGND VGND VPWR VPWR _01364_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_170_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20301_ net6499 net6471 VGND VGND VPWR VPWR _12106_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21281_ _01294_ _01295_ VGND VGND VPWR VPWR _01296_ sky130_fd_sc_hd__xor2_1
Xwire4409 net4410 VGND VGND VPWR VPWR net4409 sky130_fd_sc_hd__clkbuf_1
X_23020_ net4949 net4740 VGND VGND VPWR VPWR _02890_ sky130_fd_sc_hd__nand2_2
XFILLER_0_13_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20232_ net10 net11 _12043_ VGND VGND VPWR VPWR _12050_ sky130_fd_sc_hd__and3_1
Xwire3708 net3709 VGND VGND VPWR VPWR net3708 sky130_fd_sc_hd__clkbuf_1
Xwire3719 net3720 VGND VGND VPWR VPWR net3719 sky130_fd_sc_hd__buf_1
X_20163_ _11988_ _11989_ net1439 VGND VGND VPWR VPWR _11990_ sky130_fd_sc_hd__a21oi_1
X_24971_ _04740_ VGND VGND VPWR VPWR _00765_ sky130_fd_sc_hd__clkbuf_1
X_20094_ _11913_ _11922_ VGND VGND VPWR VPWR _11923_ sky130_fd_sc_hd__or2_1
XFILLER_0_196_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23922_ _03782_ _03785_ VGND VGND VPWR VPWR _03786_ sky130_fd_sc_hd__xnor2_1
X_23853_ net4617 net4891 VGND VGND VPWR VPWR _03718_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22804_ pid_d.kp\[14\] _02690_ net2036 VGND VGND VPWR VPWR _02710_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23784_ net1163 _03649_ VGND VGND VPWR VPWR _03650_ sky130_fd_sc_hd__xnor2_2
X_20996_ _01009_ _01010_ net1732 VGND VGND VPWR VPWR _01012_ sky130_fd_sc_hd__a21o_1
XFILLER_0_177_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25523_ clknet_leaf_48_clk _00403_ net8756 VGND VGND VPWR VPWR svm0.counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_22735_ net3718 net106 VGND VGND VPWR VPWR _02668_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25454_ clknet_leaf_112_clk _00337_ net8362 VGND VGND VPWR VPWR cordic0.vec\[1\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_22666_ net5650 net3085 net178 net8888 VGND VGND VPWR VPWR _00582_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24405_ _04261_ _04262_ VGND VGND VPWR VPWR _04263_ sky130_fd_sc_hd__xnor2_1
Xwire7002 net7003 VGND VGND VPWR VPWR net7002 sky130_fd_sc_hd__buf_1
Xfanout6206 net6213 VGND VGND VPWR VPWR net6206 sky130_fd_sc_hd__buf_1
X_21617_ _01447_ _01519_ _01442_ VGND VGND VPWR VPWR _01629_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_109_Right_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7013 net7012 VGND VGND VPWR VPWR net7013 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_47_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25385_ clknet_leaf_73_clk _00268_ net8474 VGND VGND VPWR VPWR matmul0.b\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_164_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6228 net6237 VGND VGND VPWR VPWR net6228 sky130_fd_sc_hd__buf_1
Xwire7024 net7025 VGND VGND VPWR VPWR net7024 sky130_fd_sc_hd__clkbuf_1
X_22597_ _02573_ VGND VGND VPWR VPWR _00558_ sky130_fd_sc_hd__clkbuf_1
Xwire7035 net7038 VGND VGND VPWR VPWR net7035 sky130_fd_sc_hd__buf_1
XFILLER_0_62_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout5505 net5519 VGND VGND VPWR VPWR net5505 sky130_fd_sc_hd__buf_1
Xwire7046 net7043 VGND VGND VPWR VPWR net7046 sky130_fd_sc_hd__buf_1
X_24336_ net634 net633 _04194_ _04105_ VGND VGND VPWR VPWR _04195_ sky130_fd_sc_hd__a211o_1
Xwire6312 net6311 VGND VGND VPWR VPWR net6312 sky130_fd_sc_hd__buf_2
XFILLER_0_90_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21548_ _01558_ _01559_ VGND VGND VPWR VPWR _01560_ sky130_fd_sc_hd__xnor2_1
Xwire6323 net6320 VGND VGND VPWR VPWR net6323 sky130_fd_sc_hd__buf_1
XFILLER_0_105_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire7068 net7069 VGND VGND VPWR VPWR net7068 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7079 net7073 VGND VGND VPWR VPWR net7079 sky130_fd_sc_hd__buf_1
XFILLER_0_105_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6345 net6346 VGND VGND VPWR VPWR net6345 sky130_fd_sc_hd__clkbuf_1
Xmax_length2043 net2044 VGND VGND VPWR VPWR net2043 sky130_fd_sc_hd__buf_1
Xfanout4826 net4832 VGND VGND VPWR VPWR net4826 sky130_fd_sc_hd__buf_1
X_24267_ net4589 net4803 VGND VGND VPWR VPWR _04127_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5622 net5620 VGND VGND VPWR VPWR net5622 sky130_fd_sc_hd__clkbuf_1
X_21479_ net5920 net5400 VGND VGND VPWR VPWR _01492_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5633 net5630 VGND VGND VPWR VPWR net5633 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6378 net6377 VGND VGND VPWR VPWR net6378 sky130_fd_sc_hd__buf_1
X_14020_ _06234_ _06242_ _06283_ VGND VGND VPWR VPWR _06284_ sky130_fd_sc_hd__a21o_1
Xwire6389 cordic0.domain\[0\] VGND VGND VPWR VPWR net6389 sky130_fd_sc_hd__clkbuf_1
X_23218_ _03060_ _03086_ VGND VGND VPWR VPWR _03088_ sky130_fd_sc_hd__nand2_1
Xwire4910 net4903 VGND VGND VPWR VPWR net4910 sky130_fd_sc_hd__clkbuf_1
Xwire5655 net5657 VGND VGND VPWR VPWR net5655 sky130_fd_sc_hd__clkbuf_1
Xwire4921 net4922 VGND VGND VPWR VPWR net4921 sky130_fd_sc_hd__clkbuf_1
Xwire5666 net5667 VGND VGND VPWR VPWR net5666 sky130_fd_sc_hd__clkbuf_1
Xwire4932 net4923 VGND VGND VPWR VPWR net4932 sky130_fd_sc_hd__clkbuf_1
X_24198_ _03986_ _03988_ _03987_ VGND VGND VPWR VPWR _04059_ sky130_fd_sc_hd__o21ai_1
Xwire5677 net5678 VGND VGND VPWR VPWR net5677 sky130_fd_sc_hd__clkbuf_1
Xmax_length1375 net1376 VGND VGND VPWR VPWR net1375 sky130_fd_sc_hd__clkbuf_1
Xwire4954 net4955 VGND VGND VPWR VPWR net4954 sky130_fd_sc_hd__clkbuf_1
Xwire5699 net5700 VGND VGND VPWR VPWR net5699 sky130_fd_sc_hd__clkbuf_1
X_23149_ _03015_ _03016_ _03018_ VGND VGND VPWR VPWR _03019_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_105_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4976 net4965 VGND VGND VPWR VPWR net4976 sky130_fd_sc_hd__buf_1
Xwire4987 net4980 VGND VGND VPWR VPWR net4987 sky130_fd_sc_hd__buf_1
Xwire4998 net4996 VGND VGND VPWR VPWR net4998 sky130_fd_sc_hd__buf_1
XFILLER_0_101_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15971_ net2649 net2626 VGND VGND VPWR VPWR _08039_ sky130_fd_sc_hd__nor2_1
XFILLER_0_175_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17710_ pid_q.prev_int\[1\] net1218 net1452 net5182 VGND VGND VPWR VPWR _00415_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14922_ net4192 net4187 net4182 net4180 VGND VGND VPWR VPWR _06996_ sky130_fd_sc_hd__o22a_1
X_18690_ _10534_ _10535_ VGND VGND VPWR VPWR _10536_ sky130_fd_sc_hd__xnor2_1
Xhold60 pid_d.curr_error\[9\] VGND VGND VPWR VPWR net9013 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 matmul0.matmul_stage_inst.a\[13\] VGND VGND VPWR VPWR net9024 sky130_fd_sc_hd__dlygate4sd3_1
X_17641_ svm0.tA\[14\] net6688 VGND VGND VPWR VPWR _09521_ sky130_fd_sc_hd__and2b_1
XFILLER_0_26_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold82 pid_d.curr_int\[8\] VGND VGND VPWR VPWR net9035 sky130_fd_sc_hd__dlygate4sd3_1
X_14853_ matmul0.a\[15\] matmul0.matmul_stage_inst.e\[15\] net3607 VGND VGND VPWR
+ VPWR _06944_ sky130_fd_sc_hd__mux2_1
Xhold93 cordic0.cos\[12\] VGND VGND VPWR VPWR net9046 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13804_ net996 _06071_ VGND VGND VPWR VPWR _06072_ sky130_fd_sc_hd__xor2_1
X_17572_ _09452_ _09453_ VGND VGND VPWR VPWR _09454_ sky130_fd_sc_hd__and2b_1
X_14784_ _06907_ VGND VGND VPWR VPWR _00165_ sky130_fd_sc_hd__clkbuf_1
X_19311_ _10985_ _11147_ _10912_ _11051_ VGND VGND VPWR VPWR _11148_ sky130_fd_sc_hd__a22o_1
X_16523_ _08581_ _08582_ VGND VGND VPWR VPWR _08583_ sky130_fd_sc_hd__or2b_1
X_13735_ _05867_ net451 VGND VGND VPWR VPWR _06004_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19242_ net3908 _10802_ _11074_ _11078_ VGND VGND VPWR VPWR _11079_ sky130_fd_sc_hd__o22a_1
Xfanout8120 net6 VGND VGND VPWR VPWR net8120 sky130_fd_sc_hd__clkbuf_2
X_16454_ _08511_ _08514_ VGND VGND VPWR VPWR _08515_ sky130_fd_sc_hd__xnor2_1
X_13666_ net322 _05935_ VGND VGND VPWR VPWR _05936_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15405_ net3584 net3577 net4098 net4096 VGND VGND VPWR VPWR _07479_ sky130_fd_sc_hd__o22a_1
X_12617_ _04889_ VGND VGND VPWR VPWR _04890_ sky130_fd_sc_hd__clkbuf_1
X_19173_ net1426 _11009_ VGND VGND VPWR VPWR _11010_ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16385_ net1248 _08400_ _08399_ VGND VGND VPWR VPWR _08447_ sky130_fd_sc_hd__a21bo_1
X_13597_ _05863_ _05865_ VGND VGND VPWR VPWR _05867_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8270 net25 VGND VGND VPWR VPWR net8270 sky130_fd_sc_hd__clkbuf_1
X_18124_ net3942 _09974_ net7135 VGND VGND VPWR VPWR _09975_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8281 net8282 VGND VGND VPWR VPWR net8281 sky130_fd_sc_hd__clkbuf_1
X_15336_ net1280 _07406_ _07408_ _07073_ _07409_ VGND VGND VPWR VPWR _07410_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_170_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout7496 net7508 VGND VGND VPWR VPWR net7496 sky130_fd_sc_hd__buf_1
Xwire8292 net8293 VGND VGND VPWR VPWR net8292 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire7580 matmul0.a_in\[15\] VGND VGND VPWR VPWR net7580 sky130_fd_sc_hd__buf_1
X_18055_ net3348 net3264 net3994 _08966_ VGND VGND VPWR VPWR _09906_ sky130_fd_sc_hd__a211o_1
Xwire7591 matmul0.a_in\[12\] VGND VGND VPWR VPWR net7591 sky130_fd_sc_hd__clkbuf_1
X_15267_ _07219_ _07265_ _07336_ _07340_ VGND VGND VPWR VPWR _07341_ sky130_fd_sc_hd__a22oi_2
XANTENNA_2 net3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout6795 net6802 VGND VGND VPWR VPWR net6795 sky130_fd_sc_hd__buf_1
XFILLER_0_124_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17006_ net4044 VGND VGND VPWR VPWR _08967_ sky130_fd_sc_hd__buf_1
X_14218_ _06466_ _06475_ VGND VGND VPWR VPWR _06477_ sky130_fd_sc_hd__or2_1
Xwire6890 net6891 VGND VGND VPWR VPWR net6890 sky130_fd_sc_hd__buf_1
X_15198_ net3583 net3581 net4169 net4164 VGND VGND VPWR VPWR _07272_ sky130_fd_sc_hd__o22a_1
XFILLER_0_22_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14149_ net1560 _06382_ net7603 net1124 VGND VGND VPWR VPWR _06410_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_6_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18957_ net6318 net6343 VGND VGND VPWR VPWR _10794_ sky130_fd_sc_hd__nand2_1
X_17908_ _09751_ _09755_ VGND VGND VPWR VPWR _09759_ sky130_fd_sc_hd__nand2_1
X_18888_ net6376 _10729_ VGND VGND VPWR VPWR _10730_ sky130_fd_sc_hd__nand2_1
XFILLER_0_174_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17839_ net7020 _09689_ VGND VGND VPWR VPWR _09690_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_178_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20850_ _12526_ _12528_ VGND VGND VPWR VPWR _00866_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19509_ net3161 _11275_ _11344_ _11345_ VGND VGND VPWR VPWR _11346_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_53_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20781_ _12548_ _12551_ VGND VGND VPWR VPWR _12552_ sky130_fd_sc_hd__xnor2_2
Xmax_length5619 net5617 VGND VGND VPWR VPWR net5619 sky130_fd_sc_hd__buf_1
XFILLER_0_53_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22520_ net3105 VGND VGND VPWR VPWR _02520_ sky130_fd_sc_hd__buf_1
XFILLER_0_14_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22451_ _02451_ _02452_ VGND VGND VPWR VPWR _02453_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_162_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21402_ net3118 _01414_ _01415_ _01304_ VGND VGND VPWR VPWR _01416_ sky130_fd_sc_hd__o22a_1
XFILLER_0_161_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25170_ clknet_leaf_54_clk _00059_ net8730 VGND VGND VPWR VPWR svm0.periodTop\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_22382_ _02380_ _02384_ VGND VGND VPWR VPWR _02385_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24121_ _03981_ _03982_ VGND VGND VPWR VPWR _03983_ sky130_fd_sc_hd__xnor2_2
X_21333_ _01343_ _01346_ VGND VGND VPWR VPWR _01347_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4206 net4207 VGND VGND VPWR VPWR net4206 sky130_fd_sc_hd__dlymetal6s2s_1
X_24052_ _03914_ VGND VGND VPWR VPWR _03915_ sky130_fd_sc_hd__inv_2
Xwire4217 net4218 VGND VGND VPWR VPWR net4217 sky130_fd_sc_hd__clkbuf_1
X_21264_ net5778 net5543 VGND VGND VPWR VPWR _01279_ sky130_fd_sc_hd__nand2_1
Xwire4228 net4229 VGND VGND VPWR VPWR net4228 sky130_fd_sc_hd__clkbuf_1
Xwire4239 net4240 VGND VGND VPWR VPWR net4239 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23003_ net5044 net4654 VGND VGND VPWR VPWR _02873_ sky130_fd_sc_hd__nand2_1
X_20215_ net8953 net8119 net8120 VGND VGND VPWR VPWR _12037_ sky130_fd_sc_hd__a21oi_1
Xwire3505 net3508 VGND VGND VPWR VPWR net3505 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_8_Left_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire3516 net3517 VGND VGND VPWR VPWR net3516 sky130_fd_sc_hd__buf_1
X_21195_ _01160_ _01188_ _01194_ VGND VGND VPWR VPWR _01211_ sky130_fd_sc_hd__and3_1
Xwire3527 _07062_ VGND VGND VPWR VPWR net3527 sky130_fd_sc_hd__buf_1
Xwire3538 _07055_ VGND VGND VPWR VPWR net3538 sky130_fd_sc_hd__clkbuf_1
Xwire2804 net2805 VGND VGND VPWR VPWR net2804 sky130_fd_sc_hd__buf_1
XFILLER_0_60_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3549 _07044_ VGND VGND VPWR VPWR net3549 sky130_fd_sc_hd__buf_1
X_20146_ net6027 _11942_ _11972_ net6078 VGND VGND VPWR VPWR _11973_ sky130_fd_sc_hd__a22o_1
Xwire2815 net2816 VGND VGND VPWR VPWR net2815 sky130_fd_sc_hd__clkbuf_2
Xwire2837 net2838 VGND VGND VPWR VPWR net2837 sky130_fd_sc_hd__buf_1
Xwire2848 _07012_ VGND VGND VPWR VPWR net2848 sky130_fd_sc_hd__buf_1
Xwire2859 _06869_ VGND VGND VPWR VPWR net2859 sky130_fd_sc_hd__buf_1
X_24954_ net8871 net135 VGND VGND VPWR VPWR _04730_ sky130_fd_sc_hd__and2b_1
X_20077_ _11850_ _11868_ _11905_ VGND VGND VPWR VPWR _11906_ sky130_fd_sc_hd__o21a_1
X_23905_ pid_q.curr_int\[5\] net3061 net2027 _03769_ VGND VGND VPWR VPWR _00670_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24885_ _04681_ VGND VGND VPWR VPWR _00738_ sky130_fd_sc_hd__clkbuf_1
X_23836_ net5121 net5095 VGND VGND VPWR VPWR _03701_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23767_ _03493_ net2413 _03632_ VGND VGND VPWR VPWR _03633_ sky130_fd_sc_hd__a21o_1
XFILLER_0_196_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20979_ net2076 _00994_ VGND VGND VPWR VPWR _00995_ sky130_fd_sc_hd__or2_1
XFILLER_0_170_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25506_ clknet_leaf_39_clk _00386_ net8770 VGND VGND VPWR VPWR svm0.delta\[11\] sky130_fd_sc_hd__dfrtp_1
X_13520_ _05701_ _05702_ _05790_ VGND VGND VPWR VPWR _05791_ sky130_fd_sc_hd__a21o_1
Xmax_length6865 net6861 VGND VGND VPWR VPWR net6865 sky130_fd_sc_hd__clkbuf_1
X_22718_ net8108 VGND VGND VPWR VPWR _02654_ sky130_fd_sc_hd__inv_2
X_23698_ net639 _03564_ VGND VGND VPWR VPWR _03565_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13451_ net915 net913 VGND VGND VPWR VPWR _05724_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25437_ clknet_leaf_98_clk _00320_ net8384 VGND VGND VPWR VPWR matmul0.sin\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_125_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout6003 net6014 VGND VGND VPWR VPWR net6003 sky130_fd_sc_hd__buf_1
X_22649_ net700 net3077 net1388 _02609_ net8889 VGND VGND VPWR VPWR _00574_ sky130_fd_sc_hd__o311a_1
Xfanout6014 cordic0.vec\[0\]\[17\] VGND VGND VPWR VPWR net6014 sky130_fd_sc_hd__buf_1
XFILLER_0_152_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16170_ _08234_ _08235_ VGND VGND VPWR VPWR _08236_ sky130_fd_sc_hd__xnor2_1
X_13382_ _05567_ _05568_ _05571_ _05486_ _05654_ VGND VGND VPWR VPWR _05655_ sky130_fd_sc_hd__a221o_1
XFILLER_0_134_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6047 net6053 VGND VGND VPWR VPWR net6047 sky130_fd_sc_hd__buf_1
X_25368_ clknet_leaf_81_clk _00251_ net8498 VGND VGND VPWR VPWR matmul0.alpha_pass\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout6058 net6076 VGND VGND VPWR VPWR net6058 sky130_fd_sc_hd__buf_1
XFILLER_0_106_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6120 net6121 VGND VGND VPWR VPWR net6120 sky130_fd_sc_hd__clkbuf_1
X_15121_ net4162 net4158 net4221 net4219 VGND VGND VPWR VPWR _07195_ sky130_fd_sc_hd__o22a_1
XFILLER_0_180_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24319_ _04178_ _04111_ pid_q.prev_error\[9\] VGND VGND VPWR VPWR _04179_ sky130_fd_sc_hd__o21ba_1
Xwire6142 net6143 VGND VGND VPWR VPWR net6142 sky130_fd_sc_hd__buf_1
X_25299_ clknet_leaf_88_clk _00182_ net8444 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.a\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout4623 net4633 VGND VGND VPWR VPWR net4623 sky130_fd_sc_hd__buf_1
Xwire5441 net5442 VGND VGND VPWR VPWR net5441 sky130_fd_sc_hd__clkbuf_1
Xwire6186 net6187 VGND VGND VPWR VPWR net6186 sky130_fd_sc_hd__buf_1
XFILLER_0_32_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15052_ net6629 matmul0.matmul_stage_inst.d\[0\] matmul0.matmul_stage_inst.a\[0\]
+ net6582 VGND VGND VPWR VPWR _07126_ sky130_fd_sc_hd__a22o_1
Xwire5452 pid_d.mult0.a\[12\] VGND VGND VPWR VPWR net5452 sky130_fd_sc_hd__buf_1
XFILLER_0_10_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout4656 pid_q.mult0.a\[6\] VGND VGND VPWR VPWR net4656 sky130_fd_sc_hd__clkbuf_1
Xwire5463 net5464 VGND VGND VPWR VPWR net5463 sky130_fd_sc_hd__clkbuf_1
X_14003_ _06162_ _06266_ _06267_ VGND VGND VPWR VPWR _06268_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5474 net5475 VGND VGND VPWR VPWR net5474 sky130_fd_sc_hd__clkbuf_1
Xwire5485 net5486 VGND VGND VPWR VPWR net5485 sky130_fd_sc_hd__buf_1
Xwire4751 net4752 VGND VGND VPWR VPWR net4751 sky130_fd_sc_hd__clkbuf_1
X_19860_ net6066 net3201 _10790_ VGND VGND VPWR VPWR _11693_ sky130_fd_sc_hd__a21o_1
Xwire4762 net4763 VGND VGND VPWR VPWR net4762 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4784 net4785 VGND VGND VPWR VPWR net4784 sky130_fd_sc_hd__buf_1
X_18811_ _10652_ _10654_ VGND VGND VPWR VPWR _10655_ sky130_fd_sc_hd__xor2_1
Xwire4795 net4796 VGND VGND VPWR VPWR net4795 sky130_fd_sc_hd__buf_1
X_19791_ net6088 net3141 net2100 VGND VGND VPWR VPWR _11625_ sky130_fd_sc_hd__a21o_1
X_15954_ _08020_ _08021_ VGND VGND VPWR VPWR _08022_ sky130_fd_sc_hd__xnor2_1
X_18742_ net6813 net6796 VGND VGND VPWR VPWR _10587_ sky130_fd_sc_hd__nor2_1
X_14905_ net3598 _06978_ VGND VGND VPWR VPWR _06979_ sky130_fd_sc_hd__xnor2_1
X_18673_ net1431 _10483_ net1433 VGND VGND VPWR VPWR _10519_ sky130_fd_sc_hd__o21a_1
X_15885_ net2737 net3395 VGND VGND VPWR VPWR _07954_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17624_ _09451_ svm0.tB\[2\] _09504_ _09500_ VGND VGND VPWR VPWR _09505_ sky130_fd_sc_hd__o22a_1
XFILLER_0_144_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14836_ matmul0.a\[7\] matmul0.matmul_stage_inst.e\[7\] net3611 VGND VGND VPWR VPWR
+ _06935_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17555_ net4009 svm0.tC\[4\] svm0.tC\[3\] net4019 VGND VGND VPWR VPWR _09437_ sky130_fd_sc_hd__o22a_1
XFILLER_0_169_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14767_ _06850_ _06894_ VGND VGND VPWR VPWR _06895_ sky130_fd_sc_hd__nand2_1
XFILLER_0_187_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16506_ _08561_ net1244 net2784 VGND VGND VPWR VPWR _08566_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13718_ _05882_ _05884_ _05986_ VGND VGND VPWR VPWR _05987_ sky130_fd_sc_hd__o21a_1
X_17486_ net6717 VGND VGND VPWR VPWR _09376_ sky130_fd_sc_hd__inv_2
XFILLER_0_184_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14698_ net7152 _06843_ VGND VGND VPWR VPWR _06844_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19225_ net2519 _11048_ net3175 VGND VGND VPWR VPWR _11062_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16437_ net723 _08478_ VGND VGND VPWR VPWR _08498_ sky130_fd_sc_hd__or2_1
X_13649_ _05895_ _05918_ VGND VGND VPWR VPWR _05919_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19156_ _10988_ net2520 VGND VGND VPWR VPWR _10993_ sky130_fd_sc_hd__xor2_1
X_16368_ net490 _08430_ VGND VGND VPWR VPWR _08431_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18107_ _09957_ VGND VGND VPWR VPWR _09958_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15319_ _06996_ _07001_ _07004_ VGND VGND VPWR VPWR _07393_ sky130_fd_sc_hd__a21o_1
X_19087_ net3892 _10829_ net6268 VGND VGND VPWR VPWR _10924_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16299_ _08360_ _08362_ _08245_ VGND VGND VPWR VPWR _08363_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_120_clk clknet_4_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_120_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_2_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18038_ net7050 net7004 VGND VGND VPWR VPWR _09889_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20000_ _11826_ _11829_ _11830_ net3860 VGND VGND VPWR VPWR _11831_ sky130_fd_sc_hd__a211o_1
XFILLER_0_185_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19989_ _11774_ _11776_ VGND VGND VPWR VPWR _11820_ sky130_fd_sc_hd__nor2_1
XFILLER_0_158_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21951_ net5812 _01957_ _01958_ VGND VGND VPWR VPWR _01959_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_20_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20902_ net3830 net3840 VGND VGND VPWR VPWR _00918_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24670_ net9145 net1376 _04517_ VGND VGND VPWR VPWR _00687_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21882_ _01799_ net1046 VGND VGND VPWR VPWR _01891_ sky130_fd_sc_hd__xnor2_1
X_23621_ _03465_ _03463_ _03487_ VGND VGND VPWR VPWR _03488_ sky130_fd_sc_hd__a21oi_1
Xmax_length6117 net6113 VGND VGND VPWR VPWR net6117 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_179_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20833_ net2483 _00848_ VGND VGND VPWR VPWR _00849_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_194_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23552_ _03417_ _03419_ VGND VGND VPWR VPWR _03420_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_194_Right_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20764_ net2486 _12533_ _12534_ VGND VGND VPWR VPWR _12535_ sky130_fd_sc_hd__o21a_1
XFILLER_0_193_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22503_ _02438_ _02501_ _02499_ VGND VGND VPWR VPWR _02504_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23483_ net4702 net4900 VGND VGND VPWR VPWR _03352_ sky130_fd_sc_hd__nand2_1
X_20695_ net6058 net1496 _12468_ VGND VGND VPWR VPWR _12470_ sky130_fd_sc_hd__and3_1
XFILLER_0_147_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire707 _12393_ VGND VGND VPWR VPWR net707 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire718 net719 VGND VGND VPWR VPWR net718 sky130_fd_sc_hd__clkbuf_1
X_25222_ clknet_leaf_59_clk _00111_ net8693 VGND VGND VPWR VPWR svm0.vC\[10\] sky130_fd_sc_hd__dfrtp_1
Xwire729 net730 VGND VGND VPWR VPWR net729 sky130_fd_sc_hd__clkbuf_1
X_22434_ net5377 _02434_ _02435_ VGND VGND VPWR VPWR _02436_ sky130_fd_sc_hd__and3_1
XFILLER_0_190_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_99_Left_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25153_ clknet_leaf_41_clk _00042_ net8767 VGND VGND VPWR VPWR pid_q.target\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22365_ _02283_ _02302_ net1702 VGND VGND VPWR VPWR _02368_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_143_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_111_clk clknet_4_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_111_clk
+ sky130_fd_sc_hd__clkbuf_16
X_24104_ net4970 net4501 VGND VGND VPWR VPWR _03966_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21316_ _01254_ _01330_ VGND VGND VPWR VPWR _01331_ sky130_fd_sc_hd__xnor2_1
X_22296_ net5765 net5780 net5800 VGND VGND VPWR VPWR _02300_ sky130_fd_sc_hd__and3_1
X_25084_ net7499 net2396 VGND VGND VPWR VPWR _04829_ sky130_fd_sc_hd__nand2_1
Xwire4014 _09291_ VGND VGND VPWR VPWR net4014 sky130_fd_sc_hd__buf_1
Xwire4025 net4026 VGND VGND VPWR VPWR net4025 sky130_fd_sc_hd__buf_1
Xwire4036 _09156_ VGND VGND VPWR VPWR net4036 sky130_fd_sc_hd__buf_1
X_24035_ _03782_ _03784_ _03783_ VGND VGND VPWR VPWR _03898_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_131_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3302 net3303 VGND VGND VPWR VPWR net3302 sky130_fd_sc_hd__clkbuf_1
X_21247_ _00826_ _00827_ _00828_ VGND VGND VPWR VPWR _01262_ sky130_fd_sc_hd__o21ai_1
Xwire3313 net3314 VGND VGND VPWR VPWR net3313 sky130_fd_sc_hd__clkbuf_2
Xwire3324 _09023_ VGND VGND VPWR VPWR net3324 sky130_fd_sc_hd__buf_1
Xwire4069 net4070 VGND VGND VPWR VPWR net4069 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3335 _08969_ VGND VGND VPWR VPWR net3335 sky130_fd_sc_hd__clkbuf_2
Xwire3346 net3348 VGND VGND VPWR VPWR net3346 sky130_fd_sc_hd__buf_1
X_21178_ net5619 net5909 _01192_ _01193_ VGND VGND VPWR VPWR _01194_ sky130_fd_sc_hd__a31o_1
Xwire2612 _08849_ VGND VGND VPWR VPWR net2612 sky130_fd_sc_hd__buf_1
Xwire3357 net3358 VGND VGND VPWR VPWR net3357 sky130_fd_sc_hd__clkbuf_1
Xwire3368 _08792_ VGND VGND VPWR VPWR net3368 sky130_fd_sc_hd__clkbuf_2
Xwire2623 _08040_ VGND VGND VPWR VPWR net2623 sky130_fd_sc_hd__buf_1
Xwire3379 _08770_ VGND VGND VPWR VPWR net3379 sky130_fd_sc_hd__buf_1
Xwire2645 net2646 VGND VGND VPWR VPWR net2645 sky130_fd_sc_hd__buf_1
Xwire1900 _07058_ VGND VGND VPWR VPWR net1900 sky130_fd_sc_hd__clkbuf_1
X_20129_ _11934_ _11956_ VGND VGND VPWR VPWR _11957_ sky130_fd_sc_hd__xnor2_1
Xwire1911 net1912 VGND VGND VPWR VPWR net1911 sky130_fd_sc_hd__clkbuf_1
Xwire2656 net2657 VGND VGND VPWR VPWR net2656 sky130_fd_sc_hd__buf_1
Xwire1922 _06508_ VGND VGND VPWR VPWR net1922 sky130_fd_sc_hd__buf_1
Xwire2667 net2668 VGND VGND VPWR VPWR net2667 sky130_fd_sc_hd__clkbuf_1
Xwire1933 net1934 VGND VGND VPWR VPWR net1933 sky130_fd_sc_hd__buf_1
Xwire2678 _07560_ VGND VGND VPWR VPWR net2678 sky130_fd_sc_hd__buf_1
Xwire1944 _05608_ VGND VGND VPWR VPWR net1944 sky130_fd_sc_hd__clkbuf_1
Xwire2689 _07508_ VGND VGND VPWR VPWR net2689 sky130_fd_sc_hd__buf_1
X_24937_ pid_q.ki\[8\] _04718_ net1361 VGND VGND VPWR VPWR _04719_ sky130_fd_sc_hd__mux2_1
Xwire1955 _05131_ VGND VGND VPWR VPWR net1955 sky130_fd_sc_hd__buf_1
X_12951_ _05010_ _05223_ VGND VGND VPWR VPWR _05224_ sky130_fd_sc_hd__xnor2_1
Xwire1966 _04965_ VGND VGND VPWR VPWR net1966 sky130_fd_sc_hd__clkbuf_1
Xwire1977 net1978 VGND VGND VPWR VPWR net1977 sky130_fd_sc_hd__clkbuf_1
Xwire1988 net1989 VGND VGND VPWR VPWR net1988 sky130_fd_sc_hd__buf_1
Xwire1999 _04665_ VGND VGND VPWR VPWR net1999 sky130_fd_sc_hd__clkbuf_1
X_15670_ _07741_ VGND VGND VPWR VPWR _00217_ sky130_fd_sc_hd__clkbuf_1
X_24868_ pid_q.ki\[4\] net2398 _00008_ pid_q.kp\[4\] VGND VGND VPWR VPWR _04670_ sky130_fd_sc_hd__a22o_1
X_12882_ net7874 net1958 VGND VGND VPWR VPWR _05155_ sky130_fd_sc_hd__nand2_1
X_14621_ _06791_ VGND VGND VPWR VPWR _00118_ sky130_fd_sc_hd__clkbuf_1
X_23819_ _03682_ _03683_ VGND VGND VPWR VPWR _03684_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_157_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_length7352 net7353 VGND VGND VPWR VPWR net7352 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24799_ net7961 _04623_ VGND VGND VPWR VPWR _04624_ sky130_fd_sc_hd__xor2_1
Xmax_length7374 matmul0.alpha_pass\[0\] VGND VGND VPWR VPWR net7374 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17340_ _09251_ _09252_ _09213_ VGND VGND VPWR VPWR _09254_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14552_ net7278 _06727_ _06729_ VGND VGND VPWR VPWR _06730_ sky130_fd_sc_hd__o21a_2
XFILLER_0_83_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_161_Right_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13503_ svm0.state\[1\] svm0.state\[0\] VGND VGND VPWR VPWR _05776_ sky130_fd_sc_hd__nor2_1
X_17271_ net2159 net189 net1797 net9220 VGND VGND VPWR VPWR _00365_ sky130_fd_sc_hd__a22o_1
X_14483_ net7340 net5294 VGND VGND VPWR VPWR _06668_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19010_ _10845_ _10846_ VGND VGND VPWR VPWR _10847_ sky130_fd_sc_hd__nor2_1
X_16222_ _08283_ _08285_ VGND VGND VPWR VPWR _08287_ sky130_fd_sc_hd__nand2_1
X_13434_ net7866 net1577 VGND VGND VPWR VPWR _05707_ sky130_fd_sc_hd__nand2_1
XFILLER_0_180_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16153_ net2223 _08114_ _08116_ _08217_ _08218_ VGND VGND VPWR VPWR _08219_ sky130_fd_sc_hd__a311o_1
X_13365_ _05637_ _05541_ _05542_ VGND VGND VPWR VPWR _05638_ sky130_fd_sc_hd__nand3_1
Xclkbuf_leaf_102_clk clknet_4_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_102_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_140_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15104_ net4126 net4124 net4153 net4148 VGND VGND VPWR VPWR _07178_ sky130_fd_sc_hd__o22a_1
XFILLER_0_23_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16084_ _08066_ _08073_ VGND VGND VPWR VPWR _08151_ sky130_fd_sc_hd__nand2_1
X_13296_ _05558_ _05561_ VGND VGND VPWR VPWR _05569_ sky130_fd_sc_hd__or2b_1
Xwire5260 net5261 VGND VGND VPWR VPWR net5260 sky130_fd_sc_hd__clkbuf_1
Xwire5271 net5272 VGND VGND VPWR VPWR net5271 sky130_fd_sc_hd__clkbuf_1
X_19912_ net2097 _11696_ _11743_ VGND VGND VPWR VPWR _11744_ sky130_fd_sc_hd__o21ai_1
X_15035_ net3496 net2808 VGND VGND VPWR VPWR _07109_ sky130_fd_sc_hd__nor2_1
Xwire5282 matmul0.beta_pass\[4\] VGND VGND VPWR VPWR net5282 sky130_fd_sc_hd__buf_1
Xwire5293 net5294 VGND VGND VPWR VPWR net5293 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4581 net4582 VGND VGND VPWR VPWR net4581 sky130_fd_sc_hd__buf_1
X_19843_ _11651_ net1747 VGND VGND VPWR VPWR _11676_ sky130_fd_sc_hd__and2b_1
Xwire4592 net4593 VGND VGND VPWR VPWR net4592 sky130_fd_sc_hd__buf_1
Xwire3880 net3881 VGND VGND VPWR VPWR net3880 sky130_fd_sc_hd__buf_1
Xwire3891 net3892 VGND VGND VPWR VPWR net3891 sky130_fd_sc_hd__clkbuf_1
X_19774_ _11606_ _11608_ VGND VGND VPWR VPWR _11609_ sky130_fd_sc_hd__xnor2_2
X_16986_ _08821_ _08930_ net4062 VGND VGND VPWR VPWR _08948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18725_ net1066 VGND VGND VPWR VPWR _10570_ sky130_fd_sc_hd__inv_2
X_15937_ _07909_ _08004_ _08005_ VGND VGND VPWR VPWR _08006_ sky130_fd_sc_hd__o21a_1
XFILLER_0_64_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15868_ net2723 net2627 VGND VGND VPWR VPWR _07937_ sky130_fd_sc_hd__nor2_1
X_18656_ net605 _10456_ VGND VGND VPWR VPWR _10503_ sky130_fd_sc_hd__nand2_1
X_17607_ _09393_ svm0.tB\[11\] _09485_ _09487_ VGND VGND VPWR VPWR _09488_ sky130_fd_sc_hd__a211o_1
X_14819_ net7438 net7166 _04884_ VGND VGND VPWR VPWR _06926_ sky130_fd_sc_hd__and3_1
X_15799_ _07863_ _07868_ VGND VGND VPWR VPWR _07869_ sky130_fd_sc_hd__xnor2_2
X_18587_ net3953 _10434_ net3924 net3299 _10220_ VGND VGND VPWR VPWR _10435_ sky130_fd_sc_hd__a221o_1
XFILLER_0_80_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17538_ net6685 svm0.tC\[15\] VGND VGND VPWR VPWR _09420_ sky130_fd_sc_hd__xor2_1
XFILLER_0_188_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17469_ net4014 _09360_ VGND VGND VPWR VPWR _09362_ sky130_fd_sc_hd__nor2_1
XFILLER_0_190_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19208_ _11030_ _11033_ _11040_ _11044_ VGND VGND VPWR VPWR _11045_ sky130_fd_sc_hd__a22o_1
X_20480_ net6804 net6763 net6523 VGND VGND VPWR VPWR _12269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19139_ _10939_ _10975_ VGND VGND VPWR VPWR _10976_ sky130_fd_sc_hd__or2b_1
XFILLER_0_42_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22150_ _02152_ _02155_ VGND VGND VPWR VPWR _02156_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21101_ net5564 net5949 VGND VGND VPWR VPWR _01117_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22081_ _02085_ _02086_ _02087_ VGND VGND VPWR VPWR _02088_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21032_ _00986_ _01047_ VGND VGND VPWR VPWR _01048_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_160_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25840_ clknet_leaf_38_clk _00713_ net8743 VGND VGND VPWR VPWR pid_q.mult0.b\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1207 _10291_ VGND VGND VPWR VPWR net1207 sky130_fd_sc_hd__buf_1
Xwire1218 net1219 VGND VGND VPWR VPWR net1218 sky130_fd_sc_hd__buf_1
Xwire1229 net1230 VGND VGND VPWR VPWR net1229 sky130_fd_sc_hd__buf_1
X_25771_ clknet_leaf_27_clk _00644_ net8650 VGND VGND VPWR VPWR pid_d.out\[12\] sky130_fd_sc_hd__dfrtp_1
X_22983_ _02859_ VGND VGND VPWR VPWR _00658_ sky130_fd_sc_hd__clkbuf_1
X_24722_ net8017 _04552_ _04555_ VGND VGND VPWR VPWR _04556_ sky130_fd_sc_hd__a21o_1
XFILLER_0_179_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21934_ net5799 net5393 VGND VGND VPWR VPWR _01942_ sky130_fd_sc_hd__nand2_2
X_24653_ net7477 net8862 net2146 VGND VGND VPWR VPWR _04507_ sky130_fd_sc_hd__a21o_1
XFILLER_0_195_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21865_ net3780 net3788 _01865_ _01872_ net3776 VGND VGND VPWR VPWR _01874_ sky130_fd_sc_hd__o32a_1
Xfanout8708 net8713 VGND VGND VPWR VPWR net8708 sky130_fd_sc_hd__buf_1
X_23604_ _03307_ net646 net640 _03469_ _03471_ VGND VGND VPWR VPWR _03472_ sky130_fd_sc_hd__a32o_1
XFILLER_0_166_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length5202 net5203 VGND VGND VPWR VPWR net5202 sky130_fd_sc_hd__clkbuf_1
X_20816_ _00823_ _00831_ VGND VGND VPWR VPWR _00832_ sky130_fd_sc_hd__xnor2_1
X_24584_ _04412_ _04439_ VGND VGND VPWR VPWR _04440_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21796_ _01718_ _01720_ _01805_ VGND VGND VPWR VPWR _01806_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4501 net4502 VGND VGND VPWR VPWR net4501 sky130_fd_sc_hd__buf_1
Xwire8825 net8826 VGND VGND VPWR VPWR net8825 sky130_fd_sc_hd__clkbuf_1
X_23535_ _03401_ _03402_ VGND VGND VPWR VPWR _03403_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8836 net8837 VGND VGND VPWR VPWR net8836 sky130_fd_sc_hd__clkbuf_1
X_20747_ _12514_ _12517_ VGND VGND VPWR VPWR _12518_ sky130_fd_sc_hd__xnor2_2
Xwire8847 net8848 VGND VGND VPWR VPWR net8847 sky130_fd_sc_hd__clkbuf_1
Xwire8858 net8859 VGND VGND VPWR VPWR net8858 sky130_fd_sc_hd__clkbuf_1
Xwire504 net505 VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire515 net516 VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23466_ _03326_ _03334_ VGND VGND VPWR VPWR _03335_ sky130_fd_sc_hd__xnor2_2
Xwire526 _10612_ VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__buf_1
Xwire537 _04115_ VGND VGND VPWR VPWR net537 sky130_fd_sc_hd__clkbuf_1
X_20678_ _12451_ _12453_ VGND VGND VPWR VPWR _12454_ sky130_fd_sc_hd__xor2_1
XFILLER_0_169_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length3844 _12499_ VGND VGND VPWR VPWR net3844 sky130_fd_sc_hd__buf_1
Xwire548 _03310_ VGND VGND VPWR VPWR net548 sky130_fd_sc_hd__clkbuf_1
X_25205_ clknet_leaf_57_clk _00094_ net8715 VGND VGND VPWR VPWR matmul0.b_in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_22417_ _02352_ _02353_ _02418_ VGND VGND VPWR VPWR _02419_ sky130_fd_sc_hd__o21ai_2
Xwire559 _01426_ VGND VGND VPWR VPWR net559 sky130_fd_sc_hd__clkbuf_1
X_23397_ net5150 net4525 VGND VGND VPWR VPWR _03267_ sky130_fd_sc_hd__nand2_1
Xmax_length3899 net3900 VGND VGND VPWR VPWR net3899 sky130_fd_sc_hd__clkbuf_1
X_25136_ clknet_leaf_51_clk _00025_ net8809 VGND VGND VPWR VPWR svm0.tC\[8\] sky130_fd_sc_hd__dfrtp_1
X_13150_ _05421_ _05422_ VGND VGND VPWR VPWR _05423_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22348_ _02348_ _02350_ VGND VGND VPWR VPWR _02351_ sky130_fd_sc_hd__xor2_2
XFILLER_0_131_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13081_ net4259 _05351_ VGND VGND VPWR VPWR _05354_ sky130_fd_sc_hd__nor2_1
X_25067_ net4424 net1994 _04812_ VGND VGND VPWR VPWR _04815_ sky130_fd_sc_hd__nor3_1
X_22279_ net2052 _02219_ _02282_ VGND VGND VPWR VPWR _02283_ sky130_fd_sc_hd__o21a_1
Xwire3110 _01609_ VGND VGND VPWR VPWR net3110 sky130_fd_sc_hd__clkbuf_1
X_24018_ net4534 net4952 VGND VGND VPWR VPWR _03881_ sky130_fd_sc_hd__nand2_1
Xwire3132 net3134 VGND VGND VPWR VPWR net3132 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold190 svm0.tA\[12\] VGND VGND VPWR VPWR net9143 sky130_fd_sc_hd__dlygate4sd3_1
Xwire3154 _11376_ VGND VGND VPWR VPWR net3154 sky130_fd_sc_hd__buf_1
Xwire2420 net2421 VGND VGND VPWR VPWR net2420 sky130_fd_sc_hd__clkbuf_2
Xwire3165 net3168 VGND VGND VPWR VPWR net3165 sky130_fd_sc_hd__buf_1
Xwire2431 _02995_ VGND VGND VPWR VPWR net2431 sky130_fd_sc_hd__buf_1
Xwire3176 net3177 VGND VGND VPWR VPWR net3176 sky130_fd_sc_hd__buf_1
Xwire2442 net2443 VGND VGND VPWR VPWR net2442 sky130_fd_sc_hd__clkbuf_1
Xwire3187 net3188 VGND VGND VPWR VPWR net3187 sky130_fd_sc_hd__clkbuf_2
X_16840_ net6423 matmul0.sin\[8\] net3366 VGND VGND VPWR VPWR _08811_ sky130_fd_sc_hd__mux2_1
Xwire2453 net2454 VGND VGND VPWR VPWR net2453 sky130_fd_sc_hd__clkbuf_1
Xwire2475 _01785_ VGND VGND VPWR VPWR net2475 sky130_fd_sc_hd__buf_1
Xwire1730 _01272_ VGND VGND VPWR VPWR net1730 sky130_fd_sc_hd__buf_1
XFILLER_0_137_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1741 _12365_ VGND VGND VPWR VPWR net1741 sky130_fd_sc_hd__clkbuf_1
X_16771_ matmul0.a_in\[5\] matmul0.a\[5\] net3378 VGND VGND VPWR VPWR _08775_ sky130_fd_sc_hd__mux2_1
Xwire2486 _12525_ VGND VGND VPWR VPWR net2486 sky130_fd_sc_hd__buf_1
XFILLER_0_189_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13983_ _06246_ _06247_ VGND VGND VPWR VPWR _06248_ sky130_fd_sc_hd__and2_1
Xwire1752 _11172_ VGND VGND VPWR VPWR net1752 sky130_fd_sc_hd__clkbuf_1
Xwire2497 _11858_ VGND VGND VPWR VPWR net2497 sky130_fd_sc_hd__clkbuf_1
Xwire1763 net1764 VGND VGND VPWR VPWR net1763 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15722_ net1852 _07658_ _07651_ VGND VGND VPWR VPWR _07793_ sky130_fd_sc_hd__o21a_1
X_18510_ _09660_ _10304_ net3229 VGND VGND VPWR VPWR _10359_ sky130_fd_sc_hd__mux2_1
Xwire1774 _10230_ VGND VGND VPWR VPWR net1774 sky130_fd_sc_hd__buf_1
XFILLER_0_73_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12934_ _05126_ net791 VGND VGND VPWR VPWR _05207_ sky130_fd_sc_hd__and2_1
Xwire1785 net1786 VGND VGND VPWR VPWR net1785 sky130_fd_sc_hd__buf_1
Xwire1796 _09203_ VGND VGND VPWR VPWR net1796 sky130_fd_sc_hd__buf_1
X_19490_ _11326_ VGND VGND VPWR VPWR _11327_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15653_ net2250 net2672 _07717_ _07724_ VGND VGND VPWR VPWR _07725_ sky130_fd_sc_hd__o211a_1
X_18441_ _10281_ _10290_ VGND VGND VPWR VPWR _10291_ sky130_fd_sc_hd__xnor2_1
X_12865_ net7931 _05057_ _05136_ VGND VGND VPWR VPWR _05138_ sky130_fd_sc_hd__a21oi_1
X_14604_ net3641 _06776_ VGND VGND VPWR VPWR _06777_ sky130_fd_sc_hd__nor2_1
X_18372_ net6825 _10222_ VGND VGND VPWR VPWR _10223_ sky130_fd_sc_hd__xnor2_2
X_15584_ net2805 net3466 VGND VGND VPWR VPWR _07656_ sky130_fd_sc_hd__nor2_1
X_12796_ _04935_ _04939_ _04916_ VGND VGND VPWR VPWR _05069_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17323_ net4032 net7943 VGND VGND VPWR VPWR _09237_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14535_ _06710_ _06711_ _06713_ VGND VGND VPWR VPWR _06714_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_172_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17254_ net2958 net174 net2163 net9165 VGND VGND VPWR VPWR _00352_ sky130_fd_sc_hd__a22o_1
X_14466_ net1990 net2887 VGND VGND VPWR VPWR _06654_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16205_ net2752 net3416 VGND VGND VPWR VPWR _08270_ sky130_fd_sc_hd__nor2_1
X_13417_ _05688_ net2944 VGND VGND VPWR VPWR _05690_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17185_ net618 _09129_ net6850 VGND VGND VPWR VPWR _09136_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14397_ net5297 net1298 net2895 net4463 _06600_ VGND VGND VPWR VPWR _06601_ sky130_fd_sc_hd__a221o_1
XFILLER_0_141_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16136_ net1516 _08103_ _08201_ VGND VGND VPWR VPWR _08202_ sky130_fd_sc_hd__o21a_1
X_13348_ net7893 _05527_ _05618_ _05620_ VGND VGND VPWR VPWR _05621_ sky130_fd_sc_hd__a211o_1
X_16067_ net2205 net1258 VGND VGND VPWR VPWR _08134_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13279_ _05550_ _05551_ VGND VGND VPWR VPWR _05552_ sky130_fd_sc_hd__nor2_1
Xwire5090 net5083 VGND VGND VPWR VPWR net5090 sky130_fd_sc_hd__buf_1
X_15018_ _07078_ VGND VGND VPWR VPWR _07092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19826_ _11656_ _11659_ VGND VGND VPWR VPWR _11660_ sky130_fd_sc_hd__xnor2_2
X_19757_ _11586_ net2099 VGND VGND VPWR VPWR _11592_ sky130_fd_sc_hd__xnor2_2
X_16969_ net6325 net6309 net6277 net6254 net6518 net6498 VGND VGND VPWR VPWR _08932_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18708_ net6772 _10553_ VGND VGND VPWR VPWR _10554_ sky130_fd_sc_hd__nand2_1
XFILLER_0_190_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19688_ net3157 _11523_ VGND VGND VPWR VPWR _11524_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_195_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18639_ net6830 net3282 VGND VGND VPWR VPWR _10486_ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21650_ net5609 net5653 VGND VGND VPWR VPWR _01661_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_59_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20601_ net8057 net6212 net1554 _12382_ VGND VGND VPWR VPWR _00508_ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21581_ net5384 _01592_ VGND VGND VPWR VPWR _01593_ sky130_fd_sc_hd__nand2_2
XFILLER_0_191_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23320_ _03186_ _03189_ VGND VGND VPWR VPWR _03190_ sky130_fd_sc_hd__xnor2_1
X_20532_ net6756 _08944_ net2490 _08924_ VGND VGND VPWR VPWR _12318_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire6708 net6705 VGND VGND VPWR VPWR net6708 sky130_fd_sc_hd__buf_1
Xwire6719 net6724 VGND VGND VPWR VPWR net6719 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23251_ _03014_ _03024_ _03019_ VGND VGND VPWR VPWR _03121_ sky130_fd_sc_hd__o21ai_1
X_20463_ net3667 _12224_ _12254_ VGND VGND VPWR VPWR _12255_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_7_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22202_ net944 net1706 VGND VGND VPWR VPWR _02207_ sky130_fd_sc_hd__xor2_2
X_23182_ _03049_ _03050_ VGND VGND VPWR VPWR _03052_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20394_ _08836_ net1501 VGND VGND VPWR VPWR _12192_ sky130_fd_sc_hd__nand2_1
X_22133_ _02137_ _02138_ VGND VGND VPWR VPWR _02139_ sky130_fd_sc_hd__or2b_1
XFILLER_0_3_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22064_ net1715 _01969_ VGND VGND VPWR VPWR _02071_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21015_ _00995_ _01030_ VGND VGND VPWR VPWR _01031_ sky130_fd_sc_hd__nand2_1
Xwire1004 _05198_ VGND VGND VPWR VPWR net1004 sky130_fd_sc_hd__clkbuf_2
Xwire1015 _04006_ VGND VGND VPWR VPWR net1015 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1026 net1027 VGND VGND VPWR VPWR net1026 sky130_fd_sc_hd__clkbuf_1
X_25823_ clknet_leaf_31_clk _00696_ net8684 VGND VGND VPWR VPWR pid_q.prev_error\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1037 _02149_ VGND VGND VPWR VPWR net1037 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1048 _01746_ VGND VGND VPWR VPWR net1048 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1059 _11526_ VGND VGND VPWR VPWR net1059 sky130_fd_sc_hd__clkbuf_1
X_25754_ clknet_leaf_13_clk _00627_ net8614 VGND VGND VPWR VPWR pid_d.kp\[12\] sky130_fd_sc_hd__dfrtp_1
X_22966_ matmul0.beta_pass\[2\] net2613 net6569 VGND VGND VPWR VPWR _02851_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24705_ _04541_ VGND VGND VPWR VPWR _04542_ sky130_fd_sc_hd__buf_1
X_21917_ _01825_ _01826_ _01923_ _01924_ VGND VGND VPWR VPWR _01925_ sky130_fd_sc_hd__a31o_1
X_25685_ clknet_leaf_5_clk _00558_ net8566 VGND VGND VPWR VPWR pid_d.curr_error\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_22897_ net342 net2033 _02790_ VGND VGND VPWR VPWR _02791_ sky130_fd_sc_hd__a21o_1
X_24636_ _04487_ _04490_ VGND VGND VPWR VPWR _04491_ sky130_fd_sc_hd__xnor2_1
X_12650_ net7362 net3030 net3695 VGND VGND VPWR VPWR _04923_ sky130_fd_sc_hd__nand3_1
Xfanout8505 net8517 VGND VGND VPWR VPWR net8505 sky130_fd_sc_hd__buf_1
X_21848_ _01845_ _01856_ VGND VGND VPWR VPWR _01857_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8600 net8601 VGND VGND VPWR VPWR net8600 sky130_fd_sc_hd__clkbuf_1
Xwire8611 net8612 VGND VGND VPWR VPWR net8611 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24567_ _04414_ _04422_ VGND VGND VPWR VPWR _04423_ sky130_fd_sc_hd__xnor2_2
X_12581_ net4309 VGND VGND VPWR VPWR _04867_ sky130_fd_sc_hd__buf_1
X_21779_ _01680_ _01683_ _01677_ VGND VGND VPWR VPWR _01789_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14320_ net6447 _06530_ _06531_ _06541_ VGND VGND VPWR VPWR _06542_ sky130_fd_sc_hd__a211o_1
X_23518_ pid_q.prev_error\[0\] pid_q.curr_error\[0\] _03385_ VGND VGND VPWR VPWR _03387_
+ sky130_fd_sc_hd__a21oi_1
Xwire7910 net7905 VGND VGND VPWR VPWR net7910 sky130_fd_sc_hd__clkbuf_1
Xwire301 _02253_ VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__clkbuf_1
Xwire8655 net8656 VGND VGND VPWR VPWR net8655 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire7921 net7922 VGND VGND VPWR VPWR net7921 sky130_fd_sc_hd__buf_1
XFILLER_0_65_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24498_ _04284_ _04354_ VGND VGND VPWR VPWR _04355_ sky130_fd_sc_hd__xnor2_2
Xwire7932 net7933 VGND VGND VPWR VPWR net7932 sky130_fd_sc_hd__buf_1
Xmax_length4364 net4365 VGND VGND VPWR VPWR net4364 sky130_fd_sc_hd__buf_1
XFILLER_0_19_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire312 net313 VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length3630 _06800_ VGND VGND VPWR VPWR net3630 sky130_fd_sc_hd__buf_1
Xwire7943 net7944 VGND VGND VPWR VPWR net7943 sky130_fd_sc_hd__buf_1
XFILLER_0_163_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire334 net335 VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__clkbuf_1
Xwire8688 net8689 VGND VGND VPWR VPWR net8688 sky130_fd_sc_hd__buf_1
XFILLER_0_46_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7954 pid_q.target\[15\] VGND VGND VPWR VPWR net7954 sky130_fd_sc_hd__buf_1
Xwire345 _02099_ VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14251_ net6458 _06505_ VGND VGND VPWR VPWR _06506_ sky130_fd_sc_hd__nand2_1
Xwire7965 net7966 VGND VGND VPWR VPWR net7965 sky130_fd_sc_hd__clkbuf_1
X_23449_ net749 net796 VGND VGND VPWR VPWR _03318_ sky130_fd_sc_hd__or2_1
Xwire356 net357 VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__clkbuf_1
Xwire7976 net7977 VGND VGND VPWR VPWR net7976 sky130_fd_sc_hd__clkbuf_1
Xwire367 net368 VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__clkbuf_2
Xwire7987 net7988 VGND VGND VPWR VPWR net7987 sky130_fd_sc_hd__clkbuf_1
Xwire378 net379 VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__clkbuf_1
X_13202_ net734 _05473_ _05474_ VGND VGND VPWR VPWR _05475_ sky130_fd_sc_hd__a21oi_2
Xwire7998 net7999 VGND VGND VPWR VPWR net7998 sky130_fd_sc_hd__clkbuf_1
Xwire389 net390 VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__clkbuf_1
X_14182_ _06440_ _06441_ VGND VGND VPWR VPWR _06442_ sky130_fd_sc_hd__and2_1
Xmax_length2973 _04962_ VGND VGND VPWR VPWR net2973 sky130_fd_sc_hd__buf_1
X_13133_ _05349_ _05350_ VGND VGND VPWR VPWR _05406_ sky130_fd_sc_hd__nand2_1
X_25119_ net9215 net2393 net1993 net5978 VGND VGND VPWR VPWR _00800_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18990_ net6295 VGND VGND VPWR VPWR _10827_ sky130_fd_sc_hd__inv_2
X_13064_ _05279_ _05335_ _05336_ VGND VGND VPWR VPWR _05337_ sky130_fd_sc_hd__a21oi_1
X_17941_ net6916 _09791_ VGND VGND VPWR VPWR _09792_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17872_ _09605_ _09610_ VGND VGND VPWR VPWR _09723_ sky130_fd_sc_hd__nand2_1
Xwire2250 net2251 VGND VGND VPWR VPWR net2250 sky130_fd_sc_hd__buf_1
X_19611_ _10996_ net6013 VGND VGND VPWR VPWR _11448_ sky130_fd_sc_hd__nor2_1
Xwire2261 _06837_ VGND VGND VPWR VPWR net2261 sky130_fd_sc_hd__clkbuf_1
Xwire2272 net2273 VGND VGND VPWR VPWR net2272 sky130_fd_sc_hd__clkbuf_1
X_16823_ net6431 matmul0.sin\[0\] net3367 VGND VGND VPWR VPWR _08802_ sky130_fd_sc_hd__mux2_1
Xwire2294 net2295 VGND VGND VPWR VPWR net2294 sky130_fd_sc_hd__buf_1
XFILLER_0_75_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1560 _06292_ VGND VGND VPWR VPWR net1560 sky130_fd_sc_hd__clkbuf_2
Xwire1571 _05686_ VGND VGND VPWR VPWR net1571 sky130_fd_sc_hd__buf_1
X_19542_ net6073 net6029 VGND VGND VPWR VPWR _11379_ sky130_fd_sc_hd__xnor2_2
X_13966_ _06229_ _06230_ VGND VGND VPWR VPWR _06231_ sky130_fd_sc_hd__xor2_1
Xwire1582 _05555_ VGND VGND VPWR VPWR net1582 sky130_fd_sc_hd__buf_1
X_16754_ net7559 matmul0.b\[13\] net3381 VGND VGND VPWR VPWR _08766_ sky130_fd_sc_hd__mux2_1
Xmax_cap3 _02716_ VGND VGND VPWR VPWR net9248 sky130_fd_sc_hd__buf_1
Xwire1593 _05215_ VGND VGND VPWR VPWR net1593 sky130_fd_sc_hd__dlymetal6s2s_1
X_12917_ net5232 _04856_ _04897_ _04889_ svm0.vC\[10\] VGND VGND VPWR VPWR _05190_
+ sky130_fd_sc_hd__a32oi_1
X_15705_ _07680_ net1266 net1104 VGND VGND VPWR VPWR _07776_ sky130_fd_sc_hd__a21bo_1
X_19473_ _11280_ _11281_ VGND VGND VPWR VPWR _11310_ sky130_fd_sc_hd__nor2_1
X_16685_ matmul0.matmul_stage_inst.mult1\[9\] VGND VGND VPWR VPWR _08716_ sky130_fd_sc_hd__inv_2
X_13897_ _06132_ _06133_ VGND VGND VPWR VPWR _06163_ sky130_fd_sc_hd__or2b_1
XFILLER_0_159_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18424_ _10211_ _10270_ _10273_ VGND VGND VPWR VPWR _10274_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_185_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12848_ _05119_ _05120_ VGND VGND VPWR VPWR _05121_ sky130_fd_sc_hd__nand2_1
X_15636_ _07680_ _07707_ VGND VGND VPWR VPWR _07708_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15567_ net574 _07639_ VGND VGND VPWR VPWR _07640_ sky130_fd_sc_hd__xnor2_1
X_18355_ net6773 _10155_ VGND VGND VPWR VPWR _10206_ sky130_fd_sc_hd__nand2_1
X_12779_ net6665 net6599 net6748 VGND VGND VPWR VPWR _05052_ sky130_fd_sc_hd__and3b_1
X_17306_ _09214_ _09217_ _09219_ net6691 VGND VGND VPWR VPWR _09220_ sky130_fd_sc_hd__a31oi_1
X_14518_ _06692_ _06698_ VGND VGND VPWR VPWR _06699_ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15498_ net4119 net4114 net4087 net4086 VGND VGND VPWR VPWR _07571_ sky130_fd_sc_hd__o22a_1
X_18286_ _10131_ _10136_ VGND VGND VPWR VPWR _10137_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_160_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14449_ net5197 net1548 net3647 net4397 _06640_ VGND VGND VPWR VPWR _06641_ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17237_ net6759 _09183_ _09184_ VGND VGND VPWR VPWR _00341_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_25_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17168_ net1921 _09119_ net8048 net6891 VGND VGND VPWR VPWR _09121_ sky130_fd_sc_hd__o211a_1
Xwire890 net891 VGND VGND VPWR VPWR net890 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16119_ net1254 net1253 VGND VGND VPWR VPWR _08185_ sky130_fd_sc_hd__nor2_2
X_17099_ net5992 net4038 net4057 _09055_ VGND VGND VPWR VPWR _09056_ sky130_fd_sc_hd__o22a_1
XFILLER_0_161_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19809_ _11641_ _11642_ VGND VGND VPWR VPWR _11643_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_193_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22820_ net3759 VGND VGND VPWR VPWR _02722_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22751_ pid_d.ki\[8\] net3072 net1696 VGND VGND VPWR VPWR _02679_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_91_clk clknet_4_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_91_clk sky130_fd_sc_hd__clkbuf_16
X_21702_ net1721 _01599_ _01712_ VGND VGND VPWR VPWR _01713_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25470_ clknet_leaf_51_clk _00350_ net8811 VGND VGND VPWR VPWR svm0.tB\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22682_ _02629_ net5580 net2448 VGND VGND VPWR VPWR _02630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24421_ _04272_ _04278_ VGND VGND VPWR VPWR _04279_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_191_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21633_ pid_d.prev_int\[4\] VGND VGND VPWR VPWR _01644_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7206 net7207 VGND VGND VPWR VPWR net7206 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24352_ _04209_ _04210_ VGND VGND VPWR VPWR _04211_ sky130_fd_sc_hd__xor2_2
Xwire7217 matmul0.alpha_pass\[13\] VGND VGND VPWR VPWR net7217 sky130_fd_sc_hd__clkbuf_1
X_21564_ _01466_ _01468_ _01467_ VGND VGND VPWR VPWR _01576_ sky130_fd_sc_hd__o21a_1
Xwire7228 net7229 VGND VGND VPWR VPWR net7228 sky130_fd_sc_hd__clkbuf_1
Xwire7239 net7240 VGND VGND VPWR VPWR net7239 sky130_fd_sc_hd__clkbuf_1
X_23303_ _03152_ _03149_ _03167_ VGND VGND VPWR VPWR _03173_ sky130_fd_sc_hd__and3b_1
XFILLER_0_173_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6505 cordic0.gm0.iter\[1\] VGND VGND VPWR VPWR net6505 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20515_ net1484 net2082 net2084 VGND VGND VPWR VPWR _12302_ sky130_fd_sc_hd__nand3_1
Xwire6516 net6515 VGND VGND VPWR VPWR net6516 sky130_fd_sc_hd__dlymetal6s2s_1
X_24283_ _04137_ _04142_ VGND VGND VPWR VPWR _04143_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_160_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21495_ net5651 _01402_ VGND VGND VPWR VPWR _01508_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6538 net6535 VGND VGND VPWR VPWR net6538 sky130_fd_sc_hd__buf_1
XFILLER_0_90_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5804 net5805 VGND VGND VPWR VPWR net5804 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire6549 net6551 VGND VGND VPWR VPWR net6549 sky130_fd_sc_hd__buf_1
X_23234_ _03097_ _03100_ _03103_ VGND VGND VPWR VPWR _03104_ sky130_fd_sc_hd__a21o_1
Xwire5815 net5809 VGND VGND VPWR VPWR net5815 sky130_fd_sc_hd__buf_1
Xwire5826 net5819 VGND VGND VPWR VPWR net5826 sky130_fd_sc_hd__clkbuf_1
X_20446_ net3354 net6369 net1229 _12239_ VGND VGND VPWR VPWR _00496_ sky130_fd_sc_hd__a22o_1
Xwire5837 net5838 VGND VGND VPWR VPWR net5837 sky130_fd_sc_hd__buf_1
Xwire5848 net5849 VGND VGND VPWR VPWR net5848 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5859 net5856 VGND VGND VPWR VPWR net5859 sky130_fd_sc_hd__buf_1
X_23165_ _03015_ _03034_ VGND VGND VPWR VPWR _03035_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_113_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20377_ _06504_ _12175_ _12098_ VGND VGND VPWR VPWR _12176_ sky130_fd_sc_hd__o21a_1
XFILLER_0_101_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22116_ _00917_ net5661 VGND VGND VPWR VPWR _02122_ sky130_fd_sc_hd__nand2_1
X_23096_ net4904 net4771 VGND VGND VPWR VPWR _02966_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22047_ net3780 net5395 _01964_ VGND VGND VPWR VPWR _02054_ sky130_fd_sc_hd__or3_1
XFILLER_0_100_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13820_ _06064_ _06073_ _06024_ VGND VGND VPWR VPWR _06087_ sky130_fd_sc_hd__a21bo_1
X_25806_ clknet_leaf_30_clk _00679_ net8675 VGND VGND VPWR VPWR pid_q.curr_int\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_23998_ pid_q.curr_int\[6\] VGND VGND VPWR VPWR _03861_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13751_ _05866_ _05872_ net404 _06017_ _06018_ VGND VGND VPWR VPWR _06019_ sky130_fd_sc_hd__o311a_1
X_25737_ clknet_leaf_12_clk _00610_ net8822 VGND VGND VPWR VPWR pid_d.ki\[11\] sky130_fd_sc_hd__dfrtp_1
X_22949_ _02386_ _02836_ _02515_ VGND VGND VPWR VPWR _02837_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_82_clk clknet_4_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_82_clk sky130_fd_sc_hd__clkbuf_16
X_12702_ net2972 VGND VGND VPWR VPWR _04975_ sky130_fd_sc_hd__clkbuf_1
X_16470_ _08471_ _08530_ VGND VGND VPWR VPWR _08531_ sky130_fd_sc_hd__xor2_1
X_13682_ _05948_ _05949_ net1923 VGND VGND VPWR VPWR _05951_ sky130_fd_sc_hd__o21ai_1
X_25668_ clknet_leaf_120_clk _00541_ net8394 VGND VGND VPWR VPWR pid_d.prev_error\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15421_ _07493_ _07494_ VGND VGND VPWR VPWR _07495_ sky130_fd_sc_hd__nor2_1
X_24619_ _04435_ _04468_ _04471_ _04473_ VGND VGND VPWR VPWR _04474_ sky130_fd_sc_hd__o211a_1
X_12633_ net5276 _04856_ _04897_ _04889_ svm0.vC\[4\] VGND VGND VPWR VPWR _04906_
+ sky130_fd_sc_hd__a32oi_1
Xfanout7601 net7611 VGND VGND VPWR VPWR net7601 sky130_fd_sc_hd__clkbuf_1
Xfanout8357 net8361 VGND VGND VPWR VPWR net8357 sky130_fd_sc_hd__buf_1
X_25599_ clknet_leaf_105_clk _00472_ net8354 VGND VGND VPWR VPWR cordic0.slte0.opB\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8430 net8429 VGND VGND VPWR VPWR net8430 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_136_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout7634 svm0.periodTop\[14\] VGND VGND VPWR VPWR net7634 sky130_fd_sc_hd__clkbuf_1
X_18140_ _09944_ _09990_ _09901_ VGND VGND VPWR VPWR _09991_ sky130_fd_sc_hd__mux2_1
X_15352_ _07424_ _07425_ VGND VGND VPWR VPWR _07426_ sky130_fd_sc_hd__xnor2_1
X_12564_ matmul0.start VGND VGND VPWR VPWR _04854_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8463 net8462 VGND VGND VPWR VPWR net8463 sky130_fd_sc_hd__buf_1
X_14303_ _06524_ VGND VGND VPWR VPWR _06525_ sky130_fd_sc_hd__buf_1
Xwire7740 net7734 VGND VGND VPWR VPWR net7740 sky130_fd_sc_hd__buf_1
XFILLER_0_123_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18071_ _09918_ _09920_ VGND VGND VPWR VPWR _09922_ sky130_fd_sc_hd__nand2_1
Xwire8485 net8486 VGND VGND VPWR VPWR net8485 sky130_fd_sc_hd__clkbuf_1
Xwire7751 net7752 VGND VGND VPWR VPWR net7751 sky130_fd_sc_hd__clkbuf_1
X_15283_ net2839 _07045_ _07050_ _07051_ VGND VGND VPWR VPWR _07357_ sky130_fd_sc_hd__or4_1
Xwire153 _06495_ VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__buf_1
XFILLER_0_53_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7773 net7774 VGND VGND VPWR VPWR net7773 sky130_fd_sc_hd__clkbuf_1
X_17022_ net7053 net1553 VGND VGND VPWR VPWR _08983_ sky130_fd_sc_hd__nor2_1
Xwire164 net165 VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_1
X_14234_ net7629 net1304 net1119 VGND VGND VPWR VPWR _06491_ sky130_fd_sc_hd__a21o_1
Xwire175 net176 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__buf_1
XFILLER_0_123_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7784 net7777 VGND VGND VPWR VPWR net7784 sky130_fd_sc_hd__buf_1
XFILLER_0_34_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7795 net7796 VGND VGND VPWR VPWR net7795 sky130_fd_sc_hd__clkbuf_1
Xmax_length3482 net3483 VGND VGND VPWR VPWR net3482 sky130_fd_sc_hd__buf_1
Xwire186 _08545_ VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_1
Xwire197 _04501_ VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14165_ _06366_ _06425_ _06395_ _06368_ VGND VGND VPWR VPWR _06426_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_22_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13116_ _05266_ _05267_ net7847 net1601 VGND VGND VPWR VPWR _05389_ sky130_fd_sc_hd__o211ai_2
X_14096_ net366 VGND VGND VPWR VPWR _06359_ sky130_fd_sc_hd__inv_2
X_18973_ net6339 net6318 VGND VGND VPWR VPWR _10810_ sky130_fd_sc_hd__or2b_1
X_13047_ _05211_ net535 _05317_ _05319_ VGND VGND VPWR VPWR _05320_ sky130_fd_sc_hd__or4bb_1
X_17924_ _09761_ _09771_ _09773_ VGND VGND VPWR VPWR _09775_ sky130_fd_sc_hd__or3_1
X_17855_ net7097 _09701_ _09702_ net7033 _09705_ VGND VGND VPWR VPWR _09706_ sky130_fd_sc_hd__a221o_1
XFILLER_0_56_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire2080 net2081 VGND VGND VPWR VPWR net2080 sky130_fd_sc_hd__clkbuf_1
Xwire2091 _12086_ VGND VGND VPWR VPWR net2091 sky130_fd_sc_hd__buf_1
XFILLER_0_191_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16806_ _08793_ VGND VGND VPWR VPWR _00301_ sky130_fd_sc_hd__clkbuf_1
X_17786_ net7022 net7036 VGND VGND VPWR VPWR _09637_ sky130_fd_sc_hd__nor2_1
X_14998_ _07008_ _07071_ VGND VGND VPWR VPWR _07072_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1390 _01300_ VGND VGND VPWR VPWR net1390 sky130_fd_sc_hd__buf_1
X_19525_ _11358_ _11361_ VGND VGND VPWR VPWR _11362_ sky130_fd_sc_hd__xor2_1
X_16737_ net7571 matmul0.b\[5\] net3702 VGND VGND VPWR VPWR _08757_ sky130_fd_sc_hd__mux2_1
X_13949_ _06213_ _06214_ VGND VGND VPWR VPWR _06215_ sky130_fd_sc_hd__and2b_1
XFILLER_0_72_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_73_clk clknet_4_10__leaf_clk VGND VGND VPWR VPWR clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_159_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19456_ net3869 _11292_ VGND VGND VPWR VPWR _11293_ sky130_fd_sc_hd__nor2_1
X_16668_ _08700_ _08701_ VGND VGND VPWR VPWR _08702_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18407_ net767 _10205_ VGND VGND VPWR VPWR _10258_ sky130_fd_sc_hd__or2b_1
X_15619_ net2675 _07690_ VGND VGND VPWR VPWR _07691_ sky130_fd_sc_hd__xnor2_1
X_19387_ net6358 _11221_ _11223_ _11220_ VGND VGND VPWR VPWR _11224_ sky130_fd_sc_hd__o211ai_1
X_16599_ _08649_ VGND VGND VPWR VPWR _00238_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18338_ net3228 _10187_ _10188_ VGND VGND VPWR VPWR _10189_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_114_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18269_ _10117_ _10118_ _10119_ VGND VGND VPWR VPWR _10120_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_62_Left_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_188_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20300_ net9160 _12104_ _12105_ VGND VGND VPWR VPWR _00484_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_86_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21280_ net5702 net5615 VGND VGND VPWR VPWR _01295_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20231_ _12049_ VGND VGND VPWR VPWR _00471_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3709 _04873_ VGND VGND VPWR VPWR net3709 sky130_fd_sc_hd__buf_1
X_20162_ net3126 _11967_ net244 VGND VGND VPWR VPWR _11989_ sky130_fd_sc_hd__o21bai_1
X_24970_ pid_q.kp\[4\] _04710_ net1359 VGND VGND VPWR VPWR _04740_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20093_ _11914_ _11846_ _11915_ _11918_ _11921_ VGND VGND VPWR VPWR _11922_ sky130_fd_sc_hd__o32a_1
XFILLER_0_196_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23921_ _03783_ _03784_ VGND VGND VPWR VPWR _03785_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_71_Left_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23852_ net4596 net4921 VGND VGND VPWR VPWR _03717_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length8427 net8428 VGND VGND VPWR VPWR net8427 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_98_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22803_ _02709_ VGND VGND VPWR VPWR _00628_ sky130_fd_sc_hd__clkbuf_1
X_23783_ _03647_ _03648_ VGND VGND VPWR VPWR _03649_ sky130_fd_sc_hd__xnor2_1
X_20995_ net1732 _01009_ _01010_ VGND VGND VPWR VPWR _01011_ sky130_fd_sc_hd__nand3_1
Xclkbuf_leaf_64_clk clknet_4_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_16
X_25522_ clknet_leaf_47_clk _00402_ net8777 VGND VGND VPWR VPWR svm0.counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_22734_ _02667_ VGND VGND VPWR VPWR _00601_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25453_ clknet_leaf_112_clk _00336_ net8539 VGND VGND VPWR VPWR cordic0.vec\[1\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_22665_ net4301 _02463_ _02617_ VGND VGND VPWR VPWR _02618_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24404_ net5175 pid_q.prev_int\[12\] VGND VGND VPWR VPWR _04262_ sky130_fd_sc_hd__xor2_1
X_21616_ _01617_ _01627_ VGND VGND VPWR VPWR _01628_ sky130_fd_sc_hd__xor2_1
XFILLER_0_180_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7003 cordic0.vec\[1\]\[7\] VGND VGND VPWR VPWR net7003 sky130_fd_sc_hd__clkbuf_1
X_25384_ clknet_leaf_74_clk _00267_ net8473 VGND VGND VPWR VPWR matmul0.b\[3\] sky130_fd_sc_hd__dfrtp_1
Xwire7014 net7012 VGND VGND VPWR VPWR net7014 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_80_Left_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22596_ net8889 _02572_ VGND VGND VPWR VPWR _02573_ sky130_fd_sc_hd__and2_1
XFILLER_0_180_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7025 net7026 VGND VGND VPWR VPWR net7025 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24335_ _03942_ _04043_ _04106_ _04044_ VGND VGND VPWR VPWR _04194_ sky130_fd_sc_hd__a211oi_1
X_21547_ net5599 net5680 VGND VGND VPWR VPWR _01559_ sky130_fd_sc_hd__nand2_1
Xwire6302 net6304 VGND VGND VPWR VPWR net6302 sky130_fd_sc_hd__buf_1
XFILLER_0_8_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7047 net7048 VGND VGND VPWR VPWR net7047 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire7069 net7072 VGND VGND VPWR VPWR net7069 sky130_fd_sc_hd__buf_1
Xwire6335 net6336 VGND VGND VPWR VPWR net6335 sky130_fd_sc_hd__buf_1
XFILLER_0_90_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5601 net5602 VGND VGND VPWR VPWR net5601 sky130_fd_sc_hd__buf_1
Xwire6346 net6347 VGND VGND VPWR VPWR net6346 sky130_fd_sc_hd__clkbuf_2
X_24266_ _04124_ _04125_ VGND VGND VPWR VPWR _04126_ sky130_fd_sc_hd__xor2_2
XFILLER_0_121_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21478_ net5383 _01490_ VGND VGND VPWR VPWR _01491_ sky130_fd_sc_hd__nand2_1
Xwire6357 net6353 VGND VGND VPWR VPWR net6357 sky130_fd_sc_hd__buf_1
XFILLER_0_161_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire5623 net5624 VGND VGND VPWR VPWR net5623 sky130_fd_sc_hd__clkbuf_1
Xwire6368 cordic0.slte0.opA\[15\] VGND VGND VPWR VPWR net6368 sky130_fd_sc_hd__buf_1
XFILLER_0_31_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_length2066 _01796_ VGND VGND VPWR VPWR net2066 sky130_fd_sc_hd__clkbuf_2
Xwire6379 net6377 VGND VGND VPWR VPWR net6379 sky130_fd_sc_hd__buf_1
X_23217_ _03060_ _03086_ VGND VGND VPWR VPWR _03087_ sky130_fd_sc_hd__or2_1
Xwire4900 net4901 VGND VGND VPWR VPWR net4900 sky130_fd_sc_hd__buf_1
XFILLER_0_105_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout4849 net4861 VGND VGND VPWR VPWR net4849 sky130_fd_sc_hd__clkbuf_1
X_20429_ _12133_ VGND VGND VPWR VPWR _12224_ sky130_fd_sc_hd__inv_2
Xwire4922 net4920 VGND VGND VPWR VPWR net4922 sky130_fd_sc_hd__buf_1
X_24197_ _04056_ _04057_ VGND VGND VPWR VPWR _04058_ sky130_fd_sc_hd__xor2_2
Xwire5667 net5668 VGND VGND VPWR VPWR net5667 sky130_fd_sc_hd__clkbuf_1
Xwire5678 net5679 VGND VGND VPWR VPWR net5678 sky130_fd_sc_hd__buf_1
X_23148_ _03015_ _03016_ _03017_ VGND VGND VPWR VPWR _03018_ sky130_fd_sc_hd__o21ai_1
Xwire4955 net4945 VGND VGND VPWR VPWR net4955 sky130_fd_sc_hd__clkbuf_1
Xwire4966 net4967 VGND VGND VPWR VPWR net4966 sky130_fd_sc_hd__clkbuf_1
Xwire4977 net4978 VGND VGND VPWR VPWR net4977 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23079_ net4949 net4722 VGND VGND VPWR VPWR _02949_ sky130_fd_sc_hd__nand2_1
X_15970_ net2708 net3416 VGND VGND VPWR VPWR _08038_ sky130_fd_sc_hd__nor2_1
X_14921_ net6610 net7425 matmul0.matmul_stage_inst.a\[6\] net6583 VGND VGND VPWR VPWR
+ _06995_ sky130_fd_sc_hd__a22o_1
Xhold50 matmul0.matmul_stage_inst.c\[10\] VGND VGND VPWR VPWR net9003 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 pid_q.target\[5\] VGND VGND VPWR VPWR net9014 sky130_fd_sc_hd__dlygate4sd3_1
X_17640_ net6689 svm0.tA\[14\] VGND VGND VPWR VPWR _09520_ sky130_fd_sc_hd__and2b_1
Xhold72 cordic0.cos\[8\] VGND VGND VPWR VPWR net9025 sky130_fd_sc_hd__dlygate4sd3_1
X_14852_ _06943_ VGND VGND VPWR VPWR _00197_ sky130_fd_sc_hd__clkbuf_1
Xhold83 matmul0.matmul_stage_inst.b\[6\] VGND VGND VPWR VPWR net9036 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold94 svm0.vC\[4\] VGND VGND VPWR VPWR net9047 sky130_fd_sc_hd__dlygate4sd3_1
X_13803_ net7807 net1568 VGND VGND VPWR VPWR _06071_ sky130_fd_sc_hd__nand2_1
X_17571_ net4003 svm0.tC\[2\] svm0.tC\[1\] net4012 VGND VGND VPWR VPWR _09453_ sky130_fd_sc_hd__o22a_1
X_14783_ matmul0.matmul_stage_inst.c\[13\] _06906_ net3698 VGND VGND VPWR VPWR _06907_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_187_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_55_clk clknet_4_11__leaf_clk VGND VGND VPWR VPWR clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_98_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19310_ net6312 net6338 VGND VGND VPWR VPWR _11147_ sky130_fd_sc_hd__nor2_1
X_13734_ _05867_ net451 _05866_ VGND VGND VPWR VPWR _06003_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16522_ _08570_ _08580_ VGND VGND VPWR VPWR _08582_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19241_ net6288 _11075_ _11077_ VGND VGND VPWR VPWR _11078_ sky130_fd_sc_hd__and3_1
X_13665_ _05869_ _05934_ VGND VGND VPWR VPWR _05935_ sky130_fd_sc_hd__xor2_1
X_16453_ _08512_ _08513_ VGND VGND VPWR VPWR _08514_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12616_ _04888_ VGND VGND VPWR VPWR _04889_ sky130_fd_sc_hd__buf_6
XFILLER_0_6_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15404_ _07345_ _07346_ _07347_ _07477_ VGND VGND VPWR VPWR _07478_ sky130_fd_sc_hd__o22a_2
XFILLER_0_156_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19172_ net2110 net2109 _11008_ VGND VGND VPWR VPWR _11009_ sky130_fd_sc_hd__a21o_1
X_16384_ net976 _08445_ VGND VGND VPWR VPWR _08446_ sky130_fd_sc_hd__xor2_2
X_13596_ _05863_ _05865_ VGND VGND VPWR VPWR _05866_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout7453 net7460 VGND VGND VPWR VPWR net7453 sky130_fd_sc_hd__buf_1
XFILLER_0_137_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15335_ _07073_ net1280 _07407_ VGND VGND VPWR VPWR _07409_ sky130_fd_sc_hd__nand3_1
Xwire8260 net8261 VGND VGND VPWR VPWR net8260 sky130_fd_sc_hd__clkbuf_1
X_18123_ net7092 _09613_ VGND VGND VPWR VPWR _09974_ sky130_fd_sc_hd__nand2_1
Xwire8271 net8272 VGND VGND VPWR VPWR net8271 sky130_fd_sc_hd__clkbuf_1
Xwire8282 net8283 VGND VGND VPWR VPWR net8282 sky130_fd_sc_hd__clkbuf_1
Xwire8293 net8294 VGND VGND VPWR VPWR net8293 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7570 matmul0.b_in\[6\] VGND VGND VPWR VPWR net7570 sky130_fd_sc_hd__clkbuf_1
X_15266_ _07219_ _07339_ VGND VGND VPWR VPWR _07340_ sky130_fd_sc_hd__and2_1
X_18054_ net7097 _09903_ _09904_ VGND VGND VPWR VPWR _09905_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_13_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7581 net7582 VGND VGND VPWR VPWR net7581 sky130_fd_sc_hd__clkbuf_1
Xwire7592 net7593 VGND VGND VPWR VPWR net7592 sky130_fd_sc_hd__clkbuf_1
X_14217_ _06466_ _06475_ VGND VGND VPWR VPWR _06476_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17005_ net7065 VGND VGND VPWR VPWR _08966_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15197_ _07269_ _07270_ VGND VGND VPWR VPWR _07271_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14148_ _06404_ _06408_ VGND VGND VPWR VPWR _06409_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_10_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14079_ net7692 net1314 VGND VGND VPWR VPWR _06342_ sky130_fd_sc_hd__nand2_1
X_18956_ net3216 net3215 VGND VGND VPWR VPWR _10793_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17907_ _09745_ _09757_ VGND VGND VPWR VPWR _09758_ sky130_fd_sc_hd__xor2_1
X_18887_ net352 _10694_ VGND VGND VPWR VPWR _10729_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_175_Right_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17838_ net7059 net7028 VGND VGND VPWR VPWR _09689_ sky130_fd_sc_hd__and2b_1
XFILLER_0_156_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17769_ _09619_ VGND VGND VPWR VPWR _09620_ sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_46_clk clknet_4_14__leaf_clk VGND VGND VPWR VPWR clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_156_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19508_ net2507 _11343_ VGND VGND VPWR VPWR _11345_ sky130_fd_sc_hd__and2b_1
XFILLER_0_76_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20780_ _12549_ _12550_ VGND VGND VPWR VPWR _12551_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19439_ net3893 _10983_ _10854_ VGND VGND VPWR VPWR _11276_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22450_ net2057 _02375_ VGND VGND VPWR VPWR _02452_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21401_ net3789 net3118 _01306_ VGND VGND VPWR VPWR _01415_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22381_ _02382_ _02383_ VGND VGND VPWR VPWR _02384_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24120_ net4624 net4802 VGND VGND VPWR VPWR _03982_ sky130_fd_sc_hd__nand2_1
X_21332_ _01344_ _01345_ VGND VGND VPWR VPWR _01346_ sky130_fd_sc_hd__xnor2_1
X_24051_ _03911_ _03913_ VGND VGND VPWR VPWR _03914_ sky130_fd_sc_hd__nand2_1
Xwire4207 _06974_ VGND VGND VPWR VPWR net4207 sky130_fd_sc_hd__buf_1
X_21263_ net5803 net5535 VGND VGND VPWR VPWR _01278_ sky130_fd_sc_hd__nand2_1
Xwire4218 _06965_ VGND VGND VPWR VPWR net4218 sky130_fd_sc_hd__clkbuf_1
Xwire4229 net4230 VGND VGND VPWR VPWR net4229 sky130_fd_sc_hd__clkbuf_1
X_23002_ net5069 net4629 VGND VGND VPWR VPWR _02872_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20214_ _12036_ VGND VGND VPWR VPWR _00467_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3517 net3518 VGND VGND VPWR VPWR net3517 sky130_fd_sc_hd__buf_1
X_21194_ net5617 _01195_ _01208_ _01209_ _01189_ VGND VGND VPWR VPWR _01210_ sky130_fd_sc_hd__a32o_1
Xwire3528 net3529 VGND VGND VPWR VPWR net3528 sky130_fd_sc_hd__buf_1
Xwire3539 net3540 VGND VGND VPWR VPWR net3539 sky130_fd_sc_hd__buf_1
XFILLER_0_21_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2805 net2806 VGND VGND VPWR VPWR net2805 sky130_fd_sc_hd__buf_1
X_20145_ net3137 _11292_ VGND VGND VPWR VPWR _11972_ sky130_fd_sc_hd__nand2_1
Xwire2816 net2817 VGND VGND VPWR VPWR net2816 sky130_fd_sc_hd__buf_1
Xwire2838 _07041_ VGND VGND VPWR VPWR net2838 sky130_fd_sc_hd__buf_1
X_24953_ _04729_ VGND VGND VPWR VPWR _00758_ sky130_fd_sc_hd__clkbuf_1
X_20076_ _11850_ _11868_ _11806_ VGND VGND VPWR VPWR _11905_ sky130_fd_sc_hd__a21bo_1
X_23904_ net7526 _03675_ net408 net7466 net1016 VGND VGND VPWR VPWR _03769_ sky130_fd_sc_hd__a221o_1
X_24884_ _04680_ net4594 net1996 VGND VGND VPWR VPWR _04681_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_142_Right_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_196_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23835_ _03698_ _03699_ VGND VGND VPWR VPWR _03700_ sky130_fd_sc_hd__xnor2_2
Xclkbuf_leaf_37_clk clknet_4_12__leaf_clk VGND VGND VPWR VPWR clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_16
X_23766_ _03493_ net2413 _03496_ VGND VGND VPWR VPWR _03632_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_71_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6833 net6831 VGND VGND VPWR VPWR net6833 sky130_fd_sc_hd__clkbuf_2
X_20978_ _00976_ _00993_ VGND VGND VPWR VPWR _00994_ sky130_fd_sc_hd__xor2_1
X_25505_ clknet_leaf_39_clk _00385_ net8770 VGND VGND VPWR VPWR svm0.delta\[10\] sky130_fd_sc_hd__dfrtp_1
X_22717_ net3718 net97 VGND VGND VPWR VPWR _02653_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_109_Left_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23697_ _03559_ _03563_ VGND VGND VPWR VPWR _03564_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13450_ _05612_ _05721_ _05722_ VGND VGND VPWR VPWR _05723_ sky130_fd_sc_hd__a21o_1
Xmax_length6899 net6900 VGND VGND VPWR VPWR net6899 sky130_fd_sc_hd__clkbuf_1
X_25436_ clknet_leaf_97_clk _00319_ net8399 VGND VGND VPWR VPWR matmul0.sin\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22648_ _00882_ net3077 VGND VGND VPWR VPWR _02609_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13381_ _05652_ _05653_ VGND VGND VPWR VPWR _05654_ sky130_fd_sc_hd__xnor2_1
X_25367_ clknet_leaf_81_clk _00250_ net8496 VGND VGND VPWR VPWR matmul0.alpha_pass\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_22579_ net3769 _02557_ _02558_ VGND VGND VPWR VPWR _02559_ sky130_fd_sc_hd__and3_1
Xwire6110 net6111 VGND VGND VPWR VPWR net6110 sky130_fd_sc_hd__buf_1
XFILLER_0_35_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15120_ net4206 net4203 VGND VGND VPWR VPWR _07194_ sky130_fd_sc_hd__or2_1
X_24318_ pid_q.curr_error\[9\] VGND VGND VPWR VPWR _04178_ sky130_fd_sc_hd__inv_2
Xwire6121 net6118 VGND VGND VPWR VPWR net6121 sky130_fd_sc_hd__buf_1
XFILLER_0_50_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout4602 net4609 VGND VGND VPWR VPWR net4602 sky130_fd_sc_hd__clkbuf_1
Xwire6143 net6144 VGND VGND VPWR VPWR net6143 sky130_fd_sc_hd__clkbuf_1
X_25298_ clknet_leaf_88_clk _00181_ net8431 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.d\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6154 net6153 VGND VGND VPWR VPWR net6154 sky130_fd_sc_hd__buf_1
Xwire5420 net5421 VGND VGND VPWR VPWR net5420 sky130_fd_sc_hd__buf_1
Xwire6165 net6166 VGND VGND VPWR VPWR net6165 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5431 net5432 VGND VGND VPWR VPWR net5431 sky130_fd_sc_hd__buf_1
X_15051_ net3560 VGND VGND VPWR VPWR _07125_ sky130_fd_sc_hd__buf_1
X_24249_ _04109_ _04031_ pid_q.prev_error\[8\] VGND VGND VPWR VPWR _04110_ sky130_fd_sc_hd__a21bo_1
Xfanout4646 net4668 VGND VGND VPWR VPWR net4646 sky130_fd_sc_hd__clkbuf_1
Xwire5442 net5443 VGND VGND VPWR VPWR net5442 sky130_fd_sc_hd__clkbuf_1
Xwire6187 net6188 VGND VGND VPWR VPWR net6187 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_160_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6198 net6199 VGND VGND VPWR VPWR net6198 sky130_fd_sc_hd__buf_1
XFILLER_0_31_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14002_ _06165_ _06209_ VGND VGND VPWR VPWR _06267_ sky130_fd_sc_hd__nand2_1
Xwire5464 net5465 VGND VGND VPWR VPWR net5464 sky130_fd_sc_hd__buf_1
XFILLER_0_120_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4730 net4731 VGND VGND VPWR VPWR net4730 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_118_Left_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire5486 net5488 VGND VGND VPWR VPWR net5486 sky130_fd_sc_hd__clkbuf_1
Xwire4752 net4744 VGND VGND VPWR VPWR net4752 sky130_fd_sc_hd__clkbuf_1
Xwire4763 net4765 VGND VGND VPWR VPWR net4763 sky130_fd_sc_hd__clkbuf_1
Xwire4774 net4775 VGND VGND VPWR VPWR net4774 sky130_fd_sc_hd__clkbuf_1
X_18810_ _10596_ _10598_ _10653_ VGND VGND VPWR VPWR _10654_ sky130_fd_sc_hd__o21ai_2
Xwire4785 net4786 VGND VGND VPWR VPWR net4785 sky130_fd_sc_hd__clkbuf_1
Xwire4796 net4797 VGND VGND VPWR VPWR net4796 sky130_fd_sc_hd__buf_1
X_19790_ net6088 net3136 _11588_ net2100 VGND VGND VPWR VPWR _11624_ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18741_ _10579_ _10585_ VGND VGND VPWR VPWR _10586_ sky130_fd_sc_hd__xnor2_1
X_15953_ net2753 net2653 VGND VGND VPWR VPWR _08021_ sky130_fd_sc_hd__nor2_1
Xinput140 pid_q_data[4] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_1
X_14904_ net4207 net4203 net4198 net4197 VGND VGND VPWR VPWR _06978_ sky130_fd_sc_hd__o22a_1
X_18672_ _10501_ _10506_ _10500_ VGND VGND VPWR VPWR _10518_ sky130_fd_sc_hd__a21oi_1
X_15884_ net2810 _07686_ VGND VGND VPWR VPWR _07953_ sky130_fd_sc_hd__nand2_1
X_17623_ net4033 svm0.tB\[0\] _09502_ VGND VGND VPWR VPWR _09504_ sky130_fd_sc_hd__o21a_1
X_14835_ _06934_ VGND VGND VPWR VPWR _00189_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_28_clk clknet_4_9__leaf_clk VGND VGND VPWR VPWR clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_187_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17554_ svm0.tC\[4\] net4010 net6728 _09435_ VGND VGND VPWR VPWR _09436_ sky130_fd_sc_hd__o2bb2a_1
XPHY_EDGE_ROW_127_Left_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14766_ _06826_ net7149 _06847_ VGND VGND VPWR VPWR _06894_ sky130_fd_sc_hd__nand3_1
X_16505_ net2791 net2772 _08564_ VGND VGND VPWR VPWR _08565_ sky130_fd_sc_hd__a21o_1
X_13717_ net7831 net1317 _05882_ _05884_ VGND VGND VPWR VPWR _05986_ sky130_fd_sc_hd__a22o_1
X_17485_ net6717 _09374_ _09375_ _09373_ VGND VGND VPWR VPWR _00398_ sky130_fd_sc_hd__a22o_1
X_14697_ net7453 _06842_ VGND VGND VPWR VPWR _06843_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19224_ net3890 VGND VGND VPWR VPWR _11061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16436_ net723 _08478_ VGND VGND VPWR VPWR _08497_ sky130_fd_sc_hd__and2_1
XFILLER_0_186_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13648_ _05916_ _05917_ VGND VGND VPWR VPWR _05918_ sky130_fd_sc_hd__and2b_1
XFILLER_0_144_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19155_ net3184 _10991_ _10876_ VGND VGND VPWR VPWR _10992_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13579_ _05781_ _05849_ VGND VGND VPWR VPWR _05850_ sky130_fd_sc_hd__or2b_1
X_16367_ _08381_ _08429_ VGND VGND VPWR VPWR _08430_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire8090 net8091 VGND VGND VPWR VPWR net8090 sky130_fd_sc_hd__clkbuf_1
X_18106_ net3234 _09956_ VGND VGND VPWR VPWR _09957_ sky130_fd_sc_hd__xnor2_1
X_15318_ _07388_ _07391_ VGND VGND VPWR VPWR _07392_ sky130_fd_sc_hd__xnor2_1
X_19086_ net3894 net6321 VGND VGND VPWR VPWR _10923_ sky130_fd_sc_hd__nand2_1
X_16298_ _08297_ _08361_ VGND VGND VPWR VPWR _08362_ sky130_fd_sc_hd__and2b_1
XFILLER_0_78_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_136_Left_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18037_ net2555 net7004 net3237 VGND VGND VPWR VPWR _09888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15249_ _07315_ _07318_ _07322_ VGND VGND VPWR VPWR _07323_ sky130_fd_sc_hd__a21o_1
XFILLER_0_111_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19988_ _11812_ _11818_ VGND VGND VPWR VPWR _11819_ sky130_fd_sc_hd__xnor2_1
X_18939_ _10763_ _10777_ VGND VGND VPWR VPWR _10778_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21950_ net2064 net1718 VGND VGND VPWR VPWR _01958_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20901_ net5513 VGND VGND VPWR VPWR _00917_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_145_Left_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21881_ _01780_ _01790_ _01889_ VGND VGND VPWR VPWR _01890_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_19_clk clknet_4_13__leaf_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23620_ _03465_ _03463_ net1020 VGND VGND VPWR VPWR _03487_ sky130_fd_sc_hd__o21a_1
X_20832_ _12548_ _12549_ _00847_ VGND VGND VPWR VPWR _00848_ sky130_fd_sc_hd__a21o_1
XFILLER_0_193_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23551_ _03322_ _03323_ _03418_ VGND VGND VPWR VPWR _03419_ sky130_fd_sc_hd__a21oi_2
X_20763_ _12530_ net2485 VGND VGND VPWR VPWR _12534_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22502_ _02447_ _02502_ VGND VGND VPWR VPWR _02503_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23482_ net4677 net4920 VGND VGND VPWR VPWR _03351_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20694_ _12142_ _12468_ net8060 VGND VGND VPWR VPWR _12469_ sky130_fd_sc_hd__o21ai_1
X_25221_ clknet_leaf_60_clk _00110_ net8669 VGND VGND VPWR VPWR svm0.vC\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire708 _11669_ VGND VGND VPWR VPWR net708 sky130_fd_sc_hd__clkbuf_2
X_22433_ _02229_ _02300_ _02433_ VGND VGND VPWR VPWR _02435_ sky130_fd_sc_hd__o21ai_1
Xwire719 _10023_ VGND VGND VPWR VPWR net719 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25152_ clknet_leaf_41_clk _00041_ net8767 VGND VGND VPWR VPWR pid_q.target\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_154_Left_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22364_ _02358_ _02366_ VGND VGND VPWR VPWR _02367_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24103_ net4521 net4953 VGND VGND VPWR VPWR _03965_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21315_ _01328_ _01329_ VGND VGND VPWR VPWR _01330_ sky130_fd_sc_hd__and2b_1
X_25083_ net4406 net1633 net235 net1629 _04828_ VGND VGND VPWR VPWR _00789_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4004 _09426_ VGND VGND VPWR VPWR net4004 sky130_fd_sc_hd__buf_1
X_22295_ _02215_ _02216_ _02298_ VGND VGND VPWR VPWR _02299_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_4_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4015 _09257_ VGND VGND VPWR VPWR net4015 sky130_fd_sc_hd__buf_1
XFILLER_0_103_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire4026 _09223_ VGND VGND VPWR VPWR net4026 sky130_fd_sc_hd__buf_1
X_24034_ _03893_ _03896_ VGND VGND VPWR VPWR _03897_ sky130_fd_sc_hd__xnor2_2
Xwire4037 _09054_ VGND VGND VPWR VPWR net4037 sky130_fd_sc_hd__buf_1
X_21246_ _01257_ _01260_ VGND VGND VPWR VPWR _01261_ sky130_fd_sc_hd__xnor2_2
Xwire4048 _08954_ VGND VGND VPWR VPWR net4048 sky130_fd_sc_hd__buf_1
XFILLER_0_13_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire3303 net3304 VGND VGND VPWR VPWR net3303 sky130_fd_sc_hd__clkbuf_1
Xwire3314 _09031_ VGND VGND VPWR VPWR net3314 sky130_fd_sc_hd__clkbuf_2
Xwire4059 _08832_ VGND VGND VPWR VPWR net4059 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3325 net3326 VGND VGND VPWR VPWR net3325 sky130_fd_sc_hd__clkbuf_2
Xwire3336 net3337 VGND VGND VPWR VPWR net3336 sky130_fd_sc_hd__buf_1
X_21177_ _01150_ _01151_ VGND VGND VPWR VPWR _01193_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3347 net3348 VGND VGND VPWR VPWR net3347 sky130_fd_sc_hd__buf_1
Xwire3358 net3359 VGND VGND VPWR VPWR net3358 sky130_fd_sc_hd__clkbuf_1
Xwire2613 _08669_ VGND VGND VPWR VPWR net2613 sky130_fd_sc_hd__buf_1
Xwire3369 net3370 VGND VGND VPWR VPWR net3369 sky130_fd_sc_hd__buf_1
Xwire2635 net2636 VGND VGND VPWR VPWR net2635 sky130_fd_sc_hd__buf_1
Xwire1901 _07033_ VGND VGND VPWR VPWR net1901 sky130_fd_sc_hd__buf_1
Xwire2646 net2647 VGND VGND VPWR VPWR net2646 sky130_fd_sc_hd__dlymetal6s2s_1
X_20128_ _11954_ _11955_ VGND VGND VPWR VPWR _11956_ sky130_fd_sc_hd__nor2_1
Xwire1912 net1913 VGND VGND VPWR VPWR net1912 sky130_fd_sc_hd__clkbuf_1
Xwire1923 _05946_ VGND VGND VPWR VPWR net1923 sky130_fd_sc_hd__buf_1
Xwire2668 net2669 VGND VGND VPWR VPWR net2668 sky130_fd_sc_hd__buf_1
Xwire1934 net1937 VGND VGND VPWR VPWR net1934 sky130_fd_sc_hd__clkbuf_1
Xwire2679 net2680 VGND VGND VPWR VPWR net2679 sky130_fd_sc_hd__buf_1
Xwire1945 _05579_ VGND VGND VPWR VPWR net1945 sky130_fd_sc_hd__buf_1
X_12950_ _05008_ _05017_ VGND VGND VPWR VPWR _05223_ sky130_fd_sc_hd__xnor2_1
X_24936_ net8868 net144 VGND VGND VPWR VPWR _04718_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_163_Left_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire1956 _05110_ VGND VGND VPWR VPWR net1956 sky130_fd_sc_hd__clkbuf_1
X_20059_ net6126 net6063 net3140 VGND VGND VPWR VPWR _11888_ sky130_fd_sc_hd__and3_1
Xwire1967 _04932_ VGND VGND VPWR VPWR net1967 sky130_fd_sc_hd__buf_1
Xwire1978 net1979 VGND VGND VPWR VPWR net1978 sky130_fd_sc_hd__buf_1
Xwire1989 net1990 VGND VGND VPWR VPWR net1989 sky130_fd_sc_hd__buf_1
X_12881_ net1336 _05100_ _05093_ VGND VGND VPWR VPWR _05154_ sky130_fd_sc_hd__a21oi_1
X_24867_ _04669_ VGND VGND VPWR VPWR _00732_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14620_ _06788_ _06790_ VGND VGND VPWR VPWR _06791_ sky130_fd_sc_hd__and2_1
X_23818_ net4560 net4957 VGND VGND VPWR VPWR _03683_ sky130_fd_sc_hd__nand2_1
X_24798_ net2883 _04621_ _04622_ VGND VGND VPWR VPWR _04623_ sky130_fd_sc_hd__or3_1
Xmax_length7375 matmul0.matmul_stage_inst.mult2\[13\] VGND VGND VPWR VPWR net7375
+ sky130_fd_sc_hd__buf_1
XFILLER_0_185_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14551_ _06711_ _06728_ net3639 VGND VGND VPWR VPWR _06729_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23749_ _03524_ _03537_ _03538_ VGND VGND VPWR VPWR _03615_ sky130_fd_sc_hd__o21ai_1
Xmax_length7397 matmul0.matmul_stage_inst.e\[2\] VGND VGND VPWR VPWR net7397 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13502_ net367 _05774_ VGND VGND VPWR VPWR _05775_ sky130_fd_sc_hd__xor2_1
Xmax_length6685 svm0.counter\[15\] VGND VGND VPWR VPWR net6685 sky130_fd_sc_hd__clkbuf_2
X_17270_ net2159 net220 net1797 net9093 VGND VGND VPWR VPWR _00364_ sky130_fd_sc_hd__a22o_1
XFILLER_0_193_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14482_ _06657_ _06663_ _06666_ _06659_ VGND VGND VPWR VPWR _06667_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_83_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length5962 net5963 VGND VGND VPWR VPWR net5962 sky130_fd_sc_hd__clkbuf_1
X_13433_ _05607_ _05610_ _05705_ VGND VGND VPWR VPWR _05706_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16221_ _08283_ _08285_ VGND VGND VPWR VPWR _08286_ sky130_fd_sc_hd__nor2_1
XFILLER_0_192_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25419_ clknet_leaf_90_clk _00302_ net8424 VGND VGND VPWR VPWR matmul0.cos\[6\] sky130_fd_sc_hd__dfrtp_1
Xfanout5111 net5135 VGND VGND VPWR VPWR net5111 sky130_fd_sc_hd__buf_1
X_16152_ _08114_ _08116_ net2733 net2223 VGND VGND VPWR VPWR _08218_ sky130_fd_sc_hd__a211oi_1
X_13364_ _05543_ net1136 net1137 VGND VGND VPWR VPWR _05637_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_106_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15103_ net4135 net4128 net4123 net4118 VGND VGND VPWR VPWR _07177_ sky130_fd_sc_hd__o22a_1
X_16083_ _08138_ _08149_ VGND VGND VPWR VPWR _08150_ sky130_fd_sc_hd__xor2_2
X_13295_ _05561_ _05558_ VGND VGND VPWR VPWR _05568_ sky130_fd_sc_hd__and2b_1
XFILLER_0_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5250 net5251 VGND VGND VPWR VPWR net5250 sky130_fd_sc_hd__buf_1
X_19911_ net2097 _11696_ net1412 VGND VGND VPWR VPWR _11743_ sky130_fd_sc_hd__a21o_1
X_15034_ net3495 VGND VGND VPWR VPWR _07108_ sky130_fd_sc_hd__clkbuf_1
Xwire5261 net5262 VGND VGND VPWR VPWR net5261 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire5272 matmul0.beta_pass\[5\] VGND VGND VPWR VPWR net5272 sky130_fd_sc_hd__buf_1
Xfanout4487 net4493 VGND VGND VPWR VPWR net4487 sky130_fd_sc_hd__buf_1
Xwire5283 net5284 VGND VGND VPWR VPWR net5283 sky130_fd_sc_hd__buf_1
Xwire5294 net5296 VGND VGND VPWR VPWR net5294 sky130_fd_sc_hd__buf_1
XFILLER_0_43_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4560 net4561 VGND VGND VPWR VPWR net4560 sky130_fd_sc_hd__buf_1
Xfanout4498 net4509 VGND VGND VPWR VPWR net4498 sky130_fd_sc_hd__buf_1
X_19842_ net1747 _11651_ VGND VGND VPWR VPWR _11675_ sky130_fd_sc_hd__or2b_1
Xwire4571 net4574 VGND VGND VPWR VPWR net4571 sky130_fd_sc_hd__clkbuf_1
Xwire4582 net4583 VGND VGND VPWR VPWR net4582 sky130_fd_sc_hd__clkbuf_1
Xwire4593 net4588 VGND VGND VPWR VPWR net4593 sky130_fd_sc_hd__clkbuf_1
Xwire3881 _10995_ VGND VGND VPWR VPWR net3881 sky130_fd_sc_hd__buf_1
X_19773_ _11534_ net1057 _11607_ VGND VGND VPWR VPWR _11608_ sky130_fd_sc_hd__o21a_1
X_16985_ _08828_ _08928_ net4062 VGND VGND VPWR VPWR _08947_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18724_ _10552_ _10559_ VGND VGND VPWR VPWR _10569_ sky130_fd_sc_hd__nor2_1
X_15936_ _07911_ _07912_ VGND VGND VPWR VPWR _08005_ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_188_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18655_ _10500_ _10501_ VGND VGND VPWR VPWR _10502_ sky130_fd_sc_hd__and2b_1
X_15867_ net3599 VGND VGND VPWR VPWR _07936_ sky130_fd_sc_hd__buf_1
XFILLER_0_189_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17606_ _09392_ svm0.tB\[11\] _09486_ net6706 VGND VGND VPWR VPWR _09487_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14818_ net9087 _06869_ _06819_ _06911_ VGND VGND VPWR VPWR _00181_ sky130_fd_sc_hd__a22o_1
X_18586_ net6900 net3981 VGND VGND VPWR VPWR _10434_ sky130_fd_sc_hd__nand2_1
X_15798_ _07865_ _07867_ VGND VGND VPWR VPWR _07868_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_176_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17537_ net9041 _09418_ _09419_ VGND VGND VPWR VPWR _00406_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_157_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14749_ net9017 net2857 _06879_ _06881_ VGND VGND VPWR VPWR _00156_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17468_ net4014 _09360_ VGND VGND VPWR VPWR _09361_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19207_ _11043_ _11033_ _11039_ VGND VGND VPWR VPWR _11044_ sky130_fd_sc_hd__or3_1
XFILLER_0_27_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16419_ net490 net571 VGND VGND VPWR VPWR _08481_ sky130_fd_sc_hd__nand2_1
X_17399_ net2573 net1461 VGND VGND VPWR VPWR _09305_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout7080 cordic0.vec\[1\]\[3\] VGND VGND VPWR VPWR net7080 sky130_fd_sc_hd__buf_1
X_19138_ net6184 net6153 VGND VGND VPWR VPWR _10975_ sky130_fd_sc_hd__nand2_1
XFILLER_0_171_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19069_ _10893_ _10897_ _10905_ VGND VGND VPWR VPWR _10906_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_8_clk clknet_4_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_70_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_196_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21100_ _01099_ _01112_ VGND VGND VPWR VPWR _01116_ sky130_fd_sc_hd__nor2_1
X_22080_ net2477 net1044 VGND VGND VPWR VPWR _02087_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21031_ _00991_ _00983_ VGND VGND VPWR VPWR _01047_ sky130_fd_sc_hd__xor2_1
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1208 net1209 VGND VGND VPWR VPWR net1208 sky130_fd_sc_hd__buf_1
Xwire1219 _09580_ VGND VGND VPWR VPWR net1219 sky130_fd_sc_hd__buf_1
X_25770_ clknet_leaf_27_clk _00643_ net8650 VGND VGND VPWR VPWR pid_d.out\[11\] sky130_fd_sc_hd__dfrtp_1
X_22982_ net5219 net528 net6568 VGND VGND VPWR VPWR _02859_ sky130_fd_sc_hd__mux2_1
X_24721_ net5283 VGND VGND VPWR VPWR _04555_ sky130_fd_sc_hd__inv_2
X_21933_ _01836_ _01841_ _01940_ VGND VGND VPWR VPWR _01941_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24652_ _04329_ _04506_ net9015 _02867_ VGND VGND VPWR VPWR _00680_ sky130_fd_sc_hd__a2bb2o_1
X_21864_ net5375 VGND VGND VPWR VPWR _01873_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23603_ _03379_ net745 _03318_ VGND VGND VPWR VPWR _03471_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_length5203 matmul0.beta_pass\[13\] VGND VGND VPWR VPWR net5203 sky130_fd_sc_hd__buf_1
X_20815_ _00825_ _00830_ VGND VGND VPWR VPWR _00831_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_195_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24583_ _04423_ _04438_ VGND VGND VPWR VPWR _04439_ sky130_fd_sc_hd__xor2_1
X_21795_ _01718_ _01720_ _01652_ VGND VGND VPWR VPWR _01805_ sky130_fd_sc_hd__a21o_1
Xwire8804 net8805 VGND VGND VPWR VPWR net8804 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23534_ net4532 net5108 VGND VGND VPWR VPWR _03402_ sky130_fd_sc_hd__nand2_1
Xwire8815 net8816 VGND VGND VPWR VPWR net8815 sky130_fd_sc_hd__clkbuf_1
X_20746_ _12515_ _12516_ VGND VGND VPWR VPWR _12517_ sky130_fd_sc_hd__xnor2_1
Xwire8826 net8814 VGND VGND VPWR VPWR net8826 sky130_fd_sc_hd__buf_1
Xwire8837 net8838 VGND VGND VPWR VPWR net8837 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8848 net8849 VGND VGND VPWR VPWR net8848 sky130_fd_sc_hd__clkbuf_1
Xwire8859 net8860 VGND VGND VPWR VPWR net8859 sky130_fd_sc_hd__clkbuf_1
Xwire505 net506 VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23465_ _03328_ net2426 VGND VGND VPWR VPWR _03334_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_174_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length4568 net4569 VGND VGND VPWR VPWR net4568 sky130_fd_sc_hd__clkbuf_1
Xwire516 _03474_ VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__clkbuf_1
X_20677_ net1077 _12452_ VGND VGND VPWR VPWR _12453_ sky130_fd_sc_hd__nand2_1
Xwire527 _09106_ VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__buf_1
Xwire538 net539 VGND VGND VPWR VPWR net538 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25204_ clknet_leaf_57_clk _00093_ net8715 VGND VGND VPWR VPWR matmul0.b_in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22416_ _02352_ _02353_ _02354_ VGND VGND VPWR VPWR _02418_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire549 net550 VGND VGND VPWR VPWR net549 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_190_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23396_ net5124 net4550 VGND VGND VPWR VPWR _03266_ sky130_fd_sc_hd__nand2_1
X_25135_ clknet_leaf_52_clk _00024_ net8806 VGND VGND VPWR VPWR svm0.tC\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22347_ net5378 _02349_ VGND VGND VPWR VPWR _02350_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13080_ net2303 _05349_ _05350_ _05352_ VGND VGND VPWR VPWR _05353_ sky130_fd_sc_hd__a31o_1
X_25066_ net510 net238 VGND VGND VPWR VPWR _04814_ sky130_fd_sc_hd__or2_1
X_22278_ net2052 _02219_ _02214_ VGND VGND VPWR VPWR _02282_ sky130_fd_sc_hd__a21bo_1
Xwire3100 _02542_ VGND VGND VPWR VPWR net3100 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24017_ net4519 net4971 VGND VGND VPWR VPWR _03880_ sky130_fd_sc_hd__nand2_1
Xwire3111 net3112 VGND VGND VPWR VPWR net3111 sky130_fd_sc_hd__buf_1
Xhold180 pid_q.prev_error\[9\] VGND VGND VPWR VPWR net9133 sky130_fd_sc_hd__dlygate4sd3_1
X_21229_ net4298 _01244_ VGND VGND VPWR VPWR _01245_ sky130_fd_sc_hd__nor2_1
Xwire3122 net3123 VGND VGND VPWR VPWR net3122 sky130_fd_sc_hd__clkbuf_2
Xhold191 pid_q.prev_error\[5\] VGND VGND VPWR VPWR net9144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3144 net3145 VGND VGND VPWR VPWR net3144 sky130_fd_sc_hd__buf_1
Xwire2410 _03962_ VGND VGND VPWR VPWR net2410 sky130_fd_sc_hd__buf_1
XFILLER_0_109_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire3155 net3156 VGND VGND VPWR VPWR net3155 sky130_fd_sc_hd__buf_1
Xwire2421 net2422 VGND VGND VPWR VPWR net2421 sky130_fd_sc_hd__clkbuf_1
Xwire3166 net3167 VGND VGND VPWR VPWR net3166 sky130_fd_sc_hd__buf_1
Xwire2432 _02937_ VGND VGND VPWR VPWR net2432 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire3177 _11061_ VGND VGND VPWR VPWR net3177 sky130_fd_sc_hd__buf_1
Xwire2443 net2444 VGND VGND VPWR VPWR net2443 sky130_fd_sc_hd__clkbuf_1
Xwire3188 _10962_ VGND VGND VPWR VPWR net3188 sky130_fd_sc_hd__clkbuf_1
Xwire2454 _02620_ VGND VGND VPWR VPWR net2454 sky130_fd_sc_hd__buf_1
Xwire3199 net3200 VGND VGND VPWR VPWR net3199 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire1720 _01700_ VGND VGND VPWR VPWR net1720 sky130_fd_sc_hd__buf_1
Xwire2465 net2466 VGND VGND VPWR VPWR net2465 sky130_fd_sc_hd__buf_1
Xwire1731 _01048_ VGND VGND VPWR VPWR net1731 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_176_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2476 net2477 VGND VGND VPWR VPWR net2476 sky130_fd_sc_hd__buf_1
X_16770_ _08774_ VGND VGND VPWR VPWR _00284_ sky130_fd_sc_hd__clkbuf_1
X_13982_ _06244_ net1305 VGND VGND VPWR VPWR _06247_ sky130_fd_sc_hd__nand2_1
Xwire2487 net2488 VGND VGND VPWR VPWR net2487 sky130_fd_sc_hd__buf_1
Xwire1742 net1743 VGND VGND VPWR VPWR net1742 sky130_fd_sc_hd__buf_1
Xwire1753 net1754 VGND VGND VPWR VPWR net1753 sky130_fd_sc_hd__buf_1
Xwire2498 net2499 VGND VGND VPWR VPWR net2498 sky130_fd_sc_hd__buf_1
Xwire1764 _10428_ VGND VGND VPWR VPWR net1764 sky130_fd_sc_hd__clkbuf_1
X_15721_ _07783_ _07791_ VGND VGND VPWR VPWR _07792_ sky130_fd_sc_hd__xnor2_2
Xwire1775 _10153_ VGND VGND VPWR VPWR net1775 sky130_fd_sc_hd__dlymetal6s2s_1
X_24919_ pid_q.ki\[2\] _04706_ net1360 VGND VGND VPWR VPWR _04707_ sky130_fd_sc_hd__mux2_1
X_12933_ _05126_ net791 VGND VGND VPWR VPWR _05206_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire1786 net1787 VGND VGND VPWR VPWR net1786 sky130_fd_sc_hd__buf_1
X_25899_ clknet_leaf_16_clk _00772_ net8627 VGND VGND VPWR VPWR pid_q.kp\[11\] sky130_fd_sc_hd__dfrtp_1
Xwire1797 net1798 VGND VGND VPWR VPWR net1797 sky130_fd_sc_hd__clkbuf_2
X_18440_ _10288_ _10289_ VGND VGND VPWR VPWR _10290_ sky130_fd_sc_hd__or2_1
X_15652_ net3393 VGND VGND VPWR VPWR _07724_ sky130_fd_sc_hd__buf_1
X_12864_ net7931 _05057_ _05136_ VGND VGND VPWR VPWR _05137_ sky130_fd_sc_hd__and3_1
Xmax_length7150 matmul0.sin\[9\] VGND VGND VPWR VPWR net7150 sky130_fd_sc_hd__clkbuf_1
X_14603_ _06774_ _06775_ VGND VGND VPWR VPWR _06776_ sky130_fd_sc_hd__xnor2_1
X_18371_ net6882 net6854 VGND VGND VPWR VPWR _10222_ sky130_fd_sc_hd__and2b_1
XFILLER_0_157_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12795_ _04935_ _04939_ VGND VGND VPWR VPWR _05068_ sky130_fd_sc_hd__or2_1
X_15583_ net3455 net3556 VGND VGND VPWR VPWR _07655_ sky130_fd_sc_hd__nor2_1
X_17322_ net6737 net7919 VGND VGND VPWR VPWR _09236_ sky130_fd_sc_hd__xor2_1
X_14534_ _06711_ _06712_ net5247 VGND VGND VPWR VPWR _06713_ sky130_fd_sc_hd__a21o_1
XFILLER_0_83_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17253_ _09185_ net187 _09190_ net9080 VGND VGND VPWR VPWR _00351_ sky130_fd_sc_hd__a22o_1
X_14465_ _06531_ VGND VGND VPWR VPWR _06653_ sky130_fd_sc_hd__buf_1
XFILLER_0_154_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16204_ _08177_ _08262_ _08268_ VGND VGND VPWR VPWR _08269_ sky130_fd_sc_hd__o21ai_1
X_13416_ net3678 net3675 VGND VGND VPWR VPWR _05689_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14396_ net8157 net3635 VGND VGND VPWR VPWR _06600_ sky130_fd_sc_hd__and2_1
X_17184_ _09133_ _09134_ VGND VGND VPWR VPWR _09135_ sky130_fd_sc_hd__xor2_1
XFILLER_0_84_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13347_ net7923 _05619_ net2294 net3675 net3679 VGND VGND VPWR VPWR _05620_ sky130_fd_sc_hd__a311oi_2
X_16135_ net1516 _08103_ _08098_ VGND VGND VPWR VPWR _08201_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13278_ _05547_ _05548_ net846 VGND VGND VPWR VPWR _05551_ sky130_fd_sc_hd__a21oi_1
X_16066_ net1525 net1258 VGND VGND VPWR VPWR _08133_ sky130_fd_sc_hd__nor2_1
Xwire5080 net5081 VGND VGND VPWR VPWR net5080 sky130_fd_sc_hd__buf_1
X_15017_ net2826 _07078_ _07090_ VGND VGND VPWR VPWR _07091_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4390 pid_d.state\[0\] VGND VGND VPWR VPWR net4390 sky130_fd_sc_hd__buf_1
X_19825_ _11657_ _11658_ net3291 VGND VGND VPWR VPWR _11659_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19756_ net6072 _11587_ _11589_ _11590_ VGND VGND VPWR VPWR _11591_ sky130_fd_sc_hd__a31o_1
X_16968_ _08846_ _08930_ net6525 VGND VGND VPWR VPWR _08931_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18707_ net6792 net2539 _10487_ net6812 VGND VGND VPWR VPWR _10553_ sky130_fd_sc_hd__a2bb2o_1
X_15919_ _07878_ _07886_ _07884_ VGND VGND VPWR VPWR _07988_ sky130_fd_sc_hd__o21a_1
X_19687_ _11519_ _11522_ VGND VGND VPWR VPWR _11523_ sky130_fd_sc_hd__xnor2_1
X_16899_ net6371 _08861_ _08862_ VGND VGND VPWR VPWR _08863_ sky130_fd_sc_hd__a21o_1
XFILLER_0_91_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18638_ net1433 _10484_ VGND VGND VPWR VPWR _10485_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_59_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18569_ net6859 _10282_ _10283_ _10287_ _10416_ VGND VGND VPWR VPWR _10417_ sky130_fd_sc_hd__a32o_1
X_20600_ _12380_ _12381_ VGND VGND VPWR VPWR _12382_ sky130_fd_sc_hd__xnor2_1
X_21580_ net3818 _01490_ VGND VGND VPWR VPWR _01592_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20531_ net3124 _12314_ _12315_ _12316_ net3334 net3332 VGND VGND VPWR VPWR _12317_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_156_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire6709 net6710 VGND VGND VPWR VPWR net6709 sky130_fd_sc_hd__clkbuf_1
X_23250_ _03116_ _03119_ VGND VGND VPWR VPWR _03120_ sky130_fd_sc_hd__or2_1
Xmax_length2407 _04009_ VGND VGND VPWR VPWR net2407 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20462_ cordic0.slte0.opA\[15\] _12250_ _12252_ VGND VGND VPWR VPWR _12254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22201_ _02141_ _02143_ _02205_ VGND VGND VPWR VPWR _02206_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23181_ _03049_ _03050_ VGND VGND VPWR VPWR _03051_ sky130_fd_sc_hd__nand2_1
X_20393_ cordic0.slte0.opA\[9\] VGND VGND VPWR VPWR _12191_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22132_ net5764 net5389 net3779 _02136_ VGND VGND VPWR VPWR _02138_ sky130_fd_sc_hd__a211o_1
XFILLER_0_112_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22063_ net1041 _02069_ VGND VGND VPWR VPWR _02070_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21014_ net2076 _00994_ VGND VGND VPWR VPWR _01030_ sky130_fd_sc_hd__nand2_1
Xwire1005 _05117_ VGND VGND VPWR VPWR net1005 sky130_fd_sc_hd__buf_1
Xwire1016 net1017 VGND VGND VPWR VPWR net1016 sky130_fd_sc_hd__clkbuf_1
Xwire1027 _03375_ VGND VGND VPWR VPWR net1027 sky130_fd_sc_hd__clkbuf_1
X_25822_ clknet_leaf_30_clk _00695_ net8686 VGND VGND VPWR VPWR pid_q.prev_error\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire1038 net1039 VGND VGND VPWR VPWR net1038 sky130_fd_sc_hd__buf_1
Xwire1049 _01480_ VGND VGND VPWR VPWR net1049 sky130_fd_sc_hd__dlymetal6s2s_1
X_25753_ clknet_leaf_12_clk _00626_ net8604 VGND VGND VPWR VPWR pid_d.kp\[11\] sky130_fd_sc_hd__dfrtp_1
X_22965_ _02850_ VGND VGND VPWR VPWR _00649_ sky130_fd_sc_hd__clkbuf_1
X_24704_ net7488 net4000 _04540_ VGND VGND VPWR VPWR _04541_ sky130_fd_sc_hd__and3_1
X_21916_ net599 _01922_ VGND VGND VPWR VPWR _01924_ sky130_fd_sc_hd__nor2_1
X_22896_ net5354 net3103 _02789_ net4328 VGND VGND VPWR VPWR _02790_ sky130_fd_sc_hd__a22o_1
X_25684_ clknet_leaf_0_clk _00557_ net8571 VGND VGND VPWR VPWR pid_d.curr_error\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_179_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24635_ net4491 _04489_ VGND VGND VPWR VPWR _04490_ sky130_fd_sc_hd__nand2_1
X_21847_ _01850_ _01855_ VGND VGND VPWR VPWR _01856_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_33_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout7805 net7814 VGND VGND VPWR VPWR net7805 sky130_fd_sc_hd__clkbuf_1
X_24566_ net2016 _04421_ VGND VGND VPWR VPWR _04422_ sky130_fd_sc_hd__xor2_1
Xwire8601 net8590 VGND VGND VPWR VPWR net8601 sky130_fd_sc_hd__buf_1
X_12580_ _04865_ VGND VGND VPWR VPWR _04866_ sky130_fd_sc_hd__clkbuf_1
Xwire8612 net8613 VGND VGND VPWR VPWR net8612 sky130_fd_sc_hd__clkbuf_1
X_21778_ net2475 _01787_ VGND VGND VPWR VPWR _01788_ sky130_fd_sc_hd__xor2_1
Xwire8634 net8635 VGND VGND VPWR VPWR net8634 sky130_fd_sc_hd__clkbuf_1
Xfanout7827 net7837 VGND VGND VPWR VPWR net7827 sky130_fd_sc_hd__buf_1
Xwire7900 net7901 VGND VGND VPWR VPWR net7900 sky130_fd_sc_hd__clkbuf_1
X_23517_ pid_q.prev_error\[0\] pid_q.curr_error\[0\] _03385_ VGND VGND VPWR VPWR _03386_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_147_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20729_ net3843 VGND VGND VPWR VPWR _12500_ sky130_fd_sc_hd__buf_1
XFILLER_0_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24497_ _04342_ _04353_ VGND VGND VPWR VPWR _04354_ sky130_fd_sc_hd__xnor2_2
Xwire7911 net7912 VGND VGND VPWR VPWR net7911 sky130_fd_sc_hd__clkbuf_1
Xwire8656 net8657 VGND VGND VPWR VPWR net8656 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire302 _10728_ VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__buf_1
XFILLER_0_163_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7922 net7924 VGND VGND VPWR VPWR net7922 sky130_fd_sc_hd__clkbuf_1
Xwire8667 net8668 VGND VGND VPWR VPWR net8667 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_108_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire313 net314 VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__clkbuf_1
Xwire324 net325 VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__buf_1
Xwire7933 net7930 VGND VGND VPWR VPWR net7933 sky130_fd_sc_hd__clkbuf_2
Xwire7944 net7945 VGND VGND VPWR VPWR net7944 sky130_fd_sc_hd__clkbuf_1
Xwire8689 net8690 VGND VGND VPWR VPWR net8689 sky130_fd_sc_hd__buf_1
X_14250_ net4238 _06504_ VGND VGND VPWR VPWR _06505_ sky130_fd_sc_hd__nor2_1
Xwire335 _03851_ VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__clkbuf_1
X_23448_ _03315_ _03316_ VGND VGND VPWR VPWR _03317_ sky130_fd_sc_hd__xnor2_1
Xmax_length3642 net3643 VGND VGND VPWR VPWR net3642 sky130_fd_sc_hd__buf_1
Xwire7955 net7956 VGND VGND VPWR VPWR net7955 sky130_fd_sc_hd__clkbuf_2
Xwire346 net347 VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7966 pid_q.target\[13\] VGND VGND VPWR VPWR net7966 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire357 net358 VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire368 net369 VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__clkbuf_1
Xwire7977 net7978 VGND VGND VPWR VPWR net7977 sky130_fd_sc_hd__clkbuf_1
X_13201_ _05472_ _05362_ _05363_ VGND VGND VPWR VPWR _05474_ sky130_fd_sc_hd__and3_1
Xwire7988 net7989 VGND VGND VPWR VPWR net7988 sky130_fd_sc_hd__clkbuf_1
Xwire379 _03866_ VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__clkbuf_1
Xwire7999 net8000 VGND VGND VPWR VPWR net7999 sky130_fd_sc_hd__clkbuf_1
X_14181_ net7627 net1123 _06407_ VGND VGND VPWR VPWR _06441_ sky130_fd_sc_hd__a21o_1
X_23379_ net4759 net4850 VGND VGND VPWR VPWR _03249_ sky130_fd_sc_hd__nand2_1
Xmax_length2974 net2975 VGND VGND VPWR VPWR net2974 sky130_fd_sc_hd__buf_1
X_13132_ net683 _05401_ _05403_ _05404_ VGND VGND VPWR VPWR _05405_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_103_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25118_ pid_d.prev_int\[6\] net2393 net1993 net9196 VGND VGND VPWR VPWR _00799_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25049_ net9229 net1632 net2395 _04799_ VGND VGND VPWR VPWR _00784_ sky130_fd_sc_hd__a22o_1
X_13063_ _05284_ _05303_ VGND VGND VPWR VPWR _05336_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17940_ net6970 net6933 VGND VGND VPWR VPWR _09791_ sky130_fd_sc_hd__nor2b_1
X_17871_ _09605_ net2141 _09721_ _09610_ VGND VGND VPWR VPWR _09722_ sky130_fd_sc_hd__a211o_1
Xwire2240 _07275_ VGND VGND VPWR VPWR net2240 sky130_fd_sc_hd__clkbuf_1
X_19610_ net6050 net4046 VGND VGND VPWR VPWR _11447_ sky130_fd_sc_hd__nor2_1
Xwire2251 _07130_ VGND VGND VPWR VPWR net2251 sky130_fd_sc_hd__buf_1
X_16822_ _08801_ VGND VGND VPWR VPWR _00309_ sky130_fd_sc_hd__clkbuf_1
Xwire2262 _06825_ VGND VGND VPWR VPWR net2262 sky130_fd_sc_hd__clkbuf_2
Xwire2273 net2274 VGND VGND VPWR VPWR net2273 sky130_fd_sc_hd__clkbuf_1
Xwire2284 _06507_ VGND VGND VPWR VPWR net2284 sky130_fd_sc_hd__buf_1
Xwire2295 _05532_ VGND VGND VPWR VPWR net2295 sky130_fd_sc_hd__clkbuf_1
Xwire1550 _06521_ VGND VGND VPWR VPWR net1550 sky130_fd_sc_hd__buf_1
X_19541_ _10790_ _11377_ VGND VGND VPWR VPWR _11378_ sky130_fd_sc_hd__xnor2_1
Xwire1561 _06175_ VGND VGND VPWR VPWR net1561 sky130_fd_sc_hd__buf_1
X_16753_ _08765_ VGND VGND VPWR VPWR _00276_ sky130_fd_sc_hd__clkbuf_1
X_13965_ net7683 net2954 net3673 VGND VGND VPWR VPWR _06230_ sky130_fd_sc_hd__and3_1
Xwire1572 _05578_ VGND VGND VPWR VPWR net1572 sky130_fd_sc_hd__buf_1
Xwire1583 net1584 VGND VGND VPWR VPWR net1583 sky130_fd_sc_hd__clkbuf_2
Xwire1594 net1595 VGND VGND VPWR VPWR net1594 sky130_fd_sc_hd__buf_1
X_15704_ net1099 _07774_ VGND VGND VPWR VPWR _07775_ sky130_fd_sc_hd__xnor2_2
X_12916_ net7256 _04892_ net3695 VGND VGND VPWR VPWR _05189_ sky130_fd_sc_hd__nand3_1
X_19472_ _11122_ _10984_ _11280_ _11281_ VGND VGND VPWR VPWR _11309_ sky130_fd_sc_hd__a211o_1
X_16684_ _08715_ VGND VGND VPWR VPWR _00257_ sky130_fd_sc_hd__clkbuf_1
X_13896_ _06091_ _06160_ _06161_ VGND VGND VPWR VPWR _06162_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_158_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18423_ net6773 _10211_ VGND VGND VPWR VPWR _10273_ sky130_fd_sc_hd__nand2_1
X_15635_ net1104 net1266 VGND VGND VPWR VPWR _07707_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_100_Left_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12847_ _05038_ _05043_ net1147 VGND VGND VPWR VPWR _05120_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_174_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18354_ _10186_ _10189_ _10204_ VGND VGND VPWR VPWR _10205_ sky130_fd_sc_hd__o21a_1
X_15566_ net674 _07638_ VGND VGND VPWR VPWR _07639_ sky130_fd_sc_hd__xnor2_1
X_12778_ net6678 net5244 net6673 VGND VGND VPWR VPWR _05051_ sky130_fd_sc_hd__and3b_1
XFILLER_0_56_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17305_ net7661 _09213_ net7643 VGND VGND VPWR VPWR _09219_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14517_ net7302 _06695_ _06697_ VGND VGND VPWR VPWR _06698_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_71_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18285_ _10132_ _10135_ VGND VGND VPWR VPWR _10136_ sky130_fd_sc_hd__xnor2_1
X_15497_ net2800 net3440 VGND VGND VPWR VPWR _07570_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17236_ net6759 _08911_ _09182_ VGND VGND VPWR VPWR _09184_ sky130_fd_sc_hd__or3_1
X_14448_ net8174 net4233 VGND VGND VPWR VPWR _06640_ sky130_fd_sc_hd__and2_1
XFILLER_0_141_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17167_ _09068_ _09119_ net6891 VGND VGND VPWR VPWR _09120_ sky130_fd_sc_hd__a21oi_1
X_14379_ _06587_ VGND VGND VPWR VPWR _00080_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire880 _08567_ VGND VGND VPWR VPWR net880 sky130_fd_sc_hd__buf_1
Xwire891 _06864_ VGND VGND VPWR VPWR net891 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16118_ net2206 net1513 VGND VGND VPWR VPWR _08184_ sky130_fd_sc_hd__nor2_1
X_17098_ net2609 net4038 VGND VGND VPWR VPWR _09055_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16049_ net2692 net2637 VGND VGND VPWR VPWR _08116_ sky130_fd_sc_hd__nor2_1
XFILLER_0_177_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19808_ net6214 net6117 VGND VGND VPWR VPWR _11642_ sky130_fd_sc_hd__xnor2_2
X_19739_ net1056 _11573_ VGND VGND VPWR VPWR _11574_ sky130_fd_sc_hd__xor2_2
X_22750_ net4304 net8928 VGND VGND VPWR VPWR _02678_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21701_ net1721 _01599_ _01595_ VGND VGND VPWR VPWR _01712_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_176_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22681_ pid_d.ki\[4\] net2439 net2994 pid_d.kp\[4\] VGND VGND VPWR VPWR _02629_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24420_ _04276_ _04277_ VGND VGND VPWR VPWR _04278_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21632_ pid_d.curr_int\[4\] net3122 net2077 _01643_ VGND VGND VPWR VPWR _00523_ sky130_fd_sc_hd__a22o_1
XFILLER_0_192_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24351_ net4581 net4805 VGND VGND VPWR VPWR _04210_ sky130_fd_sc_hd__nand2_1
X_21563_ _01571_ _01574_ VGND VGND VPWR VPWR _01575_ sky130_fd_sc_hd__xnor2_1
Xwire7207 net7213 VGND VGND VPWR VPWR net7207 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7218 net7219 VGND VGND VPWR VPWR net7218 sky130_fd_sc_hd__buf_1
XFILLER_0_7_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7229 net7230 VGND VGND VPWR VPWR net7229 sky130_fd_sc_hd__clkbuf_1
X_23302_ _03160_ _03165_ _03009_ VGND VGND VPWR VPWR _03172_ sky130_fd_sc_hd__a21o_1
X_20514_ net1484 net2084 net2082 VGND VGND VPWR VPWR _12301_ sky130_fd_sc_hd__a21o_1
XFILLER_0_173_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24282_ net1655 net1654 VGND VGND VPWR VPWR _04142_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21494_ net5427 _01506_ net5416 VGND VGND VPWR VPWR _01507_ sky130_fd_sc_hd__a21o_1
Xwire6528 net6530 VGND VGND VPWR VPWR net6528 sky130_fd_sc_hd__clkbuf_1
X_23233_ _03097_ _03100_ net2430 VGND VGND VPWR VPWR _03103_ sky130_fd_sc_hd__o21a_1
Xwire5805 net5806 VGND VGND VPWR VPWR net5805 sky130_fd_sc_hd__buf_1
Xmax_length2237 net2238 VGND VGND VPWR VPWR net2237 sky130_fd_sc_hd__clkbuf_1
X_20445_ _12235_ _12238_ VGND VGND VPWR VPWR _12239_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length2248 _07156_ VGND VGND VPWR VPWR net2248 sky130_fd_sc_hd__clkbuf_1
Xwire5827 net5828 VGND VGND VPWR VPWR net5827 sky130_fd_sc_hd__clkbuf_1
Xmax_length1514 net1515 VGND VGND VPWR VPWR net1514 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5838 net5830 VGND VGND VPWR VPWR net5838 sky130_fd_sc_hd__buf_1
Xwire5849 net5850 VGND VGND VPWR VPWR net5849 sky130_fd_sc_hd__clkbuf_1
X_23164_ _03016_ _03017_ VGND VGND VPWR VPWR _03034_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20376_ net3313 net1501 VGND VGND VPWR VPWR _12175_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_189_Right_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22115_ _02024_ _02034_ _02120_ VGND VGND VPWR VPWR _02121_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23095_ net1032 _02964_ VGND VGND VPWR VPWR _02965_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_11_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22046_ _01941_ _01952_ _02052_ VGND VGND VPWR VPWR _02053_ sky130_fd_sc_hd__a21oi_1
X_25805_ clknet_leaf_30_clk _00678_ net8673 VGND VGND VPWR VPWR pid_q.curr_int\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_23997_ pid_q.prev_int\[6\] VGND VGND VPWR VPWR _03860_ sky130_fd_sc_hd__inv_2
X_13750_ _05867_ net404 _06013_ VGND VGND VPWR VPWR _06018_ sky130_fd_sc_hd__a21bo_1
X_25736_ clknet_leaf_12_clk _00609_ net8604 VGND VGND VPWR VPWR pid_d.ki\[10\] sky130_fd_sc_hd__dfrtp_1
X_22948_ net551 net549 _02325_ VGND VGND VPWR VPWR _02836_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12701_ net2973 VGND VGND VPWR VPWR _04974_ sky130_fd_sc_hd__clkbuf_1
X_13681_ net1923 _05948_ _05949_ VGND VGND VPWR VPWR _05950_ sky130_fd_sc_hd__or3_1
XFILLER_0_39_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25667_ clknet_leaf_120_clk _00540_ net8397 VGND VGND VPWR VPWR pid_d.prev_error\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22879_ net5360 _02774_ net3066 VGND VGND VPWR VPWR _02775_ sky130_fd_sc_hd__mux2_1
X_15420_ net1865 net1864 VGND VGND VPWR VPWR _07494_ sky130_fd_sc_hd__nor2_1
X_24618_ net1651 _04472_ _04436_ VGND VGND VPWR VPWR _04473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12632_ _04904_ VGND VGND VPWR VPWR _04905_ sky130_fd_sc_hd__clkbuf_1
X_25598_ clknet_leaf_105_clk _00471_ net8354 VGND VGND VPWR VPWR cordic0.slte0.opB\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout8369 net8540 VGND VGND VPWR VPWR net8369 sky130_fd_sc_hd__buf_1
X_15351_ _07319_ net2704 VGND VGND VPWR VPWR _07425_ sky130_fd_sc_hd__xnor2_1
Xwire8431 net8429 VGND VGND VPWR VPWR net8431 sky130_fd_sc_hd__clkbuf_2
X_24549_ net1651 _04403_ _04404_ net2018 VGND VGND VPWR VPWR _04405_ sky130_fd_sc_hd__o31a_1
XFILLER_0_0_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6901 net6905 VGND VGND VPWR VPWR net6901 sky130_fd_sc_hd__clkbuf_2
Xwire8442 net8444 VGND VGND VPWR VPWR net8442 sky130_fd_sc_hd__buf_1
Xfanout7646 net7651 VGND VGND VPWR VPWR net7646 sky130_fd_sc_hd__buf_1
XFILLER_0_53_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14302_ net6446 _06523_ VGND VGND VPWR VPWR _06524_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout6923 net6931 VGND VGND VPWR VPWR net6923 sky130_fd_sc_hd__clkbuf_1
Xwire8464 net8462 VGND VGND VPWR VPWR net8464 sky130_fd_sc_hd__clkbuf_2
Xfanout7679 net7695 VGND VGND VPWR VPWR net7679 sky130_fd_sc_hd__buf_1
Xwire7730 net7731 VGND VGND VPWR VPWR net7730 sky130_fd_sc_hd__buf_1
X_18070_ _09918_ _09920_ VGND VGND VPWR VPWR _09921_ sky130_fd_sc_hd__nor2_1
X_15282_ net1543 _07355_ VGND VGND VPWR VPWR _07356_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout6945 net6958 VGND VGND VPWR VPWR net6945 sky130_fd_sc_hd__buf_1
Xwire8486 net8487 VGND VGND VPWR VPWR net8486 sky130_fd_sc_hd__buf_1
Xwire7752 net7753 VGND VGND VPWR VPWR net7752 sky130_fd_sc_hd__buf_1
Xmax_length4184 net4185 VGND VGND VPWR VPWR net4184 sky130_fd_sc_hd__buf_1
Xwire8497 net8498 VGND VGND VPWR VPWR net8497 sky130_fd_sc_hd__buf_1
Xmax_length4195 net4196 VGND VGND VPWR VPWR net4195 sky130_fd_sc_hd__buf_1
Xwire154 _06489_ VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__buf_1
Xwire7774 net7775 VGND VGND VPWR VPWR net7774 sky130_fd_sc_hd__clkbuf_2
X_17021_ net1917 _08981_ net8043 VGND VGND VPWR VPWR _08982_ sky130_fd_sc_hd__o21a_1
X_14233_ _06466_ _06475_ _06463_ VGND VGND VPWR VPWR _06490_ sky130_fd_sc_hd__a21bo_1
Xwire165 net166 VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_1
Xwire176 net177 VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_1
Xwire187 net188 VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__buf_1
Xwire7796 net7799 VGND VGND VPWR VPWR net7796 sky130_fd_sc_hd__clkbuf_1
Xwire198 net199 VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14164_ _06368_ _06395_ _06394_ VGND VGND VPWR VPWR _06425_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_0_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_156_Right_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13115_ _05266_ _05267_ VGND VGND VPWR VPWR _05388_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14095_ _06356_ _06357_ VGND VGND VPWR VPWR _06358_ sky130_fd_sc_hd__xor2_1
X_18972_ _10793_ _10808_ VGND VGND VPWR VPWR _10809_ sky130_fd_sc_hd__xor2_1
X_13046_ _05318_ _05316_ VGND VGND VPWR VPWR _05319_ sky130_fd_sc_hd__nand2_1
X_17923_ _09761_ _09771_ _09773_ VGND VGND VPWR VPWR _09774_ sky130_fd_sc_hd__o21a_1
XFILLER_0_147_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17854_ _09703_ _09704_ net3256 VGND VGND VPWR VPWR _09705_ sky130_fd_sc_hd__o21a_1
Xwire2070 net2071 VGND VGND VPWR VPWR net2070 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2081 _12318_ VGND VGND VPWR VPWR net2081 sky130_fd_sc_hd__clkbuf_1
X_16805_ net9241 matmul0.cos\[5\] _08792_ VGND VGND VPWR VPWR _08793_ sky130_fd_sc_hd__mux2_1
Xwire2092 _11805_ VGND VGND VPWR VPWR net2092 sky130_fd_sc_hd__buf_1
X_17785_ net7006 net7051 VGND VGND VPWR VPWR _09636_ sky130_fd_sc_hd__or2b_1
X_14997_ net1287 net1286 VGND VGND VPWR VPWR _07071_ sky130_fd_sc_hd__xnor2_1
Xwire1380 _04071_ VGND VGND VPWR VPWR net1380 sky130_fd_sc_hd__buf_1
X_19524_ _11359_ net3158 _11360_ VGND VGND VPWR VPWR _11361_ sky130_fd_sc_hd__o21ai_2
Xwire1391 _01277_ VGND VGND VPWR VPWR net1391 sky130_fd_sc_hd__buf_1
X_16736_ _08756_ VGND VGND VPWR VPWR _00268_ sky130_fd_sc_hd__clkbuf_1
X_13948_ _06159_ _06212_ _06211_ VGND VGND VPWR VPWR _06214_ sky130_fd_sc_hd__a21o_1
X_19455_ net6099 net6050 VGND VGND VPWR VPWR _11292_ sky130_fd_sc_hd__nand2_1
XFILLER_0_158_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16667_ matmul0.matmul_stage_inst.mult2\[7\] matmul0.matmul_stage_inst.mult1\[7\]
+ VGND VGND VPWR VPWR _08701_ sky130_fd_sc_hd__xor2_1
X_13879_ net449 _06144_ _06145_ VGND VGND VPWR VPWR _06146_ sky130_fd_sc_hd__o21a_1
X_18406_ _10205_ net767 VGND VGND VPWR VPWR _10257_ sky130_fd_sc_hd__and2b_1
X_15618_ net4072 _07685_ _07687_ net3527 _07689_ VGND VGND VPWR VPWR _07690_ sky130_fd_sc_hd__a221o_1
X_19386_ net2509 _11157_ VGND VGND VPWR VPWR _11223_ sky130_fd_sc_hd__nand2_1
X_16598_ svm0.delta\[0\] net2614 VGND VGND VPWR VPWR _08649_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18337_ _10121_ net1776 VGND VGND VPWR VPWR _10188_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15549_ net1854 net1853 VGND VGND VPWR VPWR _07622_ sky130_fd_sc_hd__xor2_1
XFILLER_0_44_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18268_ _10117_ _10118_ net2547 VGND VGND VPWR VPWR _10119_ sky130_fd_sc_hd__o21a_1
XFILLER_0_86_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17219_ net2187 _09167_ net3324 VGND VGND VPWR VPWR _09168_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18199_ net3233 _10048_ _10044_ _10046_ VGND VGND VPWR VPWR _10050_ sky130_fd_sc_hd__a211o_1
XFILLER_0_25_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20230_ _12048_ net6415 net2936 VGND VGND VPWR VPWR _12049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20161_ net3126 _11967_ net244 VGND VGND VPWR VPWR _11988_ sky130_fd_sc_hd__or3b_1
XPHY_EDGE_ROW_123_Right_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20092_ net3861 _11915_ _11920_ VGND VGND VPWR VPWR _11921_ sky130_fd_sc_hd__and3_1
XFILLER_0_196_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23920_ net4592 net4905 VGND VGND VPWR VPWR _03784_ sky130_fd_sc_hd__nand2_1
Xmax_length8406 net8407 VGND VGND VPWR VPWR net8406 sky130_fd_sc_hd__buf_1
X_23851_ net4639 net4868 VGND VGND VPWR VPWR _03716_ sky130_fd_sc_hd__nand2_1
Xmax_length8417 net8418 VGND VGND VPWR VPWR net8417 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22802_ pid_d.kp\[13\] _02688_ net2036 VGND VGND VPWR VPWR _02709_ sky130_fd_sc_hd__mux2_1
X_23782_ _03548_ _03550_ VGND VGND VPWR VPWR _03648_ sky130_fd_sc_hd__and2b_1
X_20994_ _01007_ _01008_ net1734 VGND VGND VPWR VPWR _01010_ sky130_fd_sc_hd__a21bo_1
X_25521_ clknet_leaf_47_clk _00401_ net8777 VGND VGND VPWR VPWR svm0.counter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22733_ pid_d.ki\[2\] _02666_ net1688 VGND VGND VPWR VPWR _02667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22664_ net3089 _02598_ _02600_ VGND VGND VPWR VPWR _02617_ sky130_fd_sc_hd__a21oi_1
X_25452_ clknet_leaf_112_clk _00335_ net8341 VGND VGND VPWR VPWR cordic0.vec\[1\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24403_ _04259_ _04260_ VGND VGND VPWR VPWR _04261_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21615_ _01625_ _01626_ VGND VGND VPWR VPWR _01627_ sky130_fd_sc_hd__nand2_1
X_25383_ clknet_leaf_73_clk _00266_ net8476 VGND VGND VPWR VPWR matmul0.b\[2\] sky130_fd_sc_hd__dfrtp_1
X_22595_ pid_d.curr_error\[7\] net1388 net3087 VGND VGND VPWR VPWR _02572_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24334_ _03944_ _04168_ VGND VGND VPWR VPWR _04193_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21546_ net5685 net5592 VGND VGND VPWR VPWR _01558_ sky130_fd_sc_hd__nand2_1
Xwire7037 net7038 VGND VGND VPWR VPWR net7037 sky130_fd_sc_hd__buf_1
Xwire7048 net7049 VGND VGND VPWR VPWR net7048 sky130_fd_sc_hd__clkbuf_1
Xwire6303 net6304 VGND VGND VPWR VPWR net6303 sky130_fd_sc_hd__buf_1
Xwire6314 net6313 VGND VGND VPWR VPWR net6314 sky130_fd_sc_hd__buf_1
XFILLER_0_117_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6325 net6326 VGND VGND VPWR VPWR net6325 sky130_fd_sc_hd__buf_1
X_24265_ net4554 net4853 VGND VGND VPWR VPWR _04125_ sky130_fd_sc_hd__nand2_1
Xwire6336 net6333 VGND VGND VPWR VPWR net6336 sky130_fd_sc_hd__buf_1
Xfanout4806 net4814 VGND VGND VPWR VPWR net4806 sky130_fd_sc_hd__clkbuf_1
Xwire5602 net5606 VGND VGND VPWR VPWR net5602 sky130_fd_sc_hd__buf_1
X_21477_ net5961 net5943 VGND VGND VPWR VPWR _01490_ sky130_fd_sc_hd__xor2_1
Xwire6347 net6348 VGND VGND VPWR VPWR net6347 sky130_fd_sc_hd__clkbuf_1
Xmax_length2045 _02544_ VGND VGND VPWR VPWR net2045 sky130_fd_sc_hd__buf_1
Xwire5613 net5611 VGND VGND VPWR VPWR net5613 sky130_fd_sc_hd__clkbuf_2
Xmax_length1300 net1301 VGND VGND VPWR VPWR net1300 sky130_fd_sc_hd__clkbuf_1
Xwire5624 net5620 VGND VGND VPWR VPWR net5624 sky130_fd_sc_hd__clkbuf_1
X_23216_ _03053_ _03056_ VGND VGND VPWR VPWR _03086_ sky130_fd_sc_hd__xnor2_1
Xwire6369 cordic0.slte0.opA\[13\] VGND VGND VPWR VPWR net6369 sky130_fd_sc_hd__clkbuf_2
Xwire5635 net5634 VGND VGND VPWR VPWR net5635 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_15_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20428_ cordic0.slte0.opA\[11\] _12222_ _12223_ _12221_ VGND VGND VPWR VPWR _00494_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_160_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire4901 net4902 VGND VGND VPWR VPWR net4901 sky130_fd_sc_hd__clkbuf_1
Xwire5646 net5647 VGND VGND VPWR VPWR net5646 sky130_fd_sc_hd__buf_1
X_24196_ net4603 net4803 VGND VGND VPWR VPWR _04057_ sky130_fd_sc_hd__nand2_1
Xwire4912 net4913 VGND VGND VPWR VPWR net4912 sky130_fd_sc_hd__buf_1
Xwire5657 net5650 VGND VGND VPWR VPWR net5657 sky130_fd_sc_hd__buf_1
Xmax_length1355 net1356 VGND VGND VPWR VPWR net1355 sky130_fd_sc_hd__buf_1
Xwire5668 pid_d.mult0.b\[15\] VGND VGND VPWR VPWR net5668 sky130_fd_sc_hd__clkbuf_1
Xwire4934 net4935 VGND VGND VPWR VPWR net4934 sky130_fd_sc_hd__buf_1
Xwire5679 net5680 VGND VGND VPWR VPWR net5679 sky130_fd_sc_hd__buf_1
Xmax_length1377 net1378 VGND VGND VPWR VPWR net1377 sky130_fd_sc_hd__buf_1
X_23147_ net5140 net4681 VGND VGND VPWR VPWR _03017_ sky130_fd_sc_hd__nand2_1
X_20359_ net949 _12159_ VGND VGND VPWR VPWR _12160_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4967 net4968 VGND VGND VPWR VPWR net4967 sky130_fd_sc_hd__buf_1
Xwire4978 net4979 VGND VGND VPWR VPWR net4978 sky130_fd_sc_hd__clkbuf_1
Xwire4989 net4990 VGND VGND VPWR VPWR net4989 sky130_fd_sc_hd__clkbuf_1
X_23078_ _02947_ _02875_ _02887_ VGND VGND VPWR VPWR _02948_ sky130_fd_sc_hd__a21oi_1
X_22029_ _02024_ _02035_ VGND VGND VPWR VPWR _02036_ sky130_fd_sc_hd__xnor2_1
X_14920_ net6630 matmul0.matmul_stage_inst.d\[6\] net7411 net6532 VGND VGND VPWR VPWR
+ _06994_ sky130_fd_sc_hd__a22o_1
Xhold40 pid_d.curr_error\[13\] VGND VGND VPWR VPWR net8993 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 pid_q.target\[4\] VGND VGND VPWR VPWR net9004 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 pid_q.curr_int\[15\] VGND VGND VPWR VPWR net9015 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 matmul0.matmul_stage_inst.d\[12\] VGND VGND VPWR VPWR net9026 sky130_fd_sc_hd__dlygate4sd3_1
X_14851_ matmul0.a\[14\] matmul0.matmul_stage_inst.e\[14\] net3607 VGND VGND VPWR
+ VPWR _06943_ sky130_fd_sc_hd__mux2_1
Xhold84 pid_d.curr_error\[1\] VGND VGND VPWR VPWR net9037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 net149 VGND VGND VPWR VPWR net9048 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ net1923 _06068_ _06069_ VGND VGND VPWR VPWR _06070_ sky130_fd_sc_hd__o21a_1
X_17570_ net4019 svm0.tC\[3\] svm0.tC\[2\] net4003 VGND VGND VPWR VPWR _09452_ sky130_fd_sc_hd__a22o_1
X_14782_ _06817_ net7148 _06904_ _06905_ net7457 VGND VGND VPWR VPWR _06906_ sky130_fd_sc_hd__o32a_1
XFILLER_0_39_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16521_ _08570_ _08580_ VGND VGND VPWR VPWR _08581_ sky130_fd_sc_hd__nor2_1
X_13733_ _05992_ _06001_ VGND VGND VPWR VPWR _06002_ sky130_fd_sc_hd__xnor2_1
X_25719_ clknet_leaf_11_clk _00592_ net8602 VGND VGND VPWR VPWR pid_d.mult0.a\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19240_ _11076_ _11072_ net6273 VGND VGND VPWR VPWR _11077_ sky130_fd_sc_hd__a21o_1
X_16452_ net2622 net2631 VGND VGND VPWR VPWR _08513_ sky130_fd_sc_hd__nor2_1
X_13664_ _05872_ net451 VGND VGND VPWR VPWR _05934_ sky130_fd_sc_hd__xor2_1
Xfanout8122 net6 VGND VGND VPWR VPWR net8122 sky130_fd_sc_hd__dlymetal6s2s_1
X_15403_ _07206_ _07476_ VGND VGND VPWR VPWR _07477_ sky130_fd_sc_hd__and2_1
X_12615_ net6664 net6673 net6678 VGND VGND VPWR VPWR _04888_ sky130_fd_sc_hd__and3b_1
X_19171_ net2112 net2111 net2110 net2109 VGND VGND VPWR VPWR _11008_ sky130_fd_sc_hd__o2bb2a_1
X_16383_ net1252 net1087 net1079 VGND VGND VPWR VPWR _08445_ sky130_fd_sc_hd__mux2_1
X_13595_ net577 _05845_ _05864_ VGND VGND VPWR VPWR _05865_ sky130_fd_sc_hd__a21oi_1
Xfanout7443 net7450 VGND VGND VPWR VPWR net7443 sky130_fd_sc_hd__buf_1
Xwire8250 net8251 VGND VGND VPWR VPWR net8250 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18122_ net7089 net3263 _09694_ VGND VGND VPWR VPWR _09973_ sky130_fd_sc_hd__a21o_1
X_15334_ net1280 _07406_ _07407_ VGND VGND VPWR VPWR _07408_ sky130_fd_sc_hd__a21o_1
Xwire8261 net26 VGND VGND VPWR VPWR net8261 sky130_fd_sc_hd__clkbuf_1
Xwire8272 net8273 VGND VGND VPWR VPWR net8272 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire8283 net8284 VGND VGND VPWR VPWR net8283 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire8294 net21 VGND VGND VPWR VPWR net8294 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire7560 matmul0.b_in\[13\] VGND VGND VPWR VPWR net7560 sky130_fd_sc_hd__clkbuf_1
X_18053_ net7097 net3976 _09902_ VGND VGND VPWR VPWR _09904_ sky130_fd_sc_hd__nor3_1
X_15265_ _07264_ _07338_ VGND VGND VPWR VPWR _07339_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_53_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7571 net7572 VGND VGND VPWR VPWR net7571 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7582 net7583 VGND VGND VPWR VPWR net7582 sky130_fd_sc_hd__clkbuf_1
Xwire7593 net7594 VGND VGND VPWR VPWR net7593 sky130_fd_sc_hd__clkbuf_1
X_17004_ net7080 _08964_ _08965_ _08963_ VGND VGND VPWR VPWR _00327_ sky130_fd_sc_hd__a22o_1
Xfanout6797 net6805 VGND VGND VPWR VPWR net6797 sky130_fd_sc_hd__buf_1
X_14216_ _06470_ _06474_ VGND VGND VPWR VPWR _06475_ sky130_fd_sc_hd__xnor2_1
Xwire6870 cordic0.vec\[1\]\[13\] VGND VGND VPWR VPWR net6870 sky130_fd_sc_hd__clkbuf_1
X_15196_ net3552 net2757 net2794 net2819 VGND VGND VPWR VPWR _07270_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14147_ _06406_ _06407_ VGND VGND VPWR VPWR _06408_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14078_ net7666 net1123 VGND VGND VPWR VPWR _06341_ sky130_fd_sc_hd__and2_1
X_18955_ net3910 _10791_ VGND VGND VPWR VPWR _10792_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_184_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13029_ _05159_ _05300_ _05301_ VGND VGND VPWR VPWR _05302_ sky130_fd_sc_hd__o21ai_2
X_17906_ _09746_ _09739_ VGND VGND VPWR VPWR _09757_ sky130_fd_sc_hd__nand2_1
X_18886_ _10699_ _10727_ VGND VGND VPWR VPWR _10728_ sky130_fd_sc_hd__xnor2_1
X_17837_ _09678_ _09687_ VGND VGND VPWR VPWR _09688_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_179_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17768_ net7123 net7104 VGND VGND VPWR VPWR _09619_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_16_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16719_ _08745_ VGND VGND VPWR VPWR _00262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19507_ _11343_ net2507 VGND VGND VPWR VPWR _11344_ sky130_fd_sc_hd__or2b_1
X_17699_ _09574_ VGND VGND VPWR VPWR _09575_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19438_ _10971_ _11274_ net6183 VGND VGND VPWR VPWR _11275_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19369_ net6176 net6308 net6257 VGND VGND VPWR VPWR _11206_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21400_ _01309_ _01412_ _01413_ VGND VGND VPWR VPWR _01414_ sky130_fd_sc_hd__o21a_1
XFILLER_0_84_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22380_ net2057 _02315_ VGND VGND VPWR VPWR _02383_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21331_ net5731 net5576 VGND VGND VPWR VPWR _01345_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24050_ _03788_ _03793_ _03912_ VGND VGND VPWR VPWR _03913_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21262_ _00850_ _00857_ VGND VGND VPWR VPWR _01277_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4208 net4209 VGND VGND VPWR VPWR net4208 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_64_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire4219 net4220 VGND VGND VPWR VPWR net4219 sky130_fd_sc_hd__dlymetal6s2s_1
X_23001_ net5016 net4685 VGND VGND VPWR VPWR _02871_ sky130_fd_sc_hd__nand2_2
XFILLER_0_163_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20213_ _12035_ cordic0.slte0.opB\[2\] net2937 VGND VGND VPWR VPWR _12036_ sky130_fd_sc_hd__mux2_1
X_21193_ net3839 _01194_ _01188_ VGND VGND VPWR VPWR _01209_ sky130_fd_sc_hd__a21o_1
Xwire3507 _07096_ VGND VGND VPWR VPWR net3507 sky130_fd_sc_hd__buf_1
Xwire3518 net3519 VGND VGND VPWR VPWR net3518 sky130_fd_sc_hd__buf_1
Xwire3529 _07062_ VGND VGND VPWR VPWR net3529 sky130_fd_sc_hd__buf_1
X_20144_ _11887_ _11969_ _11970_ VGND VGND VPWR VPWR _11971_ sky130_fd_sc_hd__a21oi_1
Xwire2806 net2807 VGND VGND VPWR VPWR net2806 sky130_fd_sc_hd__buf_1
Xwire2817 net2818 VGND VGND VPWR VPWR net2817 sky130_fd_sc_hd__clkbuf_1
Xwire2828 _07080_ VGND VGND VPWR VPWR net2828 sky130_fd_sc_hd__buf_1
Xwire2839 _07040_ VGND VGND VPWR VPWR net2839 sky130_fd_sc_hd__buf_1
X_24952_ pid_q.ki\[13\] _04728_ net1637 VGND VGND VPWR VPWR _04729_ sky130_fd_sc_hd__mux2_1
X_20075_ _11897_ _11903_ VGND VGND VPWR VPWR _11904_ sky130_fd_sc_hd__xnor2_2
X_23903_ net7504 _03766_ _03767_ VGND VGND VPWR VPWR _03768_ sky130_fd_sc_hd__and3_1
X_24883_ net4479 net2397 net3699 net4476 VGND VGND VPWR VPWR _04680_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23834_ net5149 net3749 net3743 VGND VGND VPWR VPWR _03699_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_196_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_196_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23765_ _03532_ _03534_ _03630_ VGND VGND VPWR VPWR _03631_ sky130_fd_sc_hd__o21ai_1
X_20977_ _00983_ _00986_ _00992_ VGND VGND VPWR VPWR _00993_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_131_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6823 net6824 VGND VGND VPWR VPWR net6823 sky130_fd_sc_hd__clkbuf_1
X_25504_ clknet_leaf_39_clk _00384_ net8770 VGND VGND VPWR VPWR svm0.delta\[9\] sky130_fd_sc_hd__dfrtp_1
X_22716_ _02652_ VGND VGND VPWR VPWR _00598_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23696_ net744 _03562_ VGND VGND VPWR VPWR _03563_ sky130_fd_sc_hd__xor2_1
Xmax_length6867 net6868 VGND VGND VPWR VPWR net6867 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_length6889 net6887 VGND VGND VPWR VPWR net6889 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25435_ clknet_leaf_96_clk _00318_ net8445 VGND VGND VPWR VPWR matmul0.sin\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22647_ net805 net3077 net1697 _02608_ net8892 VGND VGND VPWR VPWR _00573_ sky130_fd_sc_hd__o311a_1
XFILLER_0_165_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13380_ _05554_ net1132 VGND VGND VPWR VPWR _05653_ sky130_fd_sc_hd__nand2_1
X_25366_ clknet_leaf_81_clk _00249_ net8495 VGND VGND VPWR VPWR matmul0.alpha_pass\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_22578_ net7317 _02554_ VGND VGND VPWR VPWR _02558_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire6111 net6109 VGND VGND VPWR VPWR net6111 sky130_fd_sc_hd__buf_1
X_24317_ _04105_ _04106_ _04168_ VGND VGND VPWR VPWR _04177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire6133 net6132 VGND VGND VPWR VPWR net6133 sky130_fd_sc_hd__buf_1
X_21529_ pid_d.prev_int\[3\] _01436_ _01437_ net5982 VGND VGND VPWR VPWR _01541_ sky130_fd_sc_hd__a31o_1
X_25297_ clknet_leaf_92_clk _00180_ net8429 VGND VGND VPWR VPWR matmul0.matmul_stage_inst.d\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire6144 net6145 VGND VGND VPWR VPWR net6144 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire6155 net6153 VGND VGND VPWR VPWR net6155 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire5421 net5422 VGND VGND VPWR VPWR net5421 sky130_fd_sc_hd__clkbuf_1
Xwire6166 net6168 VGND VGND VPWR VPWR net6166 sky130_fd_sc_hd__buf_1
X_15050_ _07075_ net1285 _07123_ VGND VGND VPWR VPWR _07124_ sky130_fd_sc_hd__a21o_1
XFILLER_0_50_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24248_ pid_q.curr_error\[8\] VGND VGND VPWR VPWR _04109_ sky130_fd_sc_hd__inv_2
Xwire5443 net5436 VGND VGND VPWR VPWR net5443 sky130_fd_sc_hd__buf_1
XFILLER_0_50_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14001_ _06165_ _06209_ VGND VGND VPWR VPWR _06266_ sky130_fd_sc_hd__nor2_1
Xwire6199 net6194 VGND VGND VPWR VPWR net6199 sky130_fd_sc_hd__buf_1
Xwire5454 net5455 VGND VGND VPWR VPWR net5454 sky130_fd_sc_hd__buf_1
Xwire4720 net4715 VGND VGND VPWR VPWR net4720 sky130_fd_sc_hd__clkbuf_1
Xwire5465 net5466 VGND VGND VPWR VPWR net5465 sky130_fd_sc_hd__buf_1
Xwire4731 net4732 VGND VGND VPWR VPWR net4731 sky130_fd_sc_hd__clkbuf_1
X_24179_ _04037_ _03957_ _04039_ VGND VGND VPWR VPWR _04040_ sky130_fd_sc_hd__a21o_1
Xwire5476 net5477 VGND VGND VPWR VPWR net5476 sky130_fd_sc_hd__buf_1
Xwire4742 net4743 VGND VGND VPWR VPWR net4742 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire5498 net5499 VGND VGND VPWR VPWR net5498 sky130_fd_sc_hd__buf_1
Xwire4764 net4765 VGND VGND VPWR VPWR net4764 sky130_fd_sc_hd__clkbuf_1
Xwire4775 net4777 VGND VGND VPWR VPWR net4775 sky130_fd_sc_hd__buf_1
Xwire4786 net4779 VGND VGND VPWR VPWR net4786 sky130_fd_sc_hd__clkbuf_1
Xwire4797 pid_q.mult0.b\[15\] VGND VGND VPWR VPWR net4797 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18740_ _10581_ _10584_ VGND VGND VPWR VPWR _10585_ sky130_fd_sc_hd__xor2_1
X_15952_ net2652 net2748 VGND VGND VPWR VPWR _08020_ sky130_fd_sc_hd__nor2_1
Xinput130 pid_q_data[0] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_1
Xinput141 pid_q_data[5] VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_1
X_14903_ net6612 net7420 matmul0.matmul_stage_inst.a\[10\] net6583 VGND VGND VPWR
+ VPWR _06977_ sky130_fd_sc_hd__a22o_1
X_18671_ net3923 _10516_ VGND VGND VPWR VPWR _10517_ sky130_fd_sc_hd__nor2_1
X_15883_ net2810 _07601_ net3397 net2737 VGND VGND VPWR VPWR _07952_ sky130_fd_sc_hd__a2bb2o_1
X_17622_ _09494_ _09499_ _09501_ _09502_ VGND VGND VPWR VPWR _09503_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_37_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14834_ matmul0.a\[6\] matmul0.matmul_stage_inst.e\[6\] net3611 VGND VGND VPWR VPWR
+ _06934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_187_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17553_ svm0.tC\[5\] VGND VGND VPWR VPWR _09435_ sky130_fd_sc_hd__inv_2
XFILLER_0_188_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14765_ net9034 net2858 net2865 _06893_ VGND VGND VPWR VPWR _00160_ sky130_fd_sc_hd__a22o_1
X_16504_ net2245 net2204 _08456_ net1244 VGND VGND VPWR VPWR _08564_ sky130_fd_sc_hd__o31a_1
X_13716_ _05888_ _05892_ _05893_ VGND VGND VPWR VPWR _05985_ sky130_fd_sc_hd__o21a_1
X_17484_ net6717 net2576 VGND VGND VPWR VPWR _09375_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14696_ net7153 _06839_ VGND VGND VPWR VPWR _06842_ sky130_fd_sc_hd__or2_2
X_19223_ _11048_ _11058_ _11059_ VGND VGND VPWR VPWR _11060_ sky130_fd_sc_hd__o21a_1
X_16435_ _08428_ _08480_ _08493_ _08483_ _08495_ VGND VGND VPWR VPWR _08496_ sky130_fd_sc_hd__o221a_1
X_13647_ _05914_ _05915_ VGND VGND VPWR VPWR _05917_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19154_ net6295 net3909 VGND VGND VPWR VPWR _10991_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16366_ _08427_ _08428_ VGND VGND VPWR VPWR _08429_ sky130_fd_sc_hd__nand2_1
X_13578_ _05783_ _05848_ VGND VGND VPWR VPWR _05849_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire8080 net8081 VGND VGND VPWR VPWR net8080 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18105_ net3949 _09877_ VGND VGND VPWR VPWR _09956_ sky130_fd_sc_hd__nor2_1
Xwire8091 net99 VGND VGND VPWR VPWR net8091 sky130_fd_sc_hd__clkbuf_1
X_15317_ _07389_ _07390_ VGND VGND VPWR VPWR _07391_ sky130_fd_sc_hd__xnor2_1
X_19085_ _10910_ net1757 VGND VGND VPWR VPWR _10922_ sky130_fd_sc_hd__nor2_1
X_16297_ net491 _08299_ VGND VGND VPWR VPWR _08361_ sky130_fd_sc_hd__nor2_1
Xfanout6572 net6579 VGND VGND VPWR VPWR net6572 sky130_fd_sc_hd__buf_1
XFILLER_0_152_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18036_ net7131 _09886_ VGND VGND VPWR VPWR _09887_ sky130_fd_sc_hd__and2_1
X_15248_ _07319_ net2704 _07321_ VGND VGND VPWR VPWR _07322_ sky130_fd_sc_hd__a21o_1
Xfanout5860 pid_d.mult0.b\[4\] VGND VGND VPWR VPWR net5860 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5882 net5885 VGND VGND VPWR VPWR net5882 sky130_fd_sc_hd__buf_1
XFILLER_0_10_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15179_ net1545 _07251_ _07252_ VGND VGND VPWR VPWR _07253_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_1_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19987_ _11816_ _11817_ VGND VGND VPWR VPWR _11818_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18938_ _10774_ _10776_ VGND VGND VPWR VPWR _10777_ sky130_fd_sc_hd__and2b_1
.ends

