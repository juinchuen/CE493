* NGSPICE file created from pid.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0683 ps=0.86 w=0.65 l=0.15
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X1 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X3 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_381_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VGND A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.0683 ps=0.86 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 VGND A1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_510_47# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X2 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X3 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X4 a_79_21# A2 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.162 ps=1.33 w=1 l=0.15
X5 a_297_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X6 a_79_21# C1 a_510_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.114 ps=1 w=0.65 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 a_215_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.106 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
X0 VGND A a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 Y a_38_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_38_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_820_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR a_38_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X5 VGND A a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND B a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND B a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y B a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_38_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_38_297# B a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VGND A a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_902_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_820_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_902_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 VPWR A a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 Y a_38_297# a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 Y a_38_297# a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 a_38_47# B a_38_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_38_47# B a_38_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 a_38_297# B a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X21 a_38_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 VPWR B a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X23 a_38_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X24 a_902_47# a_38_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 a_902_47# a_38_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 Y B a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_38_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 a_820_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VPWR A a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 VGND A a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 VPWR A a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 a_902_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X33 a_820_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 Y a_38_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X35 a_902_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X36 a_38_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 VPWR A a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X38 VPWR a_38_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X39 VPWR B a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
X0 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_806_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_806_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_806_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 X B a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 X a_112_47# a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_806_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND A a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 X B a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 VGND A a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_806_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.272 ps=2.56 w=1 l=0.15
X15 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X17 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X19 a_806_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR B a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 VPWR B a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X24 a_806_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 a_806_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X28 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 a_806_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.257 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X30 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 VPWR A a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 X a_112_47# a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X35 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 a_806_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X38 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X39 VPWR A a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
X0 X a_299_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X1 VPWR a_193_47# a_299_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 VGND a_193_47# a_299_93# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X6 X a_299_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
X0 a_219_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.157 ps=1.17 w=0.42 l=0.15
X1 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.157 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VPWR A a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 X a_219_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_301_297# a_27_53# a_219_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5 X a_219_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X6 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_219_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.167 ps=1.43 w=0.42 l=0.15
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.139 ps=1.08 w=0.42 l=0.15
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.12 ps=1.09 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.43 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.09 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X2 a_193_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 Y A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 a_109_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
X0 a_27_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_560_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2 VGND B a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0991 ps=0.955 w=0.65 l=0.15
X3 Y B a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y a_27_297# a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_474_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X7 VGND A a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_27_47# B a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_27_297# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VPWR B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X12 a_474_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_560_47# a_27_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14 VPWR A a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X15 Y a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X16 VPWR a_27_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X17 a_560_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 a_77_199# B2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.06 as=0.127 ps=1.04 w=0.65 l=0.15
X1 a_323_297# A2 a_227_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X2 a_227_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_227_47# B1 a_77_199# VNB sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.133 ps=1.06 w=0.65 l=0.15
X4 VGND a_77_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VPWR B1 a_539_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.205 ps=1.41 w=1 l=0.15
X6 a_227_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X7 VPWR a_77_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X8 a_77_199# A3 a_323_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X9 VGND A2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.107 ps=0.98 w=0.65 l=0.15
X10 a_227_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_539_297# B2 a_77_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.195 ps=1.39 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
X0 a_222_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X1 VPWR A1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X2 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_222_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.186 ps=1.41 w=0.42 l=0.15
X4 VGND A2 a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X5 a_448_47# a_222_93# a_79_199# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_79_199# a_222_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X7 a_544_297# A2 a_79_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8 a_448_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.41 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X17 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X18 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X19 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
X0 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_470_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_470_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_470_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.106 ps=0.975 w=0.65 l=0.15
X6 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X8 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X10 a_470_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.162 ps=1.33 w=1 l=0.15
X11 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 VPWR B a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X13 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VGND A a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X16 X a_112_47# a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 a_470_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X18 X B a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14 ps=1.28 w=1 l=0.15
X1 VGND A3 a_383_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X2 a_309_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0715 pd=0.87 as=0.153 ps=1.12 w=0.65 l=0.15
X3 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.153 pd=1.12 as=0.0747 ps=0.88 w=0.65 l=0.15
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X5 a_383_47# A2 a_309_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0715 ps=0.87 w=0.65 l=0.15
X6 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X7 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
X0 a_121_297# B a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_39_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=1 w=0.65 l=0.15
X2 VPWR a_39_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_39_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.156 ps=1.36 w=1 l=0.15
X4 VGND a_39_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.156 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VGND A a_39_297# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=1 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_39_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 a_223_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 Y A1 a_658_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR B1_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X3 a_223_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.145 ps=1.29 w=1 l=0.15
X4 Y a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 VGND A2 a_658_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_223_297# a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X7 Y a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.123 ps=1.03 w=0.65 l=0.15
X8 VPWR A2 a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 a_658_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.201 ps=1.27 w=0.65 l=0.15
X10 VPWR A1 a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_223_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 a_658_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X13 Y a_27_47# a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X14 a_223_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X15 VPWR A2 a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.155 ps=1.31 w=1 l=0.15
X16 VPWR A1 a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X17 a_658_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X18 VGND B1_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.27 ps=2.13 w=0.65 l=0.15
X19 a_223_297# a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X20 a_658_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X21 VGND A2 a_658_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X22 VGND a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.27 as=0.091 ps=0.93 w=0.65 l=0.15
X23 VGND a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X24 Y A1 a_658_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X25 Y a_27_47# a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
X0 VPWR A1 a_485_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_485_297# a_297_93# a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 a_297_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.108 ps=1.01 w=0.42 l=0.15
X3 a_581_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.01 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_79_21# a_297_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6 VGND A2 a_581_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.51 as=0.14 ps=1.28 w=1 l=0.15
X8 a_297_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.182 ps=1.51 w=0.42 l=0.15
X9 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X10 a_485_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
X0 a_298_297# a_27_413# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1 a_215_297# a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.136 ps=1.1 w=0.65 l=0.15
X2 a_298_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.258 ps=1.45 w=0.65 l=0.15
X4 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6 a_382_47# A1 a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.136 pd=1.1 as=0.111 ps=1.37 w=0.42 l=0.15
X8 VPWR A1 a_298_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND A2 a_382_47# VNB sky130_fd_pr__nfet_01v8 ad=0.258 pd=1.45 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_47# C a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y A a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.107 ps=0.98 w=0.65 l=0.15
X5 a_277_47# B a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_206_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.146 ps=1.34 w=0.42 l=0.15
X1 a_206_369# A2_N a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X2 VGND B2 a_489_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_585_369# B2 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0672 ps=0.74 w=0.42 l=0.15
X4 a_489_47# a_206_369# a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_489_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VPWR A2_N a_206_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.209 pd=1.35 as=0.129 ps=1.18 w=0.42 l=0.15
X7 a_76_199# a_206_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.209 ps=1.35 w=0.42 l=0.15
X8 a_205_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0662 pd=0.735 as=0.0986 ps=0.98 w=0.42 l=0.15
X9 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X10 VPWR B1 a_585_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.0986 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X1 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.157 ps=1.32 w=1 l=0.15
X3 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.965 w=0.65 l=0.15
X6 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X8 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X9 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X10 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X13 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.117 ps=1.01 w=0.65 l=0.15
X1 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.41 pd=1.82 as=0.135 ps=1.27 w=1 l=0.15
X2 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.175 ps=1.35 w=1 l=0.15
X4 a_277_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_27_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.41 ps=1.82 w=1 l=0.15
X10 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.18 ps=1.36 w=1 l=0.15
X11 a_277_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X13 Y A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.0975 ps=0.95 w=0.65 l=0.15
X14 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.172 ps=1.83 w=0.65 l=0.15
X2 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X3 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X4 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X5 a_326_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.127 ps=1.04 w=0.65 l=0.15
X6 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.635 pd=3.27 as=0.195 ps=1.39 w=1 l=0.15
X7 Y C1 a_326_47# VNB sky130_fd_pr__nfet_01v8 ad=0.393 pd=2.51 as=0.0683 ps=0.86 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
X0 VGND A2 a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0683 ps=0.86 w=0.65 l=0.15
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A1 a_114_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X3 a_114_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.185 ps=1.87 w=0.65 l=0.15
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X8 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X10 a_285_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
X11 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR a_80_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1 X a_80_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 VGND a_80_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.111 pd=0.99 as=0.091 ps=0.93 w=0.65 l=0.15
X3 a_386_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X4 X a_80_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X5 a_80_199# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.162 pd=1.15 as=0.111 ps=0.99 w=0.65 l=0.15
X6 a_386_297# B1 a_80_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_458_47# A1 a_80_199# VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.162 ps=1.15 w=0.65 l=0.15
X8 VPWR A1 a_386_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X9 VGND A2 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.123 ps=1.03 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
X0 VPWR a_212_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_297_47# a_27_413# a_212_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_212_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.229 ps=1.75 w=1 l=0.15
X3 X a_212_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_212_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0767 ps=0.785 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VPWR B a_212_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.229 pd=1.75 as=0.0609 ps=0.71 w=0.42 l=0.15
X7 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND a_212_413# X VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
X0 VPWR a_29_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_29_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.151 ps=1.35 w=1 l=0.15
X2 VPWR A a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3 VGND a_29_311# X VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_184_53# B a_112_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 VPWR C a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.151 pd=1.35 as=0.0744 ps=0.815 w=0.42 l=0.15
X6 X a_29_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.13 ps=1.11 w=0.65 l=0.15
X7 a_112_53# A a_29_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_29_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 VGND C a_184_53# VNB sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.11 as=0.0536 ps=0.675 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
X0 VPWR A a_49_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VGND a_285_47# a_391_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.5
X2 X a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VGND A a_49_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VPWR a_285_47# a_391_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.5
X5 a_285_47# a_49_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X6 a_285_47# a_49_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X7 X a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.108 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122 ps=1.08 w=0.65 l=0.15
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.0536 ps=0.675 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 a_78_199# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2 a_493_297# A2 a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X3 VPWR a_78_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.373 pd=1.75 as=0.28 ps=2.56 w=1 l=0.15
X4 VGND A2 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X5 a_78_199# B2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.117 ps=1.24 w=1 l=0.15
X6 a_215_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_215_47# B2 a_78_199# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_292_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.117 pd=1.24 as=0.373 ps=1.75 w=1 l=0.15
X9 VGND a_78_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 VPWR a_1059_315# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X8 VGND a_1059_315# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X11 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X12 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X13 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X14 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X16 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X18 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X19 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X20 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X21 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X22 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X23 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X24 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X25 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 a_388_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.25 as=0.153 ps=1.3 w=1 l=0.15
X1 a_105_352# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_297_47# a_105_352# Y VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VPWR A1 a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.127 ps=1.25 w=1 l=0.15
X5 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X6 VPWR B1_N a_105_352# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X7 Y a_105_352# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.178 ps=1.4 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
X0 Q a_1062_300# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.142 ps=1.28 w=1 l=0.15
X1 a_1020_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0657 ps=0.725 w=0.36 l=0.15
X2 a_572_47# a_193_47# a_475_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X3 VPWR a_1062_300# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0913 ps=0.855 w=0.42 l=0.15
X4 a_634_183# a_475_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.149 ps=1.22 w=0.64 l=0.15
X5 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.109 ps=1.36 w=0.42 l=0.15
X7 a_475_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X8 VGND a_1062_300# a_1020_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.41 as=0.066 ps=0.745 w=0.42 l=0.15
X9 VPWR a_634_183# a_568_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 Q a_1062_300# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0926 ps=0.935 w=0.65 l=0.15
X11 a_568_413# a_27_47# a_475_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0662 ps=0.735 w=0.42 l=0.15
X12 a_634_183# a_475_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X13 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0913 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_891_413# a_27_47# a_634_183# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X16 Q a_1062_300# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.106 ps=0.975 w=0.65 l=0.15
X17 VGND a_891_413# a_1062_300# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X18 VPWR a_1062_300# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X19 VGND a_1062_300# Q VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 Q a_1062_300# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X22 VGND a_1062_300# Q VNB sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X24 VPWR a_891_413# a_1062_300# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.28 ps=2.56 w=1 l=0.15
X25 a_891_413# a_193_47# a_634_183# VNB sky130_fd_pr__nfet_01v8 ad=0.0657 pd=0.725 as=0.0989 ps=0.995 w=0.36 l=0.15
X26 a_475_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0672 ps=0.74 w=0.42 l=0.15
X27 VGND a_634_183# a_572_47# VNB sky130_fd_pr__nfet_01v8 ad=0.149 pd=1.22 as=0.0687 ps=0.76 w=0.42 l=0.15
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X29 VPWR a_1062_300# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
X0 X a_61_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.167 ps=1.39 w=1 l=0.15
X1 VPWR a_61_75# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X2 VPWR B a_61_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VGND B a_147_75# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 X a_61_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.112 ps=1.04 w=0.65 l=0.15
X5 VGND a_61_75# X VNB sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.127 ps=1.04 w=0.65 l=0.15
X6 a_61_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X7 a_147_75# A a_61_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 a_281_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1 a_281_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.26 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X7 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X9 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.127 ps=1.04 w=0.65 l=0.15
X10 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.198 ps=1.26 w=0.65 l=0.15
X11 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.127 ps=1.04 w=0.65 l=0.15
X12 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 Y A3 a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.195 ps=1.39 w=1 l=0.15
X15 a_27_297# A2 a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
X0 a_297_47# a_27_47# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.103 ps=1 w=0.65 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0.103 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X6 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X8 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.128 ps=1.03 w=0.42 l=0.15
X9 a_193_413# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X11 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X11 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X18 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
X0 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_475_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_762_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.31 ps=1.62 w=1 l=0.15
X5 a_475_47# B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.091 ps=0.93 w=0.65 l=0.15
X6 VGND A2 a_475_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X10 a_80_21# A2 a_762_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_80_21# B1 a_475_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X12 a_80_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15 ps=1.3 w=1 l=0.15
X13 a_475_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.117 ps=1.01 w=0.65 l=0.15
X14 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 VPWR A1 a_934_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X16 a_934_297# A2 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X17 VPWR B1 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=1.62 as=0.14 ps=1.28 w=1 l=0.15
X18 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND A1 a_475_47# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.117 ps=1.01 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
X0 Y a_251_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y a_251_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X5 VGND a_251_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 VPWR B_N a_251_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X8 VGND B_N a_251_21# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_27_297# a_251_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 a_79_21# A1 a_348_47# VNB sky130_fd_pr__nfet_01v8 ad=0.115 pd=1 as=0.133 ps=1.06 w=0.65 l=0.15
X1 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.26 as=0.091 ps=0.93 w=0.65 l=0.15
X3 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 a_79_21# C1 a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5 VPWR A2 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X6 a_299_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.195 ps=1.39 w=1 l=0.15
X7 a_585_297# B1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8 a_348_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.06 as=0.2 ps=1.26 w=0.65 l=0.15
X9 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.115 ps=1 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
X0 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
X0 a_28_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 a_462_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 Y B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_462_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_28_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 a_462_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X7 Y B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y A1 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X11 a_28_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.145 ps=1.29 w=1 l=0.15
X12 VPWR A2 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X14 VGND A2 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X15 a_28_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X16 VPWR A1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X17 a_28_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 VGND A2 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X19 VPWR A2 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.155 ps=1.31 w=1 l=0.15
X20 a_28_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X21 Y A1 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X22 a_462_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X23 VPWR A1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 Y A1 a_478_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.377 ps=1.75 w=1 l=0.15
X2 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.305 ps=1.61 w=1 l=0.15
X3 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.335 ps=1.67 w=1 l=0.15
X4 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.138 ps=1.27 w=1 l=0.15
X5 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.377 pd=1.75 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_478_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_478_47# A2 a_730_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VGND A3 a_730_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12 ps=1.02 w=0.65 l=0.15
X10 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_730_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.02 as=0.205 ps=1.93 w=0.65 l=0.15
X16 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.15 ps=1.3 w=1 l=0.15
X18 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X19 a_730_47# A2 a_478_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
X0 VPWR A a_94_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.198 pd=1.39 as=0.305 ps=2.61 w=1 l=0.15
X1 a_294_47# B a_185_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.128 ps=1.04 w=0.65 l=0.15
X2 a_185_47# A a_94_47# VNB sky130_fd_pr__nfet_01v8 ad=0.128 pd=1.04 as=0.198 ps=1.91 w=0.65 l=0.15
X3 VPWR a_94_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND C a_294_47# VNB sky130_fd_pr__nfet_01v8 ad=0.138 pd=1.08 as=0.0683 ps=0.86 w=0.65 l=0.15
X5 a_94_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.198 ps=1.39 w=1 l=0.15
X6 X a_94_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.177 ps=1.36 w=1 l=0.15
X7 X a_94_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 VPWR C a_94_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.177 pd=1.36 as=0.14 ps=1.28 w=1 l=0.15
X9 X a_94_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138 ps=1.08 w=0.65 l=0.15
X10 VGND a_94_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X11 VPWR a_94_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND a_94_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X13 X a_94_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VPWR a_277_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_277_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 X a_277_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X5 a_277_47# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X6 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND a_277_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND a_277_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_193_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_361_47# A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 X a_277_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VGND A3 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X15 X a_277_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X16 a_277_47# A1 a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 a_445_47# A2 a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VGND B1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_27_297# B1 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X21 VPWR a_277_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.5 pd=3 as=0.135 ps=1.27 w=1 l=0.15
X22 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X23 a_277_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 Y A1 a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.119 ps=1.01 w=0.65 l=0.15
X1 a_181_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.0683 ps=0.86 w=0.65 l=0.15
X2 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.106 ps=0.975 w=0.65 l=0.15
X3 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.162 ps=1.33 w=1 l=0.15
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.153 ps=1.3 w=1 l=0.15
X6 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_467_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_467_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A1 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_109_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND A2 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
X0 VGND C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_277_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_27_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X8 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_277_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 a_300_297# a_27_413# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=0.15
X3 Y a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.102 ps=0.99 w=0.65 l=0.15
X4 VPWR A1 a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 a_384_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.143 ps=1.09 w=0.65 l=0.15
X6 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.111 ps=1.37 w=0.42 l=0.15
X7 a_300_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
X0 VGND A2 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X1 Y B1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 VPWR A1 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15
X4 a_29_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y A2 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND A1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X7 a_112_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X8 a_112_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.14 ps=1.28 w=1 l=0.15
X9 a_29_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X11 a_29_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.127 ps=1.04 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 VPWR A1 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 a_806_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.101 ps=0.96 w=0.65 l=0.15
X3 a_110_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VPWR A1 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X10 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_47# B1 a_1314_47# VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=2.09 as=0.104 ps=0.97 w=0.65 l=0.15
X12 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X14 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X17 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.0943 ps=0.94 w=0.65 l=0.15
X19 Y C1 a_978_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 Y C1 a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X22 a_27_47# B1 a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X23 a_110_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 a_806_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.675 pd=3.35 as=0.135 ps=1.27 w=1 l=0.15
X26 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.091 ps=0.93 w=0.65 l=0.15
X27 a_978_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.091 ps=0.93 w=0.65 l=0.15
X28 a_1314_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X31 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
X0 VPWR A a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_218_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.156 ps=1.16 w=0.42 l=0.15
X2 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.156 pd=1.16 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_300_297# a_27_53# a_218_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4 X a_218_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X5 VPWR a_218_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X6 X a_218_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148 ps=1.34 w=1 l=0.15
X7 VGND a_218_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X9 VGND A a_218_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
X0 a_109_93# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 a_215_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VGND a_109_93# a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3 VGND A a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VPWR A a_369_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 a_369_297# B a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_215_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X7 a_297_297# a_109_93# a_215_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_109_93# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X9 X a_215_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.1 ps=0.985 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.91 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148 ps=1.34 w=1 l=0.15
X9 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VPWR A2 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 a_277_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2 a_79_21# B1 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3 a_277_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_361_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_277_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.127 ps=1.04 w=0.65 l=0.15
X9 a_79_21# A1 a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.107 ps=0.98 w=0.65 l=0.15
X10 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=1.67 w=1 l=0.15
X1 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0.194 pd=1.95 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VGND B a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 Y a_27_93# a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 a_229_47# a_27_93# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y a_27_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.147 ps=1.34 w=1 l=0.15
X6 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.165 ps=1.33 w=1 l=0.15
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X8 a_229_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
X0 VPWR D a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_223_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.5 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 a_515_93# a_223_47# a_429_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 a_223_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.134 pd=1.48 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X5 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X6 X a_343_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.46 w=1 l=0.15
X7 a_429_93# a_27_47# a_343_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.118 ps=1.4 w=0.42 l=0.15
X8 VGND D a_615_93# VNB sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.11 as=0.0777 ps=0.79 w=0.42 l=0.15
X9 a_343_93# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X10 a_343_93# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X11 a_615_93# C a_515_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X12 X a_343_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.82 as=0.126 ps=1.11 w=0.65 l=0.15
X13 VPWR a_223_47# a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 Y a_61_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.183 ps=1.24 w=0.65 l=0.15
X1 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_217_297# a_61_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_479_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X4 a_217_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X5 Y a_61_47# a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VPWR A1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_61_47# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=0.15
X8 VGND A2 a_637_47# VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND a_61_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 Y A1 a_479_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0683 ps=0.86 w=0.65 l=0.15
X11 VGND B1_N a_61_47# VNB sky130_fd_pr__nfet_01v8 ad=0.183 pd=1.24 as=0.126 ps=1.44 w=0.42 l=0.15
X12 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X13 a_637_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X1 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_215_297# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_392_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0452 pd=0.635 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 a_465_297# B a_392_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.064 pd=0.725 as=0.0452 ps=0.635 w=0.42 l=0.15
X6 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR A a_465_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.064 ps=0.725 w=0.42 l=0.15
X8 a_297_297# a_109_53# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.064 ps=0.725 w=0.42 l=0.15
X11 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 a_286_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2 a_286_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.185 ps=1.87 w=0.65 l=0.15
X3 Y A2 a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 VGND A1 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.185 ps=1.87 w=0.65 l=0.15
X6 VGND A2 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7 a_487_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 a_27_47# B1 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10 VPWR A1 a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X13 a_487_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X14 a_286_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X15 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_449_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_449_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X15 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
X0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X7 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X13 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X14 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X16 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X17 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X18 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X19 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X20 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X21 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X22 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X23 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.92 as=0.107 ps=0.98 w=0.65 l=0.15
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.213 ps=1.42 w=1 l=0.15
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.127 ps=1.04 w=0.65 l=0.15
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
X0 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X1 Y a_27_93# a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_206_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X3 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X5 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR A1 a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.16 ps=1.32 w=1 l=0.15
X1 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.4 ps=1.8 w=1 l=0.15
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0894 ps=0.925 w=0.65 l=0.15
X3 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_470_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=1.8 as=0.138 ps=1.27 w=1 l=0.15
X6 a_384_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X7 a_384_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.104 ps=0.97 w=0.65 l=0.15
X8 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_455_297# B1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X2 a_28_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 a_821_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4 a_28_297# C1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 a_455_297# C1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.091 ps=0.93 w=0.65 l=0.15
X7 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 VPWR A2 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.2 ps=1.4 w=1 l=0.15
X9 Y D1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X10 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X11 VGND D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X13 a_821_297# B1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X15 Y D1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.117 ps=1.01 w=0.65 l=0.15
X17 a_1205_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X18 a_28_297# C1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14 ps=1.28 w=1 l=0.15
X19 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.127 ps=1.04 w=0.65 l=0.15
X20 a_1205_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X21 a_821_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.14 ps=1.28 w=1 l=0.15
X22 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X23 Y A1 a_1205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X24 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X25 VPWR A1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.145 ps=1.29 w=1 l=0.15
X26 Y A1 a_1205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.182 ps=1.86 w=0.65 l=0.15
X27 a_1205_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.02 as=0.091 ps=0.93 w=0.65 l=0.15
X28 a_28_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X29 VGND A2 a_1205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X30 a_455_297# B1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 a_821_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2 pd=1.4 as=0.15 ps=1.3 w=1 l=0.15
X32 a_1205_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X33 VGND A2 a_1205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.122 ps=1.02 w=0.65 l=0.15
X34 VPWR A1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.14 ps=1.28 w=1 l=0.15
X35 a_821_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X36 VPWR A2 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X37 a_455_297# C1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X38 a_821_297# B1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X39 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 VGND a_415_21# a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_415_21# A2_N a_717_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_717_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 VGND A2_N a_415_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_193_47# a_415_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR a_193_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_193_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_193_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_415_21# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X11 a_415_21# A2_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 X a_193_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_27_297# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_193_47# B2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 VGND B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 VGND a_193_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 VGND A1_N a_415_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VGND a_193_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_109_47# B2 a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 a_193_47# a_415_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 VPWR a_193_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 a_27_297# a_415_21# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X23 X a_193_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR A1_N a_717_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X26 a_717_297# A2_N a_415_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_109_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
X0 a_408_47# B a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_408_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y a_27_47# a_408_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.176 pd=1.39 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VGND C a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6 a_218_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.12 ps=1.04 w=0.65 l=0.15
X7 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_218_47# B a_408_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.176 ps=1.39 w=1 l=0.15
X12 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.04 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 VGND A2 a_485_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 VPWR A1 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 a_37_297# B1 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_485_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_292_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X7 VPWR A2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8 a_485_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X11 a_37_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 Y A1 a_485_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X13 Y C1 a_37_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X14 a_292_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X15 a_292_297# B1 a_37_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_297# a_419_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND a_419_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VGND a_419_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 Y a_419_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X11 Y a_419_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VGND B_N a_419_21# VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.182 ps=1.86 w=0.65 l=0.15
X13 Y a_419_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VPWR B_N a_419_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.27 ps=2.54 w=1 l=0.15
X15 a_27_297# a_419_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 Y a_419_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 a_56_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR A2 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
X3 a_139_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.266 ps=2.12 w=0.65 l=0.15
X4 a_311_297# B1 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X5 Y C1 a_311_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X6 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X7 Y A1 a_139_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 a_465_47# A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VGND A4 a_561_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X2 VPWR A3 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3 a_297_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4 a_297_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X5 VPWR A1 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_381_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.184 ps=1.22 w=0.65 l=0.15
X7 a_297_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9 a_79_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.184 pd=1.22 as=0.161 ps=1.14 w=0.65 l=0.15
X10 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.161 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_561_47# A3 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
X0 Y C a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X6 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X10 a_281_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
X0 a_121_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X1 VPWR a_35_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2 X a_35_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_35_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.115 ps=1 w=0.65 l=0.15
X4 X a_35_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR a_35_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 X a_35_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.177 ps=1.36 w=1 l=0.15
X7 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.177 pd=1.36 as=0.105 ps=1.21 w=1 l=0.15
X9 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.115 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 VGND A2 a_660_47# VNB sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X1 VGND C1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X2 a_414_297# C1 a_334_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X3 VGND a_85_193# X VNB sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X4 a_334_297# D1 a_85_193# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X5 a_516_297# B1 a_414_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X6 a_516_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7 a_660_47# A1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X8 a_85_193# D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X9 VPWR A1 a_516_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X10 a_85_193# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X11 VPWR a_85_193# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
X0 VGND B1_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VGND A2 a_478_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.106 ps=0.975 w=0.65 l=0.15
X2 a_478_47# a_27_93# a_174_21# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_478_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X6 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X7 VPWR A1 a_574_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X8 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR B1_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X10 a_574_297# A2 a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X11 a_174_21# a_27_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.395 ps=1.79 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X11 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
X0 a_27_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_27_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y A a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y A a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_27_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_27_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 a_445_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12 a_445_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_445_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X17 a_445_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X23 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.26 ps=1.45 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.4 ps=1.8 w=1 l=0.15
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.205 pd=1.93 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=1.8 as=0.135 ps=1.27 w=1 l=0.15
X5 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_109_297# C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 Y B1 a_383_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_301_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_301_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND B2 a_383_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y A1 a_735_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_27_297# B2 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VPWR A1 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND A2 a_735_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_301_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.176 ps=1.84 w=0.65 l=0.15
X12 VPWR A2 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X13 a_383_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X14 a_383_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_735_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X16 a_27_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X17 a_301_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X18 a_735_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_27_297# B1 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 Y A1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.109 ps=0.985 w=0.65 l=0.15
X4 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_949_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X8 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y C1 a_949_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15 ps=1.3 w=1 l=0.15
X10 a_781_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_27_297# B1 a_781_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 Y A1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_781_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_1301_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.15 ps=1.3 w=1 l=0.15
X16 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 Y C1 a_781_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.14 ps=1.28 w=1 l=0.15
X18 a_109_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_109_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 a_109_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0878 ps=0.92 w=0.65 l=0.15
X24 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=0.985 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X27 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X28 a_27_297# B1 a_1301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X29 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0894 ps=0.925 w=0.65 l=0.15
X30 a_109_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X31 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
X0 a_176_21# a_27_47# a_626_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X1 a_626_297# B a_542_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X3 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_542_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X8 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X12 a_176_21# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X13 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 a_397_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR B1_N a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X2 Y A2 a_397_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 VGND A2 a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VGND A1 a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_28_297# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X6 Y a_28_297# a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VPWR a_28_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 a_397_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X9 a_229_47# a_28_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 Y a_28_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X11 a_229_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_229_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VPWR A1 a_397_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
X0 VPWR S a_591_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X1 a_591_369# A0 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.131 ps=1.05 w=0.64 l=0.15
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.41 as=0.135 ps=1.27 w=1 l=0.15
X3 a_79_21# A1 a_306_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.131 pd=1.05 as=0.229 ps=1.36 w=0.64 l=0.15
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND S a_578_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0578 ps=0.695 w=0.42 l=0.15
X6 a_306_369# a_257_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.229 pd=1.36 as=0.178 ps=1.41 w=0.64 l=0.15
X7 a_79_21# A0 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=0.173 pd=1.25 as=0.0683 ps=0.745 w=0.42 l=0.15
X8 a_288_47# a_257_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X9 a_257_199# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_578_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.173 ps=1.25 w=0.42 l=0.15
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 a_257_199# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.173 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 VPWR A3 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X2 a_352_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.115 pd=1 as=0.21 ps=1.29 w=0.65 l=0.15
X3 a_549_47# A1 a_21_199# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.08 as=0.107 ps=0.98 w=0.65 l=0.15
X4 X a_21_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_21_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.21 pd=1.29 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_665_47# A2 a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.14 ps=1.08 w=0.65 l=0.15
X7 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X8 a_299_297# B1 a_21_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_21_199# B2 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND A3 a_665_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VPWR a_21_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 X a_21_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_21_199# B1 a_352_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.115 ps=1 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_27_47# a_415_21# a_193_297# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VPWR A2_N a_415_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_415_21# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X3 a_415_21# A2_N a_717_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_193_297# a_415_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR a_193_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_193_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_109_297# B2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_193_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_717_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_717_47# A2_N a_415_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 X a_193_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_27_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 VGND a_193_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 VGND A1_N a_717_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VGND a_193_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 a_193_297# a_415_21# a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 VPWR a_193_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR a_415_21# a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X23 X a_193_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR A1_N a_415_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 a_109_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X26 a_415_21# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 VGND B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
X0 VPWR a_30_53# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.315 pd=2.63 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND a_30_53# X VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 X a_30_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148 ps=1.34 w=1 l=0.15
X3 a_112_297# C a_30_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4 X a_30_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X5 VGND A a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_30_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VGND C a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_184_297# B a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X9 VPWR A a_184_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
X0 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X1 a_471_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.42 pd=2.84 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_27_47# C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=1.67 w=1 l=0.15
X8 a_277_47# B a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X9 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.135 ps=1.27 w=1 l=0.15
X10 Y A a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_277_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X13 a_471_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0894 ps=0.925 w=0.65 l=0.15
X1 a_191_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X2 VPWR A a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.119 ps=1.01 w=0.65 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_297_297# B a_191_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X6 a_109_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
X0 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 a_27_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_27_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=1.77 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X9 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.385 ps=1.77 w=1 l=0.15
X14 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X21 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X24 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 a_445_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_445_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X28 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X31 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 a_471_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_471_47# B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_471_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A1 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X5 a_471_47# B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_471_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_1241_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X10 a_27_47# B2 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VPWR B1 a_553_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND A2 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_553_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X14 a_27_47# B2 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 VGND A2 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 VGND A1 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X19 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 a_1241_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VPWR B1 a_553_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR A1 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 Y B2 a_553_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 a_1241_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X26 a_553_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_471_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X28 Y A2 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 a_553_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 a_27_47# B1 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X31 VGND A1 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X32 Y B2 a_553_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 a_1241_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 a_27_47# B1 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X35 a_553_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 Y A2 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X38 a_471_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X39 a_471_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 a_316_297# C1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.172 ps=1.35 w=1 l=0.15
X1 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.03 as=0.481 ps=2.78 w=0.65 l=0.15
X2 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.02 as=0.125 ps=1.03 w=0.65 l=0.15
X3 a_420_297# B1 a_316_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=1.58 as=0.185 ps=1.37 w=1 l=0.15
X4 VPWR A1 a_420_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.29 ps=1.58 w=1 l=0.15
X5 VGND A2 a_568_47# VNB sky130_fd_pr__nfet_01v8 ad=0.192 pd=1.89 as=0.0845 ps=0.91 w=0.65 l=0.15
X6 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.192 pd=1.24 as=0.12 ps=1.02 w=0.65 l=0.15
X7 a_420_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.138 ps=1.27 w=1 l=0.15
X8 a_217_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.755 ps=3.51 w=1 l=0.15
X9 a_568_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0845 pd=0.91 as=0.192 ps=1.24 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X2 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.338 pd=1.67 as=0.135 ps=1.27 w=1 l=0.15
X5 a_1249_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_1249_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.252 pd=1.5 as=0.338 ps=1.67 w=1 l=0.15
X12 a_803_47# A2 a_1249_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X16 a_803_47# A2 a_1249_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X20 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X21 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 a_1249_47# A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.133 ps=1.06 w=0.65 l=0.15
X23 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 a_1249_47# A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.252 ps=1.5 w=1 l=0.15
X28 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.06 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X30 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X32 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X33 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X35 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 VGND A3 a_1249_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X37 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X38 VGND A3 a_1249_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X39 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 a_484_297# B2 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND B2 a_566_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_96_21# B1 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X8 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_484_297# B1 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_484_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND A2 a_918_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_96_21# B2 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 a_96_21# B1 a_566_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_484_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR A1 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_96_21# A1 a_918_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 VPWR A2 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X18 a_566_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X19 a_918_47# A1 a_96_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 a_566_47# B1 a_96_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 a_918_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X22 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X23 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.115 ps=1 w=0.65 l=0.15
X1 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.115 pd=1 as=0.0926 ps=0.935 w=0.65 l=0.15
X2 VPWR A1 a_307_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.105 ps=1.21 w=1 l=0.15
X3 a_307_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.233 ps=1.47 w=1 l=0.15
X4 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.233 pd=1.47 as=0.112 ps=1.23 w=1 l=0.15
X6 a_109_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.112 pd=1.23 as=0.26 ps=2.52 w=1 l=0.15
X7 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
X0 a_176_21# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 VGND D_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.5 as=0.135 ps=1.27 w=1 l=0.15
X5 a_555_297# C a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 a_176_21# a_27_53# a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.169 ps=1.5 w=1 l=0.15
X8 a_387_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.168 ps=1.5 w=0.42 l=0.15
X9 a_483_297# B a_387_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 VGND a_27_53# a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 VPWR D_N a_27_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.169 pd=1.5 as=0.109 ps=1.36 w=0.42 l=0.15
X13 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1 ps=0.985 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 Y a_33_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_225_47# a_33_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VPWR a_33_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_33_297# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.182 ps=1.86 w=0.65 l=0.15
X4 Y a_33_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A2 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 Y a_33_297# a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 Y a_33_297# a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VGND A2 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VGND A2 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 a_561_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X11 a_225_47# a_33_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VPWR A1 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_225_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_225_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 VPWR A1 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 a_561_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR B1_N a_33_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X20 a_561_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 Y A2 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X24 a_561_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 VPWR a_33_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 a_676_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.213 ps=1.42 w=1 l=0.15
X1 a_512_47# B1 a_409_47# VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.26 as=0.119 ps=1.01 w=0.65 l=0.15
X2 a_306_47# D1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.198 ps=1.91 w=0.65 l=0.15
X3 VGND A2 a_512_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.198 ps=1.26 w=0.65 l=0.15
X4 VPWR C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.218 ps=1.43 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.42 as=0.305 ps=1.61 w=1 l=0.15
X6 VPWR A1 a_676_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X7 a_512_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_409_47# C1 a_306_47# VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.119 ps=1.01 w=0.65 l=0.15
X9 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.382 pd=1.76 as=0.26 ps=2.52 w=1 l=0.15
X10 a_79_21# D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=1.43 as=0.382 ps=1.76 w=1 l=0.15
X11 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 a_1224_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VPWR A1 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.183 ps=1.37 w=1 l=0.15
X2 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_806_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.205 ps=1.28 w=0.65 l=0.15
X8 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.205 pd=1.28 as=0.14 ps=1.08 w=0.65 l=0.15
X10 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_806_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 Y A3 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 Y A3 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X19 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.119 ps=1.01 w=0.65 l=0.15
X22 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0926 ps=0.935 w=0.65 l=0.15
X24 a_806_297# A2 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X25 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.142 ps=1.28 w=1 l=0.15
X28 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.08 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 a_1224_297# A2 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 a_1224_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.135 ps=1.27 w=1 l=0.15
X32 a_806_297# A2 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 VPWR A1 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X35 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X36 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X37 a_1224_297# A2 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X38 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X39 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 Y A3 a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_449_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 Y A3 a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A1 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y B1 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_449_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.263 ps=2.57 w=1 l=0.15
X8 Y B1 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_31_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 a_27_297# A2 a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.261 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND A1 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 a_31_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14 a_31_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_31_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_449_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X20 VGND A2 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VGND A2 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 VGND A3 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0.223 pd=1.34 as=0.0878 ps=0.92 w=0.65 l=0.15
X24 a_31_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.223 ps=1.34 w=0.65 l=0.15
X25 a_27_297# A2 a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 VGND A3 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 a_31_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.127 ps=1.04 w=0.65 l=0.15
X28 a_449_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 a_31_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 a_31_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.198 ps=1.26 w=0.65 l=0.15
X1 Y A3 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.393 pd=1.78 as=0.135 ps=1.27 w=1 l=0.15
X2 a_193_297# A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.393 ps=1.78 w=1 l=0.15
X5 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.26 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 a_429_297# A2 a_345_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND A2 a_345_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.08 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.26 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_345_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.14 ps=1.08 w=0.65 l=0.15
X5 a_345_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.305 ps=1.61 w=1 l=0.15
X6 a_629_297# B2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR B1 a_629_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.19 ps=1.38 w=1 l=0.15
X8 a_79_21# B2 a_345_47# VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_345_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.123 ps=1.03 w=0.65 l=0.15
X10 a_79_21# A3 a_429_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_345_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.198 ps=1.26 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
X0 VPWR A a_304_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X1 a_304_297# B a_220_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND C a_32_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.123 ps=1.03 w=0.65 l=0.15
X3 a_220_297# C a_114_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X4 a_32_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_32_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND A a_32_297# VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.123 ps=1.03 w=0.65 l=0.15
X11 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X13 a_114_297# D a_32_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
X14 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 a_33_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VGND A1 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VGND A2 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_33_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_797_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_797_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 Y B2 a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR B1 a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_33_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VGND A1 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 a_33_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_33_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_33_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_797_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.32 w=1 l=0.15
X17 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR B1 a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND A2 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 a_33_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 a_797_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.135 ps=1.27 w=1 l=0.15
X24 Y B2 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 Y B2 a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 Y B1 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.104 ps=0.97 w=0.65 l=0.15
X27 Y B2 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X28 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 Y B1 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 a_33_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
X0 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.177 pd=1.36 as=0.14 ps=1.28 w=1 l=0.15
X1 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138 ps=1.08 w=0.65 l=0.15
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND B a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.138 pd=1.08 as=0.0683 ps=0.86 w=0.65 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.177 ps=1.36 w=1 l=0.15
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.63 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.14 ps=1.28 w=1 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.305 ps=2.61 w=1 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.139 ps=1.5 w=0.42 l=0.15
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 a_79_21# C1 a_635_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.21 ps=1.42 w=1 l=0.15
X1 VPWR A2 a_319_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.17 ps=1.34 w=1 l=0.15
X2 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.08 as=0.133 ps=1.06 w=0.65 l=0.15
X3 a_417_47# A2 a_319_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.02 as=0.111 ps=0.99 w=0.65 l=0.15
X4 a_79_21# A1 a_417_47# VNB sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.06 as=0.12 ps=1.02 w=0.65 l=0.15
X5 a_319_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.111 pd=0.99 as=0.156 ps=1.13 w=0.65 l=0.15
X6 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.24 pd=1.48 as=0.135 ps=1.27 w=1 l=0.15
X7 a_319_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.185 ps=1.37 w=1 l=0.15
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.156 pd=1.13 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_319_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.34 as=0.24 ps=1.48 w=1 l=0.15
X10 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.14 ps=1.08 w=0.65 l=0.15
X11 a_635_297# B1 a_319_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.21 ps=1.42 w=1 l=0.15
X12 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
X0 VGND B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0926 ps=0.935 w=0.65 l=0.15
X1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.142 ps=1.28 w=1 l=0.15
X2 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VGND B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_215_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.254 pd=2.08 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=2.78 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X9 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_215_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X16 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X17 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
X0 Y a_53_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.192 ps=1.38 w=1 l=0.15
X1 a_232_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.192 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A_N a_53_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VGND A_N a_53_93# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_316_47# B a_232_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.03 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 Y a_53_93# a_316_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.125 ps=1.03 w=0.65 l=0.15
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
X0 Y a_74_47# a_265_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR B_N a_74_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.39 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_265_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.157 ps=1.39 w=1 l=0.15
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X4 VGND B_N a_74_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VGND a_74_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND a_215_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VPWR a_215_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_109_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X4 a_215_297# a_109_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.165 ps=1.82 w=0.65 l=0.15
X5 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.123 ps=1.03 w=0.65 l=0.15
X6 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X8 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_109_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10 VPWR A a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND a_215_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_487_297# B a_403_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_403_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X14 VPWR a_215_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.123 ps=1.03 w=0.65 l=0.15
X16 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 a_297_297# a_109_93# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 X a_91_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X1 a_91_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X2 a_360_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.137 ps=1.07 w=0.65 l=0.15
X3 VPWR B1 a_91_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.138 ps=1.27 w=1 l=0.15
X4 a_360_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.312 ps=1.62 w=1 l=0.15
X5 VGND A2 a_360_47# VNB sky130_fd_pr__nfet_01v8 ad=0.137 pd=1.07 as=0.114 ps=1 w=0.65 l=0.15
X6 a_360_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.203 ps=1.27 w=0.65 l=0.15
X7 VPWR a_91_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.62 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND a_91_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.203 pd=1.27 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 X a_91_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.208 ps=1.94 w=0.65 l=0.15
X10 a_677_47# B1 a_360_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.119 ps=1.01 w=0.65 l=0.15
X11 a_460_297# A2 a_360_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.175 ps=1.35 w=1 l=0.15
X12 a_91_21# C1 a_677_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X13 a_91_21# A3 a_460_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.21 ps=1.42 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 a_108_21# B1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.92 as=0.107 ps=0.98 w=0.65 l=0.15
X1 a_346_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X2 X a_108_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.263 ps=2.11 w=0.65 l=0.15
X3 a_108_21# A3 a_430_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X4 a_430_297# A2 a_346_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR a_108_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.175 ps=1.35 w=1 l=0.15
X6 a_346_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND A2 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 X a_108_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.405 ps=2.81 w=1 l=0.15
X9 VPWR B1 a_108_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.213 ps=1.42 w=1 l=0.15
X10 VGND a_108_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.114 ps=1 w=0.65 l=0.15
X11 a_346_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.127 ps=1.04 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 a_75_199# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.135 ps=1.07 w=0.65 l=0.15
X1 a_208_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.03 as=0.112 ps=0.995 w=0.65 l=0.15
X2 a_315_47# A2 a_208_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.125 ps=1.03 w=0.65 l=0.15
X3 VGND B1 a_75_199# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.07 as=0.106 ps=0.975 w=0.65 l=0.15
X4 a_75_199# A1 a_315_47# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.17 w=0.65 l=0.15
X5 a_75_199# C1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.207 ps=1.41 w=1 l=0.15
X6 a_544_297# B1 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.207 pd=1.41 as=0.162 ps=1.33 w=1 l=0.15
X7 VPWR a_75_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X8 a_201_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.142 ps=1.28 w=1 l=0.15
X9 VPWR A2 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.165 ps=1.33 w=1 l=0.15
X10 a_201_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.305 ps=1.61 w=1 l=0.15
X11 VGND a_75_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_475_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR A1 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X9 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.27 pd=1.48 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X12 a_475_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 Y A2 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X14 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.27 ps=1.48 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
X0 a_109_53# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_215_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.127 ps=1.1 w=0.65 l=0.15
X2 a_109_53# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X3 VGND C a_373_53# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.1 as=0.0536 ps=0.675 w=0.42 l=0.15
X4 VGND a_215_311# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR C a_215_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X6 VPWR a_215_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_215_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X8 a_301_53# a_109_53# a_215_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_215_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_373_53# B a_301_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 VPWR a_109_53# a_215_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand4bb_2 A_N B_N C D VGND VNB VPB VPWR Y
X0 VPWR a_193_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND D a_781_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y a_193_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X6 a_591_47# C a_781_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 a_781_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_781_47# C a_591_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR B_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10 a_193_47# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.197 pd=1.78 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 Y a_193_47# a_341_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 a_591_47# a_27_47# a_341_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14 a_341_47# a_193_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_341_47# a_27_47# a_591_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X17 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 a_193_47# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.197 pd=1.78 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 VGND B_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 a_27_47# C1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_47# C1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X4 a_1163_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0959 ps=0.945 w=0.65 l=0.15
X7 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 Y A2 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_1163_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.147 ps=1.29 w=1 l=0.15
X10 a_445_47# B1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_445_47# B1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR A1 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_27_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 VGND A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0959 ps=0.945 w=0.65 l=0.15
X18 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X20 a_1163_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 a_803_47# B1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.237 pd=1.48 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR A1 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 a_803_47# B1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 Y D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.237 ps=1.48 w=1 l=0.15
X28 a_445_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 a_803_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 a_1163_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X32 Y A2 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X33 a_445_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X34 a_803_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X35 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.0878 ps=0.92 w=0.65 l=0.15
X37 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X38 Y D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X39 VGND A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 a_30_297# C1 a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14 ps=1.28 w=1 l=0.15
X1 VGND C1 a_44_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.091 ps=0.93 w=0.65 l=0.15
X2 a_44_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.266 ps=1.47 w=0.65 l=0.15
X3 VGND a_44_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VPWR A1 a_477_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.257 ps=1.51 w=1 l=0.15
X5 VPWR a_44_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 X a_44_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7 VGND B1 a_44_47# VNB sky130_fd_pr__nfet_01v8 ad=0.266 pd=1.47 as=0.109 ps=0.985 w=0.65 l=0.15
X8 X a_44_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X9 a_477_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14 ps=1.28 w=1 l=0.15
X10 a_285_297# B1 a_477_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND D1 a_44_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X12 a_770_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.182 ps=1.86 w=0.65 l=0.15
X13 X a_44_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14 a_30_297# D1 a_44_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 VGND A2 a_770_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X16 a_44_47# D1 a_30_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X17 a_477_297# B1 a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.257 pd=1.51 as=0.14 ps=1.28 w=1 l=0.15
X18 a_770_47# A1 a_44_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0926 ps=0.935 w=0.65 l=0.15
X19 a_477_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X20 VPWR a_44_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X21 a_285_297# C1 a_30_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X22 a_44_47# D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X23 a_44_47# A1 a_770_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.091 ps=0.93 w=0.65 l=0.15
X24 VGND a_44_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X25 VPWR A2 a_477_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X26 X a_44_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 a_44_47# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=0.985 as=0.102 ps=0.965 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 VGND A1 a_474_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.104 ps=0.97 w=0.65 l=0.15
X1 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 VPWR A1 a_1122_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.252 pd=1.5 as=0.14 ps=1.28 w=1 l=0.15
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.192 pd=1.89 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VPWR C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.252 ps=1.5 w=1 l=0.15
X8 a_950_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X9 a_557_47# B1 a_474_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X10 a_474_47# B1 a_748_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X11 VGND A2 a_474_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_79_21# C1 a_557_47# VNB sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.1 as=0.0683 ps=0.86 w=0.65 l=0.15
X15 a_474_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X16 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.14 ps=1.28 w=1 l=0.15
X17 a_748_47# C1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.145 ps=1.1 w=0.65 l=0.15
X18 a_474_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.127 ps=1.04 w=0.65 l=0.15
X19 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.195 ps=1.39 w=1 l=0.15
X20 a_79_21# A2 a_950_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X21 a_1122_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X22 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.305 ps=1.61 w=1 l=0.15
X1 a_467_47# C1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VGND A2 a_717_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_467_47# B1 a_717_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VGND A1 a_717_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.135 ps=1.27 w=1 l=0.15
X6 a_79_21# C1 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_717_47# B1 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VGND A3 a_717_47# VNB sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.27 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_1147_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR A1 a_1147_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_1147_297# A2 a_875_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X18 a_79_21# A3 a_875_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X19 a_875_297# A3 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X20 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 a_875_297# A2 a_1147_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X22 a_717_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.201 ps=1.27 w=0.65 l=0.15
X23 a_717_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X24 a_717_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X26 VPWR C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X21 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 a_113_297# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_113_47# A2_N a_113_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VPWR B1 a_730_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A2_N a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_730_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_471_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_471_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 Y B2 a_730_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_113_297# A2_N a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_113_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X10 VGND A1_N a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VGND B2 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VPWR a_113_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X13 a_113_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X14 Y a_113_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.4 ps=1.8 w=1 l=0.15
X15 a_730_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.153 ps=1.3 w=1 l=0.15
X16 Y a_113_297# a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.176 ps=1.84 w=0.65 l=0.15
X17 a_471_47# a_113_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VPWR A1_N a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=1.8 as=0.135 ps=1.27 w=1 l=0.15
X19 VGND B1 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0991 ps=0.955 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X16 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X24 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
X0 VPWR a_315_380# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_315_380# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X2 a_315_380# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND C_N a_27_410# VNB sky130_fd_pr__nfet_01v8 ad=0.0619 pd=0.715 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VPWR C_N a_27_410# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.32 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VPWR A a_583_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_27_410# a_315_380# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.123 ps=1.03 w=0.65 l=0.15
X7 a_583_297# B a_499_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND A a_315_380# VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_397_297# a_205_93# a_315_380# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.258 ps=2.52 w=1 l=0.15
X10 X a_315_380# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.123 ps=1.03 w=0.65 l=0.15
X11 X a_315_380# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_499_297# a_27_410# a_397_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.18 ps=1.36 w=1 l=0.15
X13 VPWR a_315_380# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14 a_205_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0619 ps=0.715 w=0.42 l=0.15
X15 a_205_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.4 as=0.123 ps=1.32 w=0.42 l=0.15
X16 VGND a_315_380# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 VGND a_315_380# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 a_315_380# a_205_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.169 ps=1.82 w=0.65 l=0.15
X19 X a_315_380# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 a_240_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_51_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VGND A1 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_51_297# B2 a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.412 pd=1.83 as=0.105 ps=1.21 w=1 l=0.15
X4 a_149_47# C1 a_51_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.201 ps=1.92 w=0.65 l=0.15
X5 a_240_47# B1 a_149_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0991 ps=0.955 w=0.65 l=0.15
X6 VPWR A1 a_512_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X7 X a_51_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
X8 a_149_47# B2 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_245_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X10 VPWR C1 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X11 a_512_297# A2 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.412 ps=1.83 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_277_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.325 ps=1.65 w=1 l=0.15
X2 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_861_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.211 ps=1.3 w=0.65 l=0.15
X4 a_27_297# B1 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_1059_47# A2 a_861_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_1059_47# A1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_277_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X9 a_27_297# C1 a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.211 pd=1.3 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VGND A3 a_861_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VGND C1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VGND B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_109_47# A1 a_1059_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 a_109_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 VPWR A3 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X21 VPWR A2 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.325 pd=1.65 as=0.135 ps=1.27 w=1 l=0.15
X22 a_109_47# C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X23 VPWR A1 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X24 a_277_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 a_277_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X26 a_109_47# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X27 a_861_47# A2 a_1059_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
X0 VGND A a_311_413# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 VPWR A a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0598 ps=0.705 w=0.42 l=0.15
X2 a_393_413# a_205_93# a_311_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X3 VGND C_N a_27_410# VNB sky130_fd_pr__nfet_01v8 ad=0.0619 pd=0.715 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VPWR C_N a_27_410# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.32 as=0.109 ps=1.36 w=0.42 l=0.15
X5 X a_311_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X6 VGND a_27_410# a_311_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0598 ps=0.705 w=0.42 l=0.15
X7 a_561_297# B a_489_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0598 pd=0.705 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 a_205_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0619 ps=0.715 w=0.42 l=0.15
X9 a_205_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.123 ps=1.32 w=0.42 l=0.15
X10 a_489_297# a_27_410# a_393_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.122 ps=1.33 w=0.42 l=0.15
X11 a_311_413# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_311_413# a_205_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0598 pd=0.705 as=0.109 ps=1.36 w=0.42 l=0.15
X13 X a_311_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.102 ps=0.99 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
X0 a_174_21# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1 a_174_21# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.331 ps=1.71 w=0.42 l=0.15
X2 a_476_47# a_27_47# a_174_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X3 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.331 pd=1.71 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.141 ps=1.33 w=1 l=0.15
X5 a_548_47# a_505_280# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X7 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8 VPWR D a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 VGND D a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 VPWR a_505_280# a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X11 a_505_280# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X12 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_505_280# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X14 a_639_47# C a_548_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.064 ps=0.725 w=0.42 l=0.15
X15 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.14 ps=1.28 w=1 l=0.15
X1 a_235_47# C1 a_163_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.0683 ps=0.86 w=0.65 l=0.15
X2 a_343_47# B1 a_235_47# VNB sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.05 as=0.127 ps=1.04 w=0.65 l=0.15
X3 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.203 pd=1.4 as=0.195 ps=1.39 w=1 l=0.15
X4 a_454_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.203 ps=1.4 w=1 l=0.15
X5 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6 VPWR A1 a_454_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.195 ps=1.39 w=1 l=0.15
X7 a_163_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X8 VGND A2 a_343_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.132 ps=1.05 w=0.65 l=0.15
X9 a_343_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.127 ps=1.04 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
X0 a_388_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.148 ps=1.34 w=0.42 l=0.15
X1 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X7 a_176_21# a_27_47# a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_472_297# B a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
X10 a_176_21# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
X0 VGND B1 a_84_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_741_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.101 ps=0.96 w=0.65 l=0.15
X2 a_84_21# A1 a_741_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0747 ps=0.88 w=0.65 l=0.15
X3 VGND A2 a_901_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR A2 a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_483_297# B1 a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.185 ps=1.87 w=0.65 l=0.15
X8 a_84_21# B1 a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.265 pd=1.47 as=0.091 ps=0.93 w=0.65 l=0.15
X10 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_483_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=2.79 as=0.135 ps=1.27 w=1 l=0.15
X12 VPWR A1 a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X14 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X15 a_84_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.265 ps=1.47 w=0.65 l=0.15
X16 a_483_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X18 a_901_47# A1 a_84_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
X0 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.107 ps=0.98 w=0.65 l=0.15
X1 VGND D a_304_47# VNB sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.28 ps=1.62 w=1 l=0.15
X3 a_198_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0619 ps=0.715 w=0.42 l=0.15
X4 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X5 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X6 a_304_47# C a_198_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X7 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0746 pd=0.775 as=0.109 ps=1.36 w=0.42 l=0.15
X8 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.62 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.175 ps=1.26 w=0.65 l=0.15
X10 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0746 ps=0.775 w=0.42 l=0.15
X11 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0619 pd=0.715 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
X0 VGND a_91_199# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VPWR A a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X3 a_91_199# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_245_297# B a_161_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_91_199# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.146 ps=1.34 w=0.42 l=0.15
X7 a_161_297# a_91_199# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
X0 a_27_47# C a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_27_47# C a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_445_47# B a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_445_47# B a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 Y A a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X14 Y A a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_803_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X17 a_803_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_445_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 a_803_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X23 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X24 a_445_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 a_803_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X30 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X31 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X1 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X2 a_475_297# A2 a_729_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3 a_729_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR A1 a_729_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 a_729_297# A2 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_475_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y A3 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X15 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.228 pd=2 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X19 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 a_585_47# B1 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.119 ps=1.01 w=0.65 l=0.15
X1 VGND A2 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.137 pd=1.07 as=0.117 ps=1.01 w=0.65 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.62 as=0.26 ps=2.52 w=1 l=0.15
X3 a_81_21# C1 a_585_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.203 pd=1.27 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_266_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.312 ps=1.62 w=1 l=0.15
X6 a_368_297# A2 a_266_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.18 ps=1.36 w=1 l=0.15
X7 a_266_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.137 ps=1.07 w=0.65 l=0.15
X8 a_266_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.203 ps=1.27 w=0.65 l=0.15
X9 a_81_21# A3 a_368_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.21 ps=1.42 w=1 l=0.15
X10 a_81_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X11 VPWR B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.138 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
X0 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND a_531_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VPWR C_N a_531_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X9 a_281_297# a_531_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X10 Y a_531_21# a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X11 VGND C_N a_531_21# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X12 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X13 Y a_531_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 a_27_47# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.368 pd=1.74 as=0.14 ps=1.28 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.231 pd=2.01 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VPWR A1 a_373_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X4 a_182_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.165 ps=1.82 w=0.65 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.195 ps=1.39 w=1 l=0.15
X6 a_182_47# B1 a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X8 a_373_297# A2 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.368 ps=1.74 w=1 l=0.15
X9 a_110_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X10 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X11 VGND A1 a_182_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 VPWR A2_N a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.42 pd=1.84 as=0.135 ps=1.27 w=1 l=0.15
X1 Y a_112_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.42 ps=1.84 w=1 l=0.15
X2 VGND B2 a_394_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_112_297# A2_N a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.241 pd=2.04 as=0.0683 ps=0.86 w=0.65 l=0.15
X4 a_112_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.179 ps=1.85 w=0.65 l=0.15
X5 a_112_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X6 VPWR B1 a_478_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X7 a_394_47# a_112_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8 a_394_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_478_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand4bb_4 A_N B_N C D VGND VNB VPB VPWR Y
X0 Y a_27_47# a_432_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y a_27_47# a_432_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_850_47# a_193_47# a_432_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND D a_1266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.555 ps=2.11 w=1 l=0.15
X8 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X10 a_432_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_432_47# a_193_47# a_850_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_432_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_432_47# a_193_47# a_850_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR a_193_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.555 pd=2.11 as=0.135 ps=1.27 w=1 l=0.15
X16 a_193_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.495 pd=2.99 as=0.135 ps=1.27 w=1 l=0.15
X17 Y a_193_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 a_193_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.322 pd=2.29 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 a_850_47# C a_1266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.189 ps=1.88 w=0.65 l=0.15
X22 a_850_47# a_193_47# a_432_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 a_850_47# C a_1266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X24 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 VGND D a_1266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 VPWR a_193_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 a_1266_47# C a_850_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 Y a_193_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 a_1266_47# C a_850_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 a_1266_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X32 a_1266_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.0878 ps=0.92 w=0.65 l=0.15
X33 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X34 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X35 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
X0 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_467_297# A4 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VPWR A1 a_1243_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_27_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 Y A4 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_27_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VGND A4 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_1243_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 VGND A4 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR A1 a_1243_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 a_467_297# A4 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 a_1243_297# A2 a_885_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y A4 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X26 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X28 a_885_297# A2 a_1243_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 a_1243_297# A2 a_885_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 a_467_297# A3 a_885_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X33 a_885_297# A2 a_1243_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X34 a_885_297# A3 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X35 a_467_297# A3 a_885_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X37 a_1243_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X38 a_885_297# A3 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X39 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 a_27_47# B2 a_549_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VGND a_549_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VPWR a_549_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_297# A2 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 a_277_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_549_297# B2 a_739_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_739_297# B2 a_549_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X9 a_739_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_549_297# B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0975 ps=0.95 w=0.65 l=0.15
X13 a_277_297# A3 a_549_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR B1 a_739_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 X a_549_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_27_47# B1 a_549_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 a_549_297# A3 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X18 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X19 VPWR a_549_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND a_549_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 X a_549_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X23 a_549_297# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X24 X a_549_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X25 X a_549_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X27 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt pid VGND VPWR clock iterate_enable measurement[0] measurement[10] measurement[11]
+ measurement[12] measurement[13] measurement[14] measurement[15] measurement[16]
+ measurement[17] measurement[18] measurement[1] measurement[2] measurement[3] measurement[4]
+ measurement[5] measurement[6] measurement[7] measurement[8] measurement[9] out_clocked[0]
+ out_clocked[10] out_clocked[11] out_clocked[12] out_clocked[13] out_clocked[14]
+ out_clocked[15] out_clocked[16] out_clocked[17] out_clocked[18] out_clocked[1] out_clocked[2]
+ out_clocked[3] out_clocked[4] out_clocked[5] out_clocked[6] out_clocked[7] out_clocked[8]
+ out_clocked[9] reg_addr[0] reg_addr[10] reg_addr[11] reg_addr[12] reg_addr[13] reg_addr[14]
+ reg_addr[15] reg_addr[16] reg_addr[17] reg_addr[18] reg_addr[1] reg_addr[2] reg_addr[3]
+ reg_addr[4] reg_addr[5] reg_addr[6] reg_addr[7] reg_addr[8] reg_addr[9] reg_data[0]
+ reg_data[10] reg_data[11] reg_data[12] reg_data[13] reg_data[14] reg_data[15] reg_data[16]
+ reg_data[17] reg_data[18] reg_data[1] reg_data[2] reg_data[3] reg_data[4] reg_data[5]
+ reg_data[6] reg_data[7] reg_data[8] reg_data[9] reset target[0] target[10] target[11]
+ target[12] target[13] target[14] target[15] target[16] target[17] target[18] target[1]
+ target[2] target[3] target[4] target[5] target[6] target[7] target[8] target[9]
+ write_enable
X_09671_ net58 _03625_ _03658_ net298 VGND VGND VPWR VPWR _00056_ sky130_fd_sc_hd__a22o_1
X_18869_ _02153_ _09313_ VGND VGND VPWR VPWR _09314_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09938_ net344 _06007_ _06194_ net341 VGND VGND VPWR VPWR _06667_ sky130_fd_sc_hd__a22oi_1
X_09869_ _04577_ _05897_ _04566_ VGND VGND VPWR VPWR _05908_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11900_ _01837_ _01838_ VGND VGND VPWR VPWR _01839_ sky130_fd_sc_hd__nor2_1
X_12880_ net232 _01908_ _01873_ net236 VGND VGND VPWR VPWR _02819_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11831_ net242 net238 _01764_ _01769_ VGND VGND VPWR VPWR _01770_ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14550_ _04542_ _04562_ VGND VGND VPWR VPWR _04563_ sky130_fd_sc_hd__nor2_1
X_11762_ prev_error\[16\] VGND VGND VPWR VPWR _01701_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13501_ _03415_ _03410_ _03414_ VGND VGND VPWR VPWR _03460_ sky130_fd_sc_hd__o21ai_1
X_10713_ _00650_ _00651_ VGND VGND VPWR VPWR _00652_ sky130_fd_sc_hd__nor2_2
X_14481_ net448 net139 VGND VGND VPWR VPWR _04487_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11693_ _01614_ _01631_ _01629_ VGND VGND VPWR VPWR _01632_ sky130_fd_sc_hd__a21oi_1
X_16220_ _01706_ _06297_ VGND VGND VPWR VPWR _06400_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_125_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13432_ _03388_ _03389_ VGND VGND VPWR VPWR _03390_ sky130_fd_sc_hd__nand2_1
X_10644_ net361 _08196_ VGND VGND VPWR VPWR _00583_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16151_ _06323_ VGND VGND VPWR VPWR _06324_ sky130_fd_sc_hd__buf_2
X_13363_ _03312_ _03307_ _03310_ VGND VGND VPWR VPWR _03316_ sky130_fd_sc_hd__nor3_1
X_10575_ _00513_ _04291_ VGND VGND VPWR VPWR _00514_ sky130_fd_sc_hd__xor2_4
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer7 _08742_ VGND VGND VPWR VPWR net571 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_122_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15102_ _05169_ VGND VGND VPWR VPWR _05170_ sky130_fd_sc_hd__inv_2
X_12314_ _02030_ _02117_ VGND VGND VPWR VPWR _02253_ sky130_fd_sc_hd__and2_1
X_16082_ _06246_ _06247_ VGND VGND VPWR VPWR _06248_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13294_ _03233_ _03245_ VGND VGND VPWR VPWR _03247_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15033_ _05091_ _05002_ VGND VGND VPWR VPWR _05095_ sky130_fd_sc_hd__or2b_1
X_12245_ _02178_ _02183_ VGND VGND VPWR VPWR _02184_ sky130_fd_sc_hd__xor2_1
XFILLER_0_121_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12176_ _02114_ _02107_ VGND VGND VPWR VPWR _02115_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11127_ _01063_ _01064_ _00982_ _01065_ VGND VGND VPWR VPWR _01066_ sky130_fd_sc_hd__a2bb2o_1
X_16984_ _07167_ _07166_ VGND VGND VPWR VPWR _07241_ sky130_fd_sc_hd__and2b_1
XFILLER_0_155_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15935_ _05675_ _05942_ VGND VGND VPWR VPWR _06087_ sky130_fd_sc_hd__and2_1
X_18723_ _08785_ _08880_ VGND VGND VPWR VPWR _09154_ sky130_fd_sc_hd__nor2_1
X_11058_ _00992_ _00993_ _00995_ VGND VGND VPWR VPWR _00997_ sky130_fd_sc_hd__nor3_1
X_10009_ net356 net353 _05600_ VGND VGND VPWR VPWR _07448_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18654_ _08828_ VGND VGND VPWR VPWR _09078_ sky130_fd_sc_hd__inv_2
X_15866_ _03888_ _02354_ _03887_ VGND VGND VPWR VPWR _06011_ sky130_fd_sc_hd__nand3_1
XFILLER_0_149_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14817_ _04845_ _04847_ _04855_ VGND VGND VPWR VPWR _04857_ sky130_fd_sc_hd__nand3_1
XFILLER_0_87_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17605_ _07920_ _07922_ VGND VGND VPWR VPWR _07924_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_99_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18585_ _09001_ _08758_ _08882_ VGND VGND VPWR VPWR _09002_ sky130_fd_sc_hd__mux2_1
X_15797_ _05927_ _05933_ _05934_ _05891_ _05929_ VGND VGND VPWR VPWR _05935_ sky130_fd_sc_hd__o32a_1
XFILLER_0_98_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17536_ _07845_ _07847_ VGND VGND VPWR VPWR _07848_ sky130_fd_sc_hd__xnor2_1
X_14748_ _04779_ _04747_ _04777_ VGND VGND VPWR VPWR _04781_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_103_Left_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17467_ _07770_ _07771_ VGND VGND VPWR VPWR _07772_ sky130_fd_sc_hd__xnor2_2
X_14679_ _04701_ _04703_ _04704_ VGND VGND VPWR VPWR _04705_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_104_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19206_ clknet_4_12_0_clock _00088_ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dfxtp_1
X_16418_ net115 _06464_ VGND VGND VPWR VPWR _06618_ sky130_fd_sc_hd__xor2_4
XFILLER_0_13_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17398_ _07303_ _07304_ _07306_ _07307_ VGND VGND VPWR VPWR _07696_ sky130_fd_sc_hd__a22o_1
X_19137_ net503 net557 net494 _09561_ VGND VGND VPWR VPWR _00123_ sky130_fd_sc_hd__o211a_1
X_16349_ _06541_ VGND VGND VPWR VPWR _06542_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19068_ net505 net544 net496 VGND VGND VPWR VPWR _09518_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18019_ _08234_ _08378_ VGND VGND VPWR VPWR _08379_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_112_Left_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout116 net118 VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__buf_2
Xfanout127 kd_2\[16\] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__buf_2
Xfanout138 net140 VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__buf_2
Xfanout149 net150 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__dlymetal6s2s_1
X_09723_ net71 _04280_ VGND VGND VPWR VPWR _04302_ sky130_fd_sc_hd__nand2_1
X_09654_ net49 _03347_ _03380_ net199 VGND VGND VPWR VPWR _00009_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10360_ _00288_ _00298_ VGND VGND VPWR VPWR _00299_ sky130_fd_sc_hd__xor2_2
XFILLER_0_131_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10291_ _09596_ _00229_ VGND VGND VPWR VPWR _00230_ sky130_fd_sc_hd__or2_1
X_12030_ _01967_ _01968_ VGND VGND VPWR VPWR _01969_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13981_ _03937_ _03952_ VGND VGND VPWR VPWR _03953_ sky130_fd_sc_hd__xnor2_1
X_15720_ _05846_ _05849_ VGND VGND VPWR VPWR _05850_ sky130_fd_sc_hd__and2_1
X_12932_ _02775_ _02866_ _02870_ VGND VGND VPWR VPWR _02871_ sky130_fd_sc_hd__o21a_1
XFILLER_0_69_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15651_ _05773_ VGND VGND VPWR VPWR _05774_ sky130_fd_sc_hd__inv_2
X_12863_ net240 _01853_ _02801_ VGND VGND VPWR VPWR _02802_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14602_ _04614_ _04617_ _04619_ VGND VGND VPWR VPWR _04620_ sky130_fd_sc_hd__o21a_1
X_18370_ net529 _08755_ _08758_ _08762_ _08764_ VGND VGND VPWR VPWR _08765_ sky130_fd_sc_hd__a32oi_1
X_11814_ prev_error\[17\] _01699_ VGND VGND VPWR VPWR _01753_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15582_ _05687_ _05690_ _05686_ VGND VGND VPWR VPWR _05698_ sky130_fd_sc_hd__o21ba_1
X_12794_ _01847_ _02546_ _02659_ VGND VGND VPWR VPWR _02733_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_157_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17321_ _07221_ _07610_ VGND VGND VPWR VPWR _07611_ sky130_fd_sc_hd__xor2_4
X_14533_ _04539_ _04543_ VGND VGND VPWR VPWR _04545_ sky130_fd_sc_hd__and2_1
X_11745_ _00956_ _01683_ VGND VGND VPWR VPWR _01684_ sky130_fd_sc_hd__or2_2
XFILLER_0_56_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17252_ net316 _06351_ _07462_ VGND VGND VPWR VPWR _07535_ sky130_fd_sc_hd__and3_1
XFILLER_0_154_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14464_ _04373_ _04468_ VGND VGND VPWR VPWR _04469_ sky130_fd_sc_hd__nand2_1
X_11676_ net399 _00514_ VGND VGND VPWR VPWR _01615_ sky130_fd_sc_hd__nand2_1
X_16203_ _06378_ _06380_ VGND VGND VPWR VPWR _06382_ sky130_fd_sc_hd__xor2_1
XFILLER_0_52_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13415_ _03371_ _03279_ VGND VGND VPWR VPWR _03372_ sky130_fd_sc_hd__nor2_1
X_17183_ _07444_ _07458_ VGND VGND VPWR VPWR _07460_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10627_ net405 _05512_ _05523_ net387 _05171_ VGND VGND VPWR VPWR _00566_ sky130_fd_sc_hd__a32o_1
X_14395_ _03895_ _04389_ _04392_ VGND VGND VPWR VPWR _04393_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16134_ _06272_ _06305_ _01796_ VGND VGND VPWR VPWR _06306_ sky130_fd_sc_hd__a21boi_4
X_13346_ _03287_ _03298_ VGND VGND VPWR VPWR _03299_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10558_ _00481_ _00482_ _00496_ VGND VGND VPWR VPWR _00497_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16065_ _06200_ _06208_ _06210_ VGND VGND VPWR VPWR _06230_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_11_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13277_ _03216_ _03218_ _03229_ VGND VGND VPWR VPWR _03230_ sky130_fd_sc_hd__o21ba_1
X_10489_ _00423_ _00421_ VGND VGND VPWR VPWR _00428_ sky130_fd_sc_hd__and2b_1
X_15016_ _05069_ _05073_ VGND VGND VPWR VPWR _05076_ sky130_fd_sc_hd__nand2_1
X_12228_ _02165_ _02166_ VGND VGND VPWR VPWR _02167_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12159_ _02080_ _02082_ _02097_ VGND VGND VPWR VPWR _02098_ sky130_fd_sc_hd__a21oi_1
X_16967_ net329 _06314_ _06318_ _07221_ VGND VGND VPWR VPWR _07222_ sky130_fd_sc_hd__nand4_1
X_18706_ _09093_ _09105_ VGND VGND VPWR VPWR _09135_ sky130_fd_sc_hd__nand2_1
X_15918_ _03856_ _03423_ _03855_ VGND VGND VPWR VPWR _06068_ sky130_fd_sc_hd__and3_1
X_16898_ _07143_ _07144_ VGND VGND VPWR VPWR _07146_ sky130_fd_sc_hd__nand2_1
X_15849_ _05990_ _05991_ VGND VGND VPWR VPWR _05992_ sky130_fd_sc_hd__nor2_1
X_18637_ _06135_ _09052_ VGND VGND VPWR VPWR _09059_ sky130_fd_sc_hd__nor2_1
X_18568_ _08981_ _08982_ VGND VGND VPWR VPWR _08983_ sky130_fd_sc_hd__or2b_1
XFILLER_0_75_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17519_ net281 _02932_ _07661_ VGND VGND VPWR VPWR _07829_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_157_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18499_ _06266_ _08852_ VGND VGND VPWR VPWR _08907_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09706_ net504 VGND VGND VPWR VPWR _04115_ sky130_fd_sc_hd__inv_4
XFILLER_0_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09637_ net50 _03358_ _03391_ net266 VGND VGND VPWR VPWR _00010_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11530_ _01467_ _01468_ VGND VGND VPWR VPWR _01469_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_136_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_137_Right_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11461_ _01337_ _01340_ _01339_ VGND VGND VPWR VPWR _01400_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13200_ _03096_ _03152_ VGND VGND VPWR VPWR _03153_ sky130_fd_sc_hd__xnor2_1
X_10412_ _00315_ _00317_ _00344_ VGND VGND VPWR VPWR _00351_ sky130_fd_sc_hd__a21bo_1
X_14180_ _04153_ _04154_ _04155_ _04067_ VGND VGND VPWR VPWR _04156_ sky130_fd_sc_hd__a211o_1
X_11392_ _01317_ _01330_ VGND VGND VPWR VPWR _01331_ sky130_fd_sc_hd__and2b_1
X_13131_ _02973_ _02972_ _02945_ VGND VGND VPWR VPWR _03078_ sky130_fd_sc_hd__a21oi_1
X_10343_ _00190_ _00279_ _00280_ _00281_ VGND VGND VPWR VPWR _00282_ sky130_fd_sc_hd__o2bb2a_1
X_13062_ _02996_ _03000_ VGND VGND VPWR VPWR _03002_ sky130_fd_sc_hd__or2b_1
X_10274_ _00211_ _00206_ VGND VGND VPWR VPWR _00213_ sky130_fd_sc_hd__or2b_1
X_12013_ _01948_ _01951_ VGND VGND VPWR VPWR _01952_ sky130_fd_sc_hd__or2_1
X_17870_ _08117_ _08118_ _08132_ VGND VGND VPWR VPWR _08215_ sky130_fd_sc_hd__o21a_1
X_16821_ _07056_ _07057_ _07060_ VGND VGND VPWR VPWR _07061_ sky130_fd_sc_hd__o21ai_1
Xfanout480 net481 VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__buf_2
XFILLER_0_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout491 net497 VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__clkbuf_2
X_16752_ net271 _06891_ _06893_ VGND VGND VPWR VPWR _06985_ sky130_fd_sc_hd__a21oi_1
X_13964_ _03930_ _03935_ VGND VGND VPWR VPWR _03936_ sky130_fd_sc_hd__and2_1
X_15703_ net457 net195 VGND VGND VPWR VPWR _05832_ sky130_fd_sc_hd__nand2_1
X_12915_ _02845_ _02848_ VGND VGND VPWR VPWR _02854_ sky130_fd_sc_hd__or2_1
X_16683_ _06547_ _06552_ VGND VGND VPWR VPWR _06910_ sky130_fd_sc_hd__xnor2_1
X_13895_ _03178_ _03861_ VGND VGND VPWR VPWR _03862_ sky130_fd_sc_hd__nand2_1
X_15634_ _05744_ _05752_ _05755_ VGND VGND VPWR VPWR _05756_ sky130_fd_sc_hd__a21o_1
X_18422_ _08814_ _08820_ _08821_ VGND VGND VPWR VPWR _08822_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12846_ _02783_ _02784_ VGND VGND VPWR VPWR _02785_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18353_ _06133_ _08616_ VGND VGND VPWR VPWR _08747_ sky130_fd_sc_hd__nor2_1
X_15565_ net472 net474 net179 net176 VGND VGND VPWR VPWR _05680_ sky130_fd_sc_hd__and4_1
XFILLER_0_68_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12777_ _02712_ _02713_ _02715_ VGND VGND VPWR VPWR _02716_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17304_ net281 _07183_ _07592_ VGND VGND VPWR VPWR _07593_ sky130_fd_sc_hd__and3_1
X_14516_ _04524_ _04525_ VGND VGND VPWR VPWR _04526_ sky130_fd_sc_hd__nor2_1
X_11728_ _01401_ _01404_ _01402_ _01403_ VGND VGND VPWR VPWR _01667_ sky130_fd_sc_hd__o211a_1
X_18284_ _08668_ _08670_ VGND VGND VPWR VPWR _08671_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15496_ _05586_ _05603_ VGND VGND VPWR VPWR _05604_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17235_ _07464_ _07465_ _07477_ _07516_ VGND VGND VPWR VPWR _07517_ sky130_fd_sc_hd__a31o_1
X_14447_ net413 net417 net170 net165 VGND VGND VPWR VPWR _04450_ sky130_fd_sc_hd__and4_1
XFILLER_0_83_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_104_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11659_ net394 net390 _00814_ _00612_ VGND VGND VPWR VPWR _01598_ sky130_fd_sc_hd__and4_1
XFILLER_0_153_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17166_ _07434_ _07440_ VGND VGND VPWR VPWR _07441_ sky130_fd_sc_hd__xor2_1
X_14378_ _04282_ _04283_ _04285_ VGND VGND VPWR VPWR _04374_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16117_ prev_error\[7\] _09577_ _02328_ _06285_ _06286_ VGND VGND VPWR VPWR _06287_
+ sky130_fd_sc_hd__a221o_2
X_13329_ kd_1\[8\] _02410_ _03280_ _03281_ VGND VGND VPWR VPWR _03282_ sky130_fd_sc_hd__a31oi_2
X_17097_ _07353_ _07364_ VGND VGND VPWR VPWR _07365_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16048_ _06198_ _06199_ _06209_ VGND VGND VPWR VPWR _06211_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17999_ _08327_ _08356_ VGND VGND VPWR VPWR _08357_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10961_ _00821_ _00807_ VGND VGND VPWR VPWR _00900_ sky130_fd_sc_hd__or2b_1
X_12700_ _02638_ VGND VGND VPWR VPWR _02639_ sky130_fd_sc_hd__clkbuf_4
X_13680_ net247 _02641_ VGND VGND VPWR VPWR _03644_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10892_ _00742_ _00725_ _00741_ VGND VGND VPWR VPWR _00831_ sky130_fd_sc_hd__and3_1
X_12631_ _02568_ _02569_ VGND VGND VPWR VPWR _02570_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15350_ _05440_ _05441_ _05426_ _05433_ VGND VGND VPWR VPWR _05443_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_26_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12562_ _02495_ _02499_ _02500_ VGND VGND VPWR VPWR _02501_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14301_ _04256_ _04286_ _04288_ VGND VGND VPWR VPWR _04289_ sky130_fd_sc_hd__o21a_1
X_11513_ _01448_ _01451_ VGND VGND VPWR VPWR _01452_ sky130_fd_sc_hd__nor2_1
Xwire111 _01778_ VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__buf_4
X_15281_ _05301_ _05361_ VGND VGND VPWR VPWR _05367_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12493_ _02428_ _02431_ VGND VGND VPWR VPWR _02432_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17020_ net324 _06334_ VGND VGND VPWR VPWR _07280_ sky130_fd_sc_hd__nand2_1
X_14232_ _04153_ _04157_ _04212_ VGND VGND VPWR VPWR _04213_ sky130_fd_sc_hd__a21oi_2
X_11444_ _01373_ _01381_ _01382_ VGND VGND VPWR VPWR _01383_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14163_ _04076_ _03940_ _04128_ VGND VGND VPWR VPWR _04138_ sky130_fd_sc_hd__a21o_2
X_11375_ _01312_ _01313_ VGND VGND VPWR VPWR _01314_ sky130_fd_sc_hd__and2_1
X_13114_ _03056_ _03059_ VGND VGND VPWR VPWR _03060_ sky130_fd_sc_hd__nor2_1
X_10326_ _00263_ _00264_ VGND VGND VPWR VPWR _00265_ sky130_fd_sc_hd__and2b_2
X_18971_ _09306_ _09323_ _09321_ VGND VGND VPWR VPWR _09426_ sky130_fd_sc_hd__a21oi_1
X_14094_ _03950_ _04047_ _04064_ VGND VGND VPWR VPWR _04066_ sky130_fd_sc_hd__nand3_1
X_13045_ _02981_ _02975_ _02980_ VGND VGND VPWR VPWR _02984_ sky130_fd_sc_hd__and3_1
X_17922_ _08269_ _08271_ VGND VGND VPWR VPWR _08272_ sky130_fd_sc_hd__and2b_1
X_10257_ _05545_ _00195_ VGND VGND VPWR VPWR _00196_ sky130_fd_sc_hd__xnor2_1
X_10188_ _09274_ _09406_ VGND VGND VPWR VPWR _09417_ sky130_fd_sc_hd__or2b_1
X_17853_ net301 _02931_ _08195_ VGND VGND VPWR VPWR _08197_ sky130_fd_sc_hd__and3_1
X_16804_ _06936_ _07042_ VGND VGND VPWR VPWR _07043_ sky130_fd_sc_hd__nor2_1
X_14996_ _04925_ _05053_ VGND VGND VPWR VPWR _05054_ sky130_fd_sc_hd__or2_1
X_17784_ _08089_ _08096_ VGND VGND VPWR VPWR _08121_ sky130_fd_sc_hd__nand2_1
X_16735_ net284 _06621_ _06881_ VGND VGND VPWR VPWR _06967_ sky130_fd_sc_hd__a21oi_1
X_13947_ _03911_ _03917_ _03918_ VGND VGND VPWR VPWR _03919_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16666_ _06890_ VGND VGND VPWR VPWR _06891_ sky130_fd_sc_hd__clkbuf_4
X_13878_ _03719_ _03750_ _03843_ VGND VGND VPWR VPWR _03844_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15617_ _05719_ _05720_ VGND VGND VPWR VPWR _05737_ sky130_fd_sc_hd__xnor2_1
X_18405_ _08800_ _08803_ net571 VGND VGND VPWR VPWR _08804_ sky130_fd_sc_hd__or3_1
XFILLER_0_147_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12829_ _02678_ _02763_ _02767_ VGND VGND VPWR VPWR _02768_ sky130_fd_sc_hd__o21a_1
XFILLER_0_69_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16597_ _06813_ _06814_ VGND VGND VPWR VPWR _06815_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15548_ _05623_ _05630_ _05632_ VGND VGND VPWR VPWR _05661_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18336_ _08682_ net530 _08727_ VGND VGND VPWR VPWR _08728_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18267_ _08651_ VGND VGND VPWR VPWR _08652_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15479_ _05502_ _05584_ VGND VGND VPWR VPWR _05585_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17218_ _07488_ _07496_ _07497_ VGND VGND VPWR VPWR _07498_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18198_ _08574_ _08575_ i_error\[6\] VGND VGND VPWR VPWR _08576_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17149_ _07405_ _07421_ VGND VGND VPWR VPWR _07422_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_130_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09971_ net339 _05336_ VGND VGND VPWR VPWR _07030_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11160_ _01085_ _01097_ VGND VGND VPWR VPWR _01099_ sky130_fd_sc_hd__and2_1
X_10111_ net344 _04841_ _04852_ VGND VGND VPWR VPWR _08570_ sky130_fd_sc_hd__and3_2
X_11091_ _00819_ _01029_ _00912_ VGND VGND VPWR VPWR _01030_ sky130_fd_sc_hd__a21bo_1
X_10042_ _07778_ _07800_ _07349_ VGND VGND VPWR VPWR _07811_ sky130_fd_sc_hd__o21ai_1
Xhold41 i_error\[0\] VGND VGND VPWR VPWR net548 sky130_fd_sc_hd__dlygate4sd3_1
X_14850_ _04887_ _04891_ _04892_ VGND VGND VPWR VPWR _04893_ sky130_fd_sc_hd__a21oi_1
Xhold52 i_error\[5\] VGND VGND VPWR VPWR net559 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13801_ net247 _02934_ _03755_ VGND VGND VPWR VPWR _03767_ sky130_fd_sc_hd__a21o_1
X_14781_ _04803_ _04806_ _04815_ VGND VGND VPWR VPWR _04817_ sky130_fd_sc_hd__or3_1
X_11993_ _01789_ _01931_ _01772_ VGND VGND VPWR VPWR _01932_ sky130_fd_sc_hd__and3b_1
X_16520_ _06715_ _06717_ _06729_ VGND VGND VPWR VPWR _06730_ sky130_fd_sc_hd__a21bo_1
X_13732_ net243 net240 _02934_ _02914_ VGND VGND VPWR VPWR _03698_ sky130_fd_sc_hd__and4_1
XFILLER_0_86_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10944_ _00786_ _00788_ VGND VGND VPWR VPWR _00883_ sky130_fd_sc_hd__xor2_1
X_16451_ _06610_ _06608_ VGND VGND VPWR VPWR _06654_ sky130_fd_sc_hd__xor2_1
XFILLER_0_129_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13663_ _03566_ _03624_ VGND VGND VPWR VPWR _03626_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10875_ _00813_ VGND VGND VPWR VPWR _00814_ sky130_fd_sc_hd__buf_2
X_15402_ _05487_ _05476_ _05485_ VGND VGND VPWR VPWR _05500_ sky130_fd_sc_hd__nand3_1
X_12614_ _02550_ _02552_ VGND VGND VPWR VPWR _02553_ sky130_fd_sc_hd__nand2_1
X_19170_ net501 net454 VGND VGND VPWR VPWR _09581_ sky130_fd_sc_hd__or2_1
X_16382_ _06451_ _06485_ VGND VGND VPWR VPWR _06578_ sky130_fd_sc_hd__nand2_1
X_13594_ _03551_ _03552_ VGND VGND VPWR VPWR _03553_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18121_ _08484_ _08490_ VGND VGND VPWR VPWR _08491_ sky130_fd_sc_hd__xnor2_2
X_15333_ _05338_ _05423_ VGND VGND VPWR VPWR _05425_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12545_ net241 _01807_ VGND VGND VPWR VPWR _02484_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18052_ _08411_ _08412_ _08348_ _08373_ VGND VGND VPWR VPWR _08415_ sky130_fd_sc_hd__o22a_1
X_15264_ _05346_ _05348_ VGND VGND VPWR VPWR _05349_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12476_ _02401_ _02403_ VGND VGND VPWR VPWR _02415_ sky130_fd_sc_hd__xor2_1
XFILLER_0_41_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17003_ net282 _07157_ VGND VGND VPWR VPWR _07262_ sky130_fd_sc_hd__nand2_1
X_14215_ _04138_ _04194_ VGND VGND VPWR VPWR _04195_ sky130_fd_sc_hd__xor2_1
XFILLER_0_151_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11427_ net377 _00408_ _01365_ VGND VGND VPWR VPWR _01366_ sky130_fd_sc_hd__a21bo_1
XANTENNA_5 _06133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15195_ net427 net433 net193 net189 VGND VGND VPWR VPWR _05273_ sky130_fd_sc_hd__and4_1
XFILLER_0_105_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14146_ _04117_ _04105_ _04056_ VGND VGND VPWR VPWR _04119_ sky130_fd_sc_hd__nand3_1
XFILLER_0_1_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11358_ _01240_ _01236_ VGND VGND VPWR VPWR _01297_ sky130_fd_sc_hd__and2b_1
X_10309_ net342 _08207_ _00247_ VGND VGND VPWR VPWR _00248_ sky130_fd_sc_hd__and3_1
X_14077_ net412 net418 net140 net134 VGND VGND VPWR VPWR _04049_ sky130_fd_sc_hd__and4_1
X_18954_ _09227_ _09267_ _09407_ VGND VGND VPWR VPWR _09408_ sky130_fd_sc_hd__o21a_1
X_11289_ _01160_ _01162_ VGND VGND VPWR VPWR _01228_ sky130_fd_sc_hd__xnor2_1
X_13028_ _02947_ _02966_ VGND VGND VPWR VPWR _02967_ sky130_fd_sc_hd__or2_1
X_17905_ _08244_ _08252_ _08253_ VGND VGND VPWR VPWR _08254_ sky130_fd_sc_hd__nor3_1
X_18885_ _09330_ _09331_ VGND VGND VPWR VPWR _09332_ sky130_fd_sc_hd__or2_1
X_17836_ net318 _07093_ VGND VGND VPWR VPWR _08178_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer17 _08917_ VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__clkbuf_1
X_17767_ _08100_ _08080_ _08101_ VGND VGND VPWR VPWR _08102_ sky130_fd_sc_hd__a21bo_1
X_14979_ _05018_ _05033_ _05034_ VGND VGND VPWR VPWR _05035_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_77_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16718_ net306 _06352_ VGND VGND VPWR VPWR _06948_ sky130_fd_sc_hd__nand2_1
X_17698_ _08003_ _08005_ VGND VGND VPWR VPWR _08026_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16649_ _06857_ _06871_ VGND VGND VPWR VPWR _06872_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18319_ _06566_ _08660_ _06559_ VGND VGND VPWR VPWR _08709_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19299_ clknet_4_8_0_clock _00039_ VGND VGND VPWR VPWR ki\[10\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_127_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09954_ _06832_ VGND VGND VPWR VPWR _06843_ sky130_fd_sc_hd__inv_2
X_09885_ net344 net341 _06073_ _05325_ VGND VGND VPWR VPWR _06084_ sky130_fd_sc_hd__and4_1
XFILLER_0_148_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10660_ _00597_ _00598_ VGND VGND VPWR VPWR _00599_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_149_Left_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10591_ _00436_ _00448_ VGND VGND VPWR VPWR _00530_ sky130_fd_sc_hd__xnor2_1
X_12330_ _02264_ _02268_ VGND VGND VPWR VPWR _02269_ sky130_fd_sc_hd__xor2_1
XFILLER_0_32_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12261_ _02192_ _02195_ _02199_ VGND VGND VPWR VPWR _02200_ sky130_fd_sc_hd__a21oi_1
X_14000_ net425 net430 net137 net136 VGND VGND VPWR VPWR _03972_ sky130_fd_sc_hd__and4_1
XFILLER_0_120_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11212_ _01087_ _01095_ VGND VGND VPWR VPWR _01151_ sky130_fd_sc_hd__xor2_1
X_12192_ _02127_ _02130_ VGND VGND VPWR VPWR _02131_ sky130_fd_sc_hd__or2_1
X_11143_ _01066_ _01074_ _01073_ VGND VGND VPWR VPWR _01082_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_128_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput86 net86 VGND VGND VPWR VPWR out_clocked[15] sky130_fd_sc_hd__clkbuf_4
Xoutput97 net97 VGND VGND VPWR VPWR out_clocked[8] sky130_fd_sc_hd__buf_2
X_15951_ _06057_ _06059_ VGND VGND VPWR VPWR _06104_ sky130_fd_sc_hd__xnor2_1
X_11074_ _00991_ _01011_ _01012_ VGND VGND VPWR VPWR _01013_ sky130_fd_sc_hd__nor3_1
X_10025_ _07393_ _07404_ VGND VGND VPWR VPWR _07624_ sky130_fd_sc_hd__xor2_1
X_14902_ _04947_ _04949_ VGND VGND VPWR VPWR _04950_ sky130_fd_sc_hd__nor2_1
X_15882_ _06024_ _06027_ VGND VGND VPWR VPWR _06028_ sky130_fd_sc_hd__or2_1
X_18670_ _06096_ _09094_ VGND VGND VPWR VPWR _09095_ sky130_fd_sc_hd__and2_1
X_17621_ _07913_ _07914_ VGND VGND VPWR VPWR _07941_ sky130_fd_sc_hd__nand2_1
X_14833_ _04760_ _04762_ _04765_ VGND VGND VPWR VPWR _04875_ sky130_fd_sc_hd__or3_1
XFILLER_0_144_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14764_ _04795_ _04798_ VGND VGND VPWR VPWR _04799_ sky130_fd_sc_hd__or2_1
X_17552_ _07861_ _07863_ _07864_ VGND VGND VPWR VPWR _07865_ sky130_fd_sc_hd__or3_1
X_11976_ _01870_ _01904_ _01914_ VGND VGND VPWR VPWR _01915_ sky130_fd_sc_hd__o21bai_1
X_16503_ net289 net286 _06409_ _06402_ VGND VGND VPWR VPWR _06712_ sky130_fd_sc_hd__and4_1
X_13715_ net267 _02222_ _02639_ net251 VGND VGND VPWR VPWR _03681_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10927_ _00864_ _00865_ VGND VGND VPWR VPWR _00866_ sky130_fd_sc_hd__xnor2_4
X_17483_ net540 _07788_ net270 VGND VGND VPWR VPWR _07790_ sky130_fd_sc_hd__and3b_1
X_14695_ net439 net155 _04517_ VGND VGND VPWR VPWR _04723_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19222_ clknet_4_5_0_clock _00104_ VGND VGND VPWR VPWR prev_error\[9\] sky130_fd_sc_hd__dfxtp_4
X_16434_ _06628_ _06632_ _06635_ VGND VGND VPWR VPWR _06636_ sky130_fd_sc_hd__a21oi_1
X_13646_ _03573_ _03606_ _03602_ VGND VGND VPWR VPWR _03607_ sky130_fd_sc_hd__a21o_1
X_10858_ _00713_ _00715_ VGND VGND VPWR VPWR _00797_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19153_ net505 net554 net495 _09570_ VGND VGND VPWR VPWR _00131_ sky130_fd_sc_hd__o211a_1
X_16365_ _06500_ _06559_ VGND VGND VPWR VPWR _06560_ sky130_fd_sc_hd__nand2_1
X_13577_ _03526_ _03535_ VGND VGND VPWR VPWR _03536_ sky130_fd_sc_hd__and2_2
XFILLER_0_125_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10789_ _00664_ _00666_ VGND VGND VPWR VPWR _00728_ sky130_fd_sc_hd__xor2_2
X_15316_ net471 net162 net157 net476 VGND VGND VPWR VPWR _05406_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_82_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18104_ _07784_ _07790_ _07791_ _08472_ VGND VGND VPWR VPWR _08473_ sky130_fd_sc_hd__o31ai_2
X_12528_ _02358_ _02462_ VGND VGND VPWR VPWR _02467_ sky130_fd_sc_hd__and2_1
X_19084_ _09523_ _00516_ _09528_ net487 VGND VGND VPWR VPWR _00098_ sky130_fd_sc_hd__o211a_1
X_16296_ _06482_ _06483_ VGND VGND VPWR VPWR _06484_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15247_ _05327_ _05328_ _05329_ VGND VGND VPWR VPWR _05330_ sky130_fd_sc_hd__o21ba_1
X_18035_ _08377_ _08396_ net331 _07183_ VGND VGND VPWR VPWR _08397_ sky130_fd_sc_hd__and4b_1
X_12459_ _02335_ _02323_ VGND VGND VPWR VPWR _02398_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15178_ _05148_ _05152_ VGND VGND VPWR VPWR _05254_ sky130_fd_sc_hd__nor2_1
X_14129_ _04098_ _04041_ _04099_ _04100_ VGND VGND VPWR VPWR _04101_ sky130_fd_sc_hd__o211a_1
Xfanout309 net310 VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__buf_2
X_18937_ _02153_ VGND VGND VPWR VPWR _09389_ sky130_fd_sc_hd__inv_2
X_09670_ net57 _03625_ _03658_ ki\[8\] VGND VGND VPWR VPWR _00055_ sky130_fd_sc_hd__a22o_1
X_18868_ _09311_ _09312_ VGND VGND VPWR VPWR _09313_ sky130_fd_sc_hd__xor2_1
XFILLER_0_27_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17819_ _08154_ _08156_ VGND VGND VPWR VPWR _08159_ sky130_fd_sc_hd__or2b_1
X_18799_ _04131_ _04193_ _09236_ VGND VGND VPWR VPWR _09237_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_15_0_clock clknet_0_clock VGND VGND VPWR VPWR clknet_4_15_0_clock sky130_fd_sc_hd__clkbuf_8
XFILLER_0_150_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09937_ net338 _06645_ VGND VGND VPWR VPWR _06656_ sky130_fd_sc_hd__nand2_1
X_09868_ _04665_ _05886_ _04599_ VGND VGND VPWR VPWR _05897_ sky130_fd_sc_hd__a21o_2
X_09799_ _04170_ _04764_ _05127_ VGND VGND VPWR VPWR _05138_ sky130_fd_sc_hd__a21o_1
X_11830_ net242 net238 _01764_ VGND VGND VPWR VPWR _01769_ sky130_fd_sc_hd__nand3_1
XFILLER_0_68_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11761_ prev_error\[17\] _01699_ VGND VGND VPWR VPWR _01700_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13500_ _03415_ _03410_ _03414_ VGND VGND VPWR VPWR _03459_ sky130_fd_sc_hd__or3_1
X_10712_ _00627_ _00649_ VGND VGND VPWR VPWR _00651_ sky130_fd_sc_hd__and2_1
X_14480_ net461 net129 _04485_ VGND VGND VPWR VPWR _04486_ sky130_fd_sc_hd__and3_1
XFILLER_0_67_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11692_ _01629_ _01630_ VGND VGND VPWR VPWR _01631_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13431_ _03376_ _03379_ _03387_ VGND VGND VPWR VPWR _03389_ sky130_fd_sc_hd__nand3_1
X_10643_ _00486_ _00581_ VGND VGND VPWR VPWR _00582_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16150_ _06321_ _06322_ VGND VGND VPWR VPWR _06323_ sky130_fd_sc_hd__nor2_1
X_13362_ _03275_ _03314_ VGND VGND VPWR VPWR _03315_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10574_ _04225_ _04269_ _04203_ VGND VGND VPWR VPWR _00513_ sky130_fd_sc_hd__o21a_4
XFILLER_0_51_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15101_ _05074_ _05076_ VGND VGND VPWR VPWR _05169_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer8 net517 VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__buf_1
X_12313_ _02250_ _02251_ VGND VGND VPWR VPWR _02252_ sky130_fd_sc_hd__nor2b_2
X_16081_ _06212_ _06213_ _06217_ VGND VGND VPWR VPWR _06247_ sky130_fd_sc_hd__o21a_1
X_13293_ _03233_ _03245_ VGND VGND VPWR VPWR _03246_ sky130_fd_sc_hd__and2_1
X_15032_ _05084_ VGND VGND VPWR VPWR _05093_ sky130_fd_sc_hd__inv_2
X_12244_ _02181_ _02182_ VGND VGND VPWR VPWR _02183_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12175_ _02103_ _02105_ VGND VGND VPWR VPWR _02114_ sky130_fd_sc_hd__or2b_1
X_11126_ net378 _09558_ _09565_ VGND VGND VPWR VPWR _01065_ sky130_fd_sc_hd__and3_1
X_16983_ net282 _06891_ VGND VGND VPWR VPWR _07240_ sky130_fd_sc_hd__nand2_1
X_18722_ _09146_ _09145_ _06138_ VGND VGND VPWR VPWR _09152_ sky130_fd_sc_hd__a21o_1
X_15934_ _06085_ _03669_ VGND VGND VPWR VPWR _06086_ sky130_fd_sc_hd__xnor2_2
X_11057_ _00992_ _00993_ _00995_ VGND VGND VPWR VPWR _00996_ sky130_fd_sc_hd__o21a_1
X_10008_ net348 _04896_ VGND VGND VPWR VPWR _07437_ sky130_fd_sc_hd__nand2_1
X_18653_ _08962_ VGND VGND VPWR VPWR _09077_ sky130_fd_sc_hd__buf_4
X_15865_ _04300_ _04301_ _05999_ _06002_ VGND VGND VPWR VPWR _06010_ sky130_fd_sc_hd__a22o_1
X_17604_ _07920_ _07922_ VGND VGND VPWR VPWR _07923_ sky130_fd_sc_hd__nand2_1
X_14816_ _04845_ _04847_ _04855_ VGND VGND VPWR VPWR _04856_ sky130_fd_sc_hd__a21o_1
X_18584_ _08754_ _08755_ VGND VGND VPWR VPWR _09001_ sky130_fd_sc_hd__nand2_1
X_15796_ _05926_ _05893_ VGND VGND VPWR VPWR _05934_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17535_ _07846_ _07482_ VGND VGND VPWR VPWR _07847_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_157_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11959_ net213 _01835_ _01807_ net217 VGND VGND VPWR VPWR _01898_ sky130_fd_sc_hd__a22oi_1
X_14747_ _04747_ _04777_ _04779_ VGND VGND VPWR VPWR _04780_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_156_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14678_ net454 net143 _04702_ VGND VGND VPWR VPWR _04704_ sky130_fd_sc_hd__and3_1
X_17466_ _07311_ _07313_ VGND VGND VPWR VPWR _07771_ sky130_fd_sc_hd__xor2_2
XFILLER_0_27_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19205_ clknet_4_12_0_clock _00087_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13629_ _03587_ _03534_ VGND VGND VPWR VPWR _03588_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16417_ _06475_ _06477_ VGND VGND VPWR VPWR _06617_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_27_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17397_ _07609_ _07612_ _07608_ VGND VGND VPWR VPWR _07695_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_6_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19136_ net503 _09051_ VGND VGND VPWR VPWR _09561_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16348_ _06537_ _06540_ VGND VGND VPWR VPWR _06541_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16279_ net115 _06464_ _06292_ _01871_ VGND VGND VPWR VPWR _06465_ sky130_fd_sc_hd__a211o_2
X_19067_ _09515_ _09517_ VGND VGND VPWR VPWR _00090_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18018_ _08376_ _08377_ VGND VGND VPWR VPWR _08378_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout117 net118 VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_4
Xfanout128 net132 VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__buf_2
Xfanout139 net140 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_4
X_09722_ _04280_ _04192_ VGND VGND VPWR VPWR _04291_ sky130_fd_sc_hd__nand2_4
XFILLER_0_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09653_ net48 _03347_ _03380_ net201 VGND VGND VPWR VPWR _00008_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_118_Right_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10290_ net338 _09583_ _09595_ VGND VGND VPWR VPWR _00229_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13980_ _03950_ _03951_ VGND VGND VPWR VPWR _03952_ sky130_fd_sc_hd__and2_1
X_12931_ _02867_ _02869_ VGND VGND VPWR VPWR _02870_ sky130_fd_sc_hd__or2b_1
X_15650_ _05760_ _05764_ net447 net195 VGND VGND VPWR VPWR _05773_ sky130_fd_sc_hd__o211a_1
X_12862_ _02598_ _02799_ _02800_ VGND VGND VPWR VPWR _02801_ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14601_ _03917_ _04618_ VGND VGND VPWR VPWR _04619_ sky130_fd_sc_hd__xnor2_1
X_11813_ _01702_ _01750_ _01751_ VGND VGND VPWR VPWR _01752_ sky130_fd_sc_hd__a21oi_4
X_15581_ _05685_ _05694_ _05696_ VGND VGND VPWR VPWR _05697_ sky130_fd_sc_hd__a21o_1
X_12793_ _02718_ _02727_ _02716_ VGND VGND VPWR VPWR _02732_ sky130_fd_sc_hd__o21a_1
X_14532_ _04527_ _04529_ _04538_ VGND VGND VPWR VPWR _04543_ sky130_fd_sc_hd__or3_1
XFILLER_0_84_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17320_ net317 _06409_ VGND VGND VPWR VPWR _07610_ sky130_fd_sc_hd__nand2_2
X_11744_ _00868_ _00955_ VGND VGND VPWR VPWR _01683_ sky130_fd_sc_hd__and2_1
XFILLER_0_139_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14463_ _04370_ _04371_ _04372_ _04343_ VGND VGND VPWR VPWR _04468_ sky130_fd_sc_hd__a22o_1
X_17251_ net302 _06803_ _07507_ _07506_ VGND VGND VPWR VPWR _07534_ sky130_fd_sc_hd__a31o_1
X_11675_ net564 net385 _00810_ _00798_ VGND VGND VPWR VPWR _01614_ sky130_fd_sc_hd__and4_1
XFILLER_0_126_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13414_ net244 _02408_ VGND VGND VPWR VPWR _03371_ sky130_fd_sc_hd__nand2_2
X_16202_ net292 _06379_ VGND VGND VPWR VPWR _06380_ sky130_fd_sc_hd__nand2_1
X_17182_ _07454_ _07457_ VGND VGND VPWR VPWR _07458_ sky130_fd_sc_hd__xor2_2
X_10626_ _00527_ _00552_ VGND VGND VPWR VPWR _00565_ sky130_fd_sc_hd__xnor2_4
X_14394_ _04309_ _04391_ VGND VGND VPWR VPWR _04392_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16133_ _06297_ _06300_ _06303_ VGND VGND VPWR VPWR _06305_ sky130_fd_sc_hd__a21oi_4
X_13345_ _03278_ _03285_ _03286_ VGND VGND VPWR VPWR _03298_ sky130_fd_sc_hd__nand3_1
XFILLER_0_106_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10557_ _00483_ _00495_ VGND VGND VPWR VPWR _00496_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16064_ _06225_ _06228_ _06223_ VGND VGND VPWR VPWR _06229_ sky130_fd_sc_hd__a21oi_2
X_13276_ _03219_ _03228_ VGND VGND VPWR VPWR _03229_ sky130_fd_sc_hd__nor2_1
X_10488_ _00348_ _00426_ VGND VGND VPWR VPWR _00427_ sky130_fd_sc_hd__nand2_2
X_15015_ net414 net419 net197 net193 VGND VGND VPWR VPWR _05075_ sky130_fd_sc_hd__and4_1
X_12227_ _02163_ _02164_ VGND VGND VPWR VPWR _02166_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12158_ _02084_ _02095_ _02096_ VGND VGND VPWR VPWR _02097_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11109_ net396 _05963_ _05974_ _06172_ net392 VGND VGND VPWR VPWR _01048_ sky130_fd_sc_hd__a32oi_2
X_12089_ _02009_ _02026_ VGND VGND VPWR VPWR _02028_ sky130_fd_sc_hd__nand2_1
X_16966_ net566 _06307_ _06308_ VGND VGND VPWR VPWR _07221_ sky130_fd_sc_hd__and3_4
X_18705_ _09119_ _09122_ _09132_ _09133_ VGND VGND VPWR VPWR _09134_ sky130_fd_sc_hd__a31o_4
X_15917_ _05953_ _06066_ VGND VGND VPWR VPWR _06067_ sky130_fd_sc_hd__nor2_1
X_16897_ _07143_ _07144_ VGND VGND VPWR VPWR _07145_ sky130_fd_sc_hd__xor2_1
XFILLER_0_79_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18636_ _09056_ _09057_ VGND VGND VPWR VPWR _09058_ sky130_fd_sc_hd__nand2_1
X_15848_ _05989_ _05978_ VGND VGND VPWR VPWR _05991_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18567_ _08970_ _08980_ VGND VGND VPWR VPWR _08982_ sky130_fd_sc_hd__nand2_1
X_15779_ _05896_ _05914_ net483 net187 VGND VGND VPWR VPWR _05915_ sky130_fd_sc_hd__and4b_1
XFILLER_0_59_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17518_ _07826_ _07825_ VGND VGND VPWR VPWR _07828_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18498_ _08905_ _08858_ VGND VGND VPWR VPWR _08906_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17449_ _07750_ _07751_ VGND VGND VPWR VPWR _07752_ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19119_ net503 _09114_ _09115_ _09549_ VGND VGND VPWR VPWR _00115_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_15_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09705_ net49 _03870_ _03903_ net568 VGND VGND VPWR VPWR _00066_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09636_ net40 _03358_ _03391_ net269 VGND VGND VPWR VPWR _00000_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11460_ _01397_ _01398_ VGND VGND VPWR VPWR _01399_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10411_ _00271_ _00349_ VGND VGND VPWR VPWR _00350_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11391_ _01323_ _01329_ VGND VGND VPWR VPWR _01330_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13130_ _02973_ _02945_ _02972_ VGND VGND VPWR VPWR _03077_ sky130_fd_sc_hd__and3_1
X_10342_ net375 _05171_ _04885_ net379 VGND VGND VPWR VPWR _00281_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_104_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13061_ _02996_ _03000_ VGND VGND VPWR VPWR _03001_ sky130_fd_sc_hd__xor2_2
XFILLER_0_131_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10273_ _00206_ _00211_ VGND VGND VPWR VPWR _00212_ sky130_fd_sc_hd__or2b_1
X_12012_ _01802_ _01821_ _01950_ VGND VGND VPWR VPWR _01951_ sky130_fd_sc_hd__o21a_1
X_16820_ _07058_ _07059_ VGND VGND VPWR VPWR _07060_ sky130_fd_sc_hd__or2b_1
XPHY_EDGE_ROW_131_Left_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout470 net472 VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__buf_2
Xfanout481 net482 VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__clkbuf_2
X_16751_ net282 _06724_ _06983_ _06981_ VGND VGND VPWR VPWR _06984_ sky130_fd_sc_hd__a31o_1
Xfanout492 net493 VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__buf_2
X_13963_ _03933_ _03934_ VGND VGND VPWR VPWR _03935_ sky130_fd_sc_hd__nor2_1
X_15702_ _05813_ _05815_ VGND VGND VPWR VPWR _05830_ sky130_fd_sc_hd__xnor2_1
X_12914_ net204 _02747_ _02852_ _02850_ VGND VGND VPWR VPWR _02853_ sky130_fd_sc_hd__a31o_1
X_13894_ _03089_ _03177_ VGND VGND VPWR VPWR _03861_ sky130_fd_sc_hd__nand2_1
X_16682_ _06649_ _06785_ VGND VGND VPWR VPWR _06908_ sky130_fd_sc_hd__xnor2_1
X_18421_ _08785_ _08788_ _08819_ _08818_ VGND VGND VPWR VPWR _08821_ sky130_fd_sc_hd__a2bb2o_1
X_15633_ _05694_ _05753_ VGND VGND VPWR VPWR _05755_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12845_ net255 _01806_ _01812_ net259 VGND VGND VPWR VPWR _02784_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_69_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18352_ _08744_ VGND VGND VPWR VPWR _08745_ sky130_fd_sc_hd__inv_2
X_15564_ _05657_ _05678_ VGND VGND VPWR VPWR _05679_ sky130_fd_sc_hd__nand2_1
X_12776_ _02623_ _02714_ VGND VGND VPWR VPWR _02715_ sky130_fd_sc_hd__or2_1
XFILLER_0_139_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17303_ _07589_ _07590_ VGND VGND VPWR VPWR _07592_ sky130_fd_sc_hd__xor2_1
X_14515_ _04523_ _04518_ _04520_ VGND VGND VPWR VPWR _04525_ sky130_fd_sc_hd__nor3_1
X_11727_ _01461_ _01507_ _01663_ _01665_ VGND VGND VPWR VPWR _01666_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15495_ _05586_ _05601_ _05602_ VGND VGND VPWR VPWR _05603_ sky130_fd_sc_hd__nand3_2
X_18283_ _06534_ _06576_ _06574_ VGND VGND VPWR VPWR _08670_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_140_Left_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17234_ _07469_ _07471_ _07475_ VGND VGND VPWR VPWR _07516_ sky130_fd_sc_hd__and3_1
XFILLER_0_142_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14446_ _04443_ _04446_ _04448_ VGND VGND VPWR VPWR _04449_ sky130_fd_sc_hd__o21ai_1
X_11658_ net390 _00814_ _00612_ net394 VGND VGND VPWR VPWR _01597_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10609_ _00531_ _00546_ VGND VGND VPWR VPWR _00548_ sky130_fd_sc_hd__and2_1
X_17165_ _07435_ _07439_ VGND VGND VPWR VPWR _07440_ sky130_fd_sc_hd__xnor2_1
X_14377_ _04343_ _04370_ _04371_ _04372_ VGND VGND VPWR VPWR _04373_ sky130_fd_sc_hd__nand4_1
XFILLER_0_153_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11589_ net390 _00323_ _01488_ VGND VGND VPWR VPWR _01528_ sky130_fd_sc_hd__nand3_1
XFILLER_0_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13328_ net241 _02332_ _03182_ VGND VGND VPWR VPWR _03281_ sky130_fd_sc_hd__and3_1
X_16116_ prev_error\[6\] _00242_ VGND VGND VPWR VPWR _06286_ sky130_fd_sc_hd__and2_1
X_17096_ _07357_ _07363_ VGND VGND VPWR VPWR _07364_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_40_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16047_ _06198_ _06199_ _06209_ VGND VGND VPWR VPWR _06210_ sky130_fd_sc_hd__or3_1
X_13259_ _03206_ _03211_ VGND VGND VPWR VPWR _03212_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17998_ net326 _07156_ _08326_ VGND VGND VPWR VPWR _08356_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16949_ net302 _06468_ _06620_ net299 VGND VGND VPWR VPWR _07202_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18619_ _08907_ _09038_ _08964_ VGND VGND VPWR VPWR _09039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10960_ net337 _00818_ VGND VGND VPWR VPWR _00899_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09619_ net57 _03102_ _03135_ net160 VGND VGND VPWR VPWR _00036_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10891_ _00791_ _00789_ VGND VGND VPWR VPWR _00830_ sky130_fd_sc_hd__xnor2_1
X_12630_ _02470_ _02567_ VGND VGND VPWR VPWR _02569_ sky130_fd_sc_hd__and2_1
XFILLER_0_155_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12561_ _02426_ _02436_ VGND VGND VPWR VPWR _02500_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14300_ _04045_ _04287_ VGND VGND VPWR VPWR _04288_ sky130_fd_sc_hd__nor2_1
X_11512_ _01447_ _01442_ _01445_ VGND VGND VPWR VPWR _01451_ sky130_fd_sc_hd__nor3_1
XFILLER_0_93_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15280_ _05355_ _05357_ _05364_ VGND VGND VPWR VPWR _05366_ sky130_fd_sc_hd__and3_1
Xwire101 _06263_ VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__buf_4
X_12492_ net259 _01764_ net111 net254 VGND VGND VPWR VPWR _02431_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_80_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14231_ _04161_ _04211_ VGND VGND VPWR VPWR _04212_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11443_ _01380_ _01375_ VGND VGND VPWR VPWR _01382_ sky130_fd_sc_hd__and2b_1
XFILLER_0_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14162_ _04134_ _04135_ VGND VGND VPWR VPWR _04136_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11374_ _01311_ _01299_ _01310_ VGND VGND VPWR VPWR _01313_ sky130_fd_sc_hd__or3_1
XFILLER_0_22_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13113_ net220 _02544_ _03057_ VGND VGND VPWR VPWR _03059_ sky130_fd_sc_hd__a21boi_1
X_10325_ _00178_ _00179_ VGND VGND VPWR VPWR _00264_ sky130_fd_sc_hd__xor2_1
XFILLER_0_132_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14093_ _03950_ _04047_ _04064_ VGND VGND VPWR VPWR _04065_ sky130_fd_sc_hd__a21o_1
X_18970_ _09405_ _09424_ VGND VGND VPWR VPWR _09425_ sky130_fd_sc_hd__xnor2_2
X_13044_ _02875_ _02982_ VGND VGND VPWR VPWR _02983_ sky130_fd_sc_hd__nand2_1
X_17921_ _08224_ _08270_ VGND VGND VPWR VPWR _08271_ sky130_fd_sc_hd__xnor2_1
X_10256_ _09175_ _00194_ VGND VGND VPWR VPWR _00195_ sky130_fd_sc_hd__xnor2_1
X_17852_ _08087_ _08194_ VGND VGND VPWR VPWR _08195_ sky130_fd_sc_hd__xor2_1
X_10187_ _09340_ _09395_ VGND VGND VPWR VPWR _09406_ sky130_fd_sc_hd__nand2_1
X_16803_ _06937_ _07036_ _07040_ VGND VGND VPWR VPWR _07042_ sky130_fd_sc_hd__o21a_1
X_17783_ _08090_ _08095_ VGND VGND VPWR VPWR _08120_ sky130_fd_sc_hd__nand2_1
X_14995_ _04921_ _04924_ VGND VGND VPWR VPWR _05053_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16734_ _06959_ _06965_ VGND VGND VPWR VPWR _06966_ sky130_fd_sc_hd__xor2_1
X_13946_ net470 net475 net118 VGND VGND VPWR VPWR _03918_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16665_ _06889_ VGND VGND VPWR VPWR _06890_ sky130_fd_sc_hd__buf_4
X_13877_ _03785_ _03809_ _03841_ _03842_ VGND VGND VPWR VPWR _03843_ sky130_fd_sc_hd__a31o_1
X_18404_ _06153_ _08802_ VGND VGND VPWR VPWR _08803_ sky130_fd_sc_hd__or2_1
X_15616_ _05727_ _05735_ VGND VGND VPWR VPWR _05736_ sky130_fd_sc_hd__and2_1
X_12828_ _02764_ _02766_ VGND VGND VPWR VPWR _02767_ sky130_fd_sc_hd__or2b_1
XFILLER_0_146_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16596_ _06726_ _06725_ VGND VGND VPWR VPWR _06814_ sky130_fd_sc_hd__and2b_1
XFILLER_0_56_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18335_ _08688_ _08726_ VGND VGND VPWR VPWR _08727_ sky130_fd_sc_hd__xnor2_1
X_15547_ _05659_ VGND VGND VPWR VPWR _05660_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12759_ net268 _01813_ VGND VGND VPWR VPWR _02698_ sky130_fd_sc_hd__and2_1
X_18266_ _06507_ _06528_ _06526_ VGND VGND VPWR VPWR _08651_ sky130_fd_sc_hd__a21oi_1
X_15478_ _05488_ _05500_ _05499_ VGND VGND VPWR VPWR _05584_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17217_ _07484_ _07487_ VGND VGND VPWR VPWR _07497_ sky130_fd_sc_hd__and2b_1
X_14429_ _04427_ _04429_ VGND VGND VPWR VPWR _04430_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18197_ _08572_ _08573_ _08494_ VGND VGND VPWR VPWR _08575_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17148_ _07407_ _07420_ VGND VGND VPWR VPWR _07421_ sky130_fd_sc_hd__xnor2_2
Xfanout8 _04137_ VGND VGND VPWR VPWR net563 sky130_fd_sc_hd__buf_4
X_09970_ net338 _06073_ _06315_ _06304_ VGND VGND VPWR VPWR _07019_ sky130_fd_sc_hd__a31o_1
XFILLER_0_150_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17079_ _07332_ _07333_ _07343_ VGND VGND VPWR VPWR _07345_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10110_ net339 _05754_ VGND VGND VPWR VPWR _08559_ sky130_fd_sc_hd__nand2_1
X_11090_ net340 _00812_ VGND VGND VPWR VPWR _01029_ sky130_fd_sc_hd__nand2_1
X_10041_ _05644_ _07789_ VGND VGND VPWR VPWR _07800_ sky130_fd_sc_hd__xor2_1
Xhold42 net83 VGND VGND VPWR VPWR net549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 i_error\[16\] VGND VGND VPWR VPWR net560 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13800_ _03760_ _03765_ VGND VGND VPWR VPWR _03766_ sky130_fd_sc_hd__nor2_1
X_11992_ net231 kd_1\[10\] VGND VGND VPWR VPWR _01931_ sky130_fd_sc_hd__or2_1
X_14780_ _04803_ _04806_ _04815_ VGND VGND VPWR VPWR _04816_ sky130_fd_sc_hd__o21ai_1
X_13731_ _03695_ _03696_ VGND VGND VPWR VPWR _03697_ sky130_fd_sc_hd__and2_1
X_10943_ _00878_ _00881_ VGND VGND VPWR VPWR _00882_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16450_ _06651_ _06652_ VGND VGND VPWR VPWR _06653_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13662_ net243 _02913_ VGND VGND VPWR VPWR _03624_ sky130_fd_sc_hd__nand2_1
X_10874_ _04236_ _04247_ VGND VGND VPWR VPWR _00813_ sky130_fd_sc_hd__xor2_4
XFILLER_0_39_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15401_ _05494_ _05498_ VGND VGND VPWR VPWR _05499_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12613_ _02540_ _02551_ VGND VGND VPWR VPWR _02552_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13593_ _03498_ _03496_ VGND VGND VPWR VPWR _03552_ sky130_fd_sc_hd__xnor2_1
X_16381_ _06534_ _06576_ VGND VGND VPWR VPWR _06577_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18120_ _08488_ _08489_ VGND VGND VPWR VPWR _08490_ sky130_fd_sc_hd__and2b_1
X_12544_ _02479_ _02482_ VGND VGND VPWR VPWR _02483_ sky130_fd_sc_hd__xor2_1
X_15332_ _05340_ _05339_ VGND VGND VPWR VPWR _05423_ sky130_fd_sc_hd__nor2_1
X_18051_ _08406_ _08410_ _08413_ VGND VGND VPWR VPWR _08414_ sky130_fd_sc_hd__and3_1
X_12475_ _02411_ _02413_ VGND VGND VPWR VPWR _02414_ sky130_fd_sc_hd__nor2_1
X_15263_ _05273_ _05272_ VGND VGND VPWR VPWR _05348_ sky130_fd_sc_hd__and2b_1
XFILLER_0_81_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17002_ _07253_ _07257_ _07259_ VGND VGND VPWR VPWR _07260_ sky130_fd_sc_hd__o21ai_1
X_14214_ _04191_ _04193_ VGND VGND VPWR VPWR _04194_ sky130_fd_sc_hd__or2_1
X_11426_ net374 _00514_ VGND VGND VPWR VPWR _01365_ sky130_fd_sc_hd__nand2_1
X_15194_ net427 net194 net189 net433 VGND VGND VPWR VPWR _05272_ sky130_fd_sc_hd__a22o_1
XANTENNA_6 _06544_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14145_ _04105_ _04056_ _04117_ VGND VGND VPWR VPWR _04118_ sky130_fd_sc_hd__a21o_1
X_11357_ _01289_ _01295_ VGND VGND VPWR VPWR _01296_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10308_ kp\[15\] _09558_ _09565_ VGND VGND VPWR VPWR _00247_ sky130_fd_sc_hd__and3_1
X_14076_ _03944_ _03946_ _03945_ VGND VGND VPWR VPWR _04048_ sky130_fd_sc_hd__o21ba_1
X_18953_ _09264_ _09265_ VGND VGND VPWR VPWR _09407_ sky130_fd_sc_hd__nand2_1
X_11288_ _01224_ _01226_ VGND VGND VPWR VPWR _01227_ sky130_fd_sc_hd__or2b_1
XFILLER_0_120_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13027_ _02961_ _02965_ VGND VGND VPWR VPWR _02966_ sky130_fd_sc_hd__and2_1
X_17904_ _08243_ _08232_ _08242_ VGND VGND VPWR VPWR _08253_ sky130_fd_sc_hd__nor3_1
X_10239_ _09472_ _00160_ _09450_ VGND VGND VPWR VPWR _00178_ sky130_fd_sc_hd__o21ai_2
X_18884_ _02119_ _02167_ _02165_ VGND VGND VPWR VPWR _09331_ sky130_fd_sc_hd__a21oi_1
X_17835_ net322 _06991_ VGND VGND VPWR VPWR _08177_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17766_ _08072_ _08074_ VGND VGND VPWR VPWR _08101_ sky130_fd_sc_hd__nand2_1
Xrebuffer18 _08897_ VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__clkbuf_1
X_14978_ _05026_ _05032_ _05020_ VGND VGND VPWR VPWR _05034_ sky130_fd_sc_hd__a21o_1
X_16717_ _06944_ _06946_ VGND VGND VPWR VPWR _06947_ sky130_fd_sc_hd__nand2_1
X_13929_ _03897_ _03898_ VGND VGND VPWR VPWR _03899_ sky130_fd_sc_hd__nor2_1
X_17697_ _08016_ _08021_ _08024_ VGND VGND VPWR VPWR _08025_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_89_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16648_ _06860_ _06866_ _06870_ VGND VGND VPWR VPWR _06871_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_146_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16579_ _06792_ _06794_ VGND VGND VPWR VPWR _06795_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_146_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18318_ _08689_ _08707_ VGND VGND VPWR VPWR _08708_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19298_ clknet_4_3_0_clock _00056_ VGND VGND VPWR VPWR ki\[9\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_155_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18249_ ki\[14\] _06311_ _06562_ _06561_ _06379_ VGND VGND VPWR VPWR _08632_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09953_ net357 net353 _04896_ _05006_ VGND VGND VPWR VPWR _06832_ sky130_fd_sc_hd__and4_1
XFILLER_0_148_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09884_ _06062_ VGND VGND VPWR VPWR _06073_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_4_11_0_clock clknet_0_clock VGND VGND VPWR VPWR clknet_4_11_0_clock sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10590_ _00483_ _00495_ VGND VGND VPWR VPWR _00529_ sky130_fd_sc_hd__xor2_2
XFILLER_0_146_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12260_ _02196_ _02198_ VGND VGND VPWR VPWR _02199_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11211_ _01148_ _01149_ VGND VGND VPWR VPWR _01150_ sky130_fd_sc_hd__and2b_1
X_12191_ _02128_ _02129_ VGND VGND VPWR VPWR _02130_ sky130_fd_sc_hd__xnor2_1
X_11142_ _01061_ _01078_ _01079_ _01080_ VGND VGND VPWR VPWR _01081_ sky130_fd_sc_hd__a211o_2
XFILLER_0_102_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput87 net87 VGND VGND VPWR VPWR out_clocked[16] sky130_fd_sc_hd__clkbuf_4
X_15950_ _06070_ _06101_ _06102_ VGND VGND VPWR VPWR _06103_ sky130_fd_sc_hd__a21o_1
X_11073_ _00989_ _00990_ _00975_ _00988_ VGND VGND VPWR VPWR _01012_ sky130_fd_sc_hd__o211a_1
Xoutput98 net98 VGND VGND VPWR VPWR out_clocked[9] sky130_fd_sc_hd__buf_2
X_10024_ _06777_ _07602_ VGND VGND VPWR VPWR _07613_ sky130_fd_sc_hd__and2_1
X_14901_ _04946_ _04938_ _04944_ VGND VGND VPWR VPWR _04949_ sky130_fd_sc_hd__and3_1
X_15881_ _05987_ _06026_ VGND VGND VPWR VPWR _06027_ sky130_fd_sc_hd__xnor2_1
X_17620_ _07936_ _07939_ _07934_ VGND VGND VPWR VPWR _07940_ sky130_fd_sc_hd__a21oi_2
X_14832_ _04871_ _04872_ VGND VGND VPWR VPWR _04873_ sky130_fd_sc_hd__nand2_1
X_17551_ _07515_ _07860_ _07854_ _07859_ VGND VGND VPWR VPWR _07864_ sky130_fd_sc_hd__o211a_1
X_14763_ _04795_ _04796_ net479 net124 VGND VGND VPWR VPWR _04798_ sky130_fd_sc_hd__and4b_1
X_11975_ net200 _01910_ _01911_ _01913_ VGND VGND VPWR VPWR _01914_ sky130_fd_sc_hd__and4_1
XFILLER_0_98_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16502_ _06626_ _06638_ VGND VGND VPWR VPWR _06710_ sky130_fd_sc_hd__xnor2_1
X_13714_ net267 _02639_ VGND VGND VPWR VPWR _03680_ sky130_fd_sc_hd__nand2_1
X_10926_ _00662_ _00754_ VGND VGND VPWR VPWR _00865_ sky130_fd_sc_hd__xor2_4
X_17482_ _07786_ _07787_ VGND VGND VPWR VPWR _07788_ sky130_fd_sc_hd__xor2_1
X_14694_ net439 net155 _04517_ VGND VGND VPWR VPWR _04722_ sky130_fd_sc_hd__and3_1
X_19221_ clknet_4_4_0_clock _00103_ VGND VGND VPWR VPWR prev_error\[8\] sky130_fd_sc_hd__dfxtp_1
X_16433_ _06471_ _06633_ VGND VGND VPWR VPWR _06635_ sky130_fd_sc_hd__xnor2_1
X_13645_ _03605_ VGND VGND VPWR VPWR _03606_ sky130_fd_sc_hd__inv_2
X_10857_ _00793_ _00795_ VGND VGND VPWR VPWR _00796_ sky130_fd_sc_hd__xor2_4
XFILLER_0_156_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19152_ net505 _09348_ VGND VGND VPWR VPWR _09570_ sky130_fd_sc_hd__nand2_1
X_16364_ net292 _06325_ VGND VGND VPWR VPWR _06559_ sky130_fd_sc_hd__nand2_1
X_13576_ _03505_ _03527_ _03534_ _03533_ _03529_ VGND VGND VPWR VPWR _03535_ sky130_fd_sc_hd__a32o_1
XFILLER_0_82_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10788_ _00642_ _00641_ _00636_ VGND VGND VPWR VPWR _00727_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_137_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18103_ _07782_ _07793_ VGND VGND VPWR VPWR _08472_ sky130_fd_sc_hd__or2b_1
X_15315_ net471 net477 net162 net157 VGND VGND VPWR VPWR _05405_ sky130_fd_sc_hd__and4_1
XFILLER_0_124_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12527_ _02464_ _02465_ VGND VGND VPWR VPWR _02466_ sky130_fd_sc_hd__or2_2
XFILLER_0_42_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19083_ net498 prev_error\[3\] VGND VGND VPWR VPWR _09528_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16295_ _06481_ _06462_ _06478_ VGND VGND VPWR VPWR _06483_ sky130_fd_sc_hd__nor3_1
XFILLER_0_23_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18034_ _06538_ _03065_ _08395_ VGND VGND VPWR VPWR _08396_ sky130_fd_sc_hd__o21ai_1
X_15246_ net453 net459 net172 net166 VGND VGND VPWR VPWR _05329_ sky130_fd_sc_hd__and4_1
XFILLER_0_140_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12458_ _02395_ _02396_ VGND VGND VPWR VPWR _02397_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11409_ _01244_ _01277_ _01276_ VGND VGND VPWR VPWR _01348_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15177_ _05231_ _05233_ VGND VGND VPWR VPWR _05253_ sky130_fd_sc_hd__or2b_1
X_12389_ _01710_ _02327_ VGND VGND VPWR VPWR _02328_ sky130_fd_sc_hd__nand2_4
XFILLER_0_22_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14128_ _04095_ _04096_ _03988_ net113 VGND VGND VPWR VPWR _04100_ sky130_fd_sc_hd__a211o_1
X_14059_ _04029_ _04030_ VGND VGND VPWR VPWR _04031_ sky130_fd_sc_hd__and2_1
X_18936_ _09383_ _09387_ VGND VGND VPWR VPWR _09388_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18867_ net210 _01930_ VGND VGND VPWR VPWR _09312_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17818_ _08145_ _08147_ _08156_ _08157_ VGND VGND VPWR VPWR _08158_ sky130_fd_sc_hd__o211ai_4
X_18798_ _09232_ _09235_ VGND VGND VPWR VPWR _09236_ sky130_fd_sc_hd__xnor2_1
X_17749_ _08071_ _08081_ VGND VGND VPWR VPWR _08082_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09936_ _06634_ VGND VGND VPWR VPWR _06645_ sky130_fd_sc_hd__clkbuf_4
X_09867_ _04423_ _04500_ _04533_ _04643_ VGND VGND VPWR VPWR _05886_ sky130_fd_sc_hd__a211o_1
X_09798_ _04775_ _04159_ VGND VGND VPWR VPWR _05127_ sky130_fd_sc_hd__or2b_2
XFILLER_0_96_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11760_ _04973_ VGND VGND VPWR VPWR _01699_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10711_ _00627_ _00649_ VGND VGND VPWR VPWR _00650_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11691_ _01628_ _01626_ VGND VGND VPWR VPWR _01630_ sky130_fd_sc_hd__and2b_1
XFILLER_0_153_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13430_ _03376_ _03379_ _03387_ VGND VGND VPWR VPWR _03388_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10642_ _00382_ _00488_ _00487_ VGND VGND VPWR VPWR _00581_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13361_ net248 _02090_ _03274_ VGND VGND VPWR VPWR _03314_ sky130_fd_sc_hd__a21oi_1
X_10573_ _00507_ _00511_ VGND VGND VPWR VPWR _00512_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15100_ _05140_ net114 _05167_ VGND VGND VPWR VPWR _05168_ sky130_fd_sc_hd__o21a_1
X_12312_ _02115_ _02113_ VGND VGND VPWR VPWR _02251_ sky130_fd_sc_hd__xnor2_1
Xrebuffer9 _08549_ VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__buf_1
X_16080_ _06177_ _06195_ _06198_ VGND VGND VPWR VPWR _06246_ sky130_fd_sc_hd__a21o_1
X_13292_ _03236_ _03240_ _03244_ VGND VGND VPWR VPWR _03245_ sky130_fd_sc_hd__a21o_1
XFILLER_0_122_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12243_ _01768_ _02180_ VGND VGND VPWR VPWR _02182_ sky130_fd_sc_hd__nand2_1
X_15031_ _05002_ _05091_ VGND VGND VPWR VPWR _05092_ sky130_fd_sc_hd__or2b_1
X_12174_ _02032_ _02112_ VGND VGND VPWR VPWR _02113_ sky130_fd_sc_hd__xor2_1
XFILLER_0_102_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11125_ net374 _09577_ _08185_ net378 VGND VGND VPWR VPWR _01064_ sky130_fd_sc_hd__a22oi_1
X_16982_ _07236_ _07237_ VGND VGND VPWR VPWR _07238_ sky130_fd_sc_hd__and2_1
X_18721_ _06138_ _09146_ _09145_ VGND VGND VPWR VPWR _09151_ sky130_fd_sc_hd__nand3_1
XFILLER_0_3_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15933_ _03554_ _03667_ _03847_ VGND VGND VPWR VPWR _06085_ sky130_fd_sc_hd__or3b_1
X_11056_ _00891_ _00994_ VGND VGND VPWR VPWR _00995_ sky130_fd_sc_hd__xnor2_1
X_10007_ _06876_ _06920_ _06942_ _06887_ VGND VGND VPWR VPWR _07426_ sky130_fd_sc_hd__a31o_1
X_18652_ _08961_ VGND VGND VPWR VPWR _09075_ sky130_fd_sc_hd__buf_4
X_15864_ _06003_ VGND VGND VPWR VPWR _06009_ sky130_fd_sc_hd__inv_2
X_17603_ _07856_ _07858_ VGND VGND VPWR VPWR _07922_ sky130_fd_sc_hd__xor2_2
X_14815_ _04752_ _04771_ VGND VGND VPWR VPWR _04855_ sky130_fd_sc_hd__xnor2_1
X_18583_ _06120_ _06028_ _06119_ VGND VGND VPWR VPWR _09000_ sky130_fd_sc_hd__and3_2
X_15795_ _05891_ _05931_ _05932_ VGND VGND VPWR VPWR _05933_ sky130_fd_sc_hd__and3_1
XFILLER_0_86_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17534_ net328 _06400_ VGND VGND VPWR VPWR _07846_ sky130_fd_sc_hd__nand2_1
X_14746_ _04661_ _04778_ VGND VGND VPWR VPWR _04779_ sky130_fd_sc_hd__nor2_1
X_11958_ net217 net213 _01835_ _01807_ VGND VGND VPWR VPWR _01897_ sky130_fd_sc_hd__and4_1
XFILLER_0_59_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10909_ _00845_ _00847_ VGND VGND VPWR VPWR _00848_ sky130_fd_sc_hd__or2b_1
X_17465_ _07697_ _07709_ VGND VGND VPWR VPWR _07770_ sky130_fd_sc_hd__or2_1
X_14677_ net454 net143 _04702_ VGND VGND VPWR VPWR _04703_ sky130_fd_sc_hd__a21oi_1
X_11889_ net230 net226 _01786_ _01799_ VGND VGND VPWR VPWR _01828_ sky130_fd_sc_hd__and4_1
XFILLER_0_157_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19204_ clknet_4_12_0_clock _00086_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dfxtp_1
X_16416_ _06613_ _06615_ VGND VGND VPWR VPWR _06616_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_129_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13628_ _03505_ _03527_ VGND VGND VPWR VPWR _03587_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_17_Left_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17396_ _07604_ _07614_ _07615_ VGND VGND VPWR VPWR _07694_ sky130_fd_sc_hd__nand3_1
X_19135_ _09559_ _09066_ _09560_ net494 VGND VGND VPWR VPWR _00122_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16347_ _06538_ _06539_ _06321_ _06322_ VGND VGND VPWR VPWR _06540_ sky130_fd_sc_hd__or4_2
XFILLER_0_14_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13559_ _03515_ _03517_ VGND VGND VPWR VPWR _03518_ sky130_fd_sc_hd__xor2_1
XFILLER_0_70_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19066_ net505 net545 net495 VGND VGND VPWR VPWR _09517_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16278_ _06273_ _02087_ _06287_ _06291_ VGND VGND VPWR VPWR _06464_ sky130_fd_sc_hd__a31o_2
XFILLER_0_30_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18017_ net327 net322 _02932_ _07570_ VGND VGND VPWR VPWR _08377_ sky130_fd_sc_hd__and4_1
X_15229_ net468 net158 net140 net486 VGND VGND VPWR VPWR _05310_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_112_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout118 kd_2\[18\] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_2
Xfanout129 kd_2\[15\] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_26_Left_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09721_ net72 net14 VGND VGND VPWR VPWR _04280_ sky130_fd_sc_hd__nand2b_2
X_18919_ _09287_ _09297_ _09294_ VGND VGND VPWR VPWR _09369_ sky130_fd_sc_hd__a21oi_1
X_09652_ net47 _03347_ _03380_ net203 VGND VGND VPWR VPWR _00007_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_35_Left_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09919_ _06238_ _06260_ VGND VGND VPWR VPWR _06458_ sky130_fd_sc_hd__xnor2_1
X_12930_ _02758_ _02837_ _02838_ _02868_ VGND VGND VPWR VPWR _02869_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_34_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12861_ net243 _01860_ _01834_ net247 VGND VGND VPWR VPWR _02800_ sky130_fd_sc_hd__a22o_1
X_14600_ _04598_ _04600_ VGND VGND VPWR VPWR _04618_ sky130_fd_sc_hd__nor2_1
X_11812_ _01701_ _04896_ VGND VGND VPWR VPWR _01751_ sky130_fd_sc_hd__nor2_1
X_15580_ _05648_ _05695_ VGND VGND VPWR VPWR _05696_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12792_ _02711_ _02730_ VGND VGND VPWR VPWR _02731_ sky130_fd_sc_hd__and2_1
XFILLER_0_157_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14531_ _04540_ _04541_ net409 net182 VGND VGND VPWR VPWR _04542_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11743_ _01131_ _01132_ VGND VGND VPWR VPWR _01682_ sky130_fd_sc_hd__or2_2
X_17250_ _07530_ _07531_ _07517_ VGND VGND VPWR VPWR _07533_ sky130_fd_sc_hd__a21oi_1
X_14462_ _04463_ _04465_ VGND VGND VPWR VPWR _04466_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11674_ _01604_ _01605_ VGND VGND VPWR VPWR _01613_ sky130_fd_sc_hd__and2_1
X_16201_ _06320_ VGND VGND VPWR VPWR _06379_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13413_ net244 _02331_ _02409_ net239 VGND VGND VPWR VPWR _03370_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17181_ _07428_ _07455_ _07456_ VGND VGND VPWR VPWR _07457_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_64_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10625_ _00556_ _00554_ VGND VGND VPWR VPWR _00564_ sky130_fd_sc_hd__xor2_1
X_14393_ net448 net128 _04307_ _04308_ VGND VGND VPWR VPWR _04391_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_4_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16132_ _06299_ _01811_ _06302_ VGND VGND VPWR VPWR _06303_ sky130_fd_sc_hd__and3_1
X_13344_ _03293_ _03295_ _03296_ VGND VGND VPWR VPWR _03297_ sky130_fd_sc_hd__a21o_1
X_10556_ _00492_ _00494_ _00490_ VGND VGND VPWR VPWR _00495_ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16063_ _09131_ _00186_ _01696_ _06226_ _09120_ VGND VGND VPWR VPWR _06228_ sky130_fd_sc_hd__a32o_1
X_13275_ _03225_ _03227_ VGND VGND VPWR VPWR _03228_ sky130_fd_sc_hd__nand2_1
X_10487_ _00346_ _00347_ VGND VGND VPWR VPWR _00426_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15014_ _05069_ _05073_ VGND VGND VPWR VPWR _05074_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12226_ _02163_ _02164_ VGND VGND VPWR VPWR _02165_ sky130_fd_sc_hd__nor2_1
X_12157_ _02080_ _02082_ VGND VGND VPWR VPWR _02096_ sky130_fd_sc_hd__xnor2_1
X_11108_ net402 _06051_ VGND VGND VPWR VPWR _01047_ sky130_fd_sc_hd__nand2_1
X_12088_ _02009_ _02026_ VGND VGND VPWR VPWR _02027_ sky130_fd_sc_hd__nor2_1
X_16965_ net333 _06314_ _06317_ _06309_ net330 VGND VGND VPWR VPWR _07220_ sky130_fd_sc_hd__a32o_1
X_15916_ _05951_ _05465_ _05950_ VGND VGND VPWR VPWR _06066_ sky130_fd_sc_hd__and3_1
X_18704_ _09104_ _09107_ _09118_ VGND VGND VPWR VPWR _09133_ sky130_fd_sc_hd__and3_1
X_11039_ net370 _08207_ VGND VGND VPWR VPWR _00978_ sky130_fd_sc_hd__nand2_1
X_16896_ _07029_ _07031_ VGND VGND VPWR VPWR _07144_ sky130_fd_sc_hd__xnor2_1
X_18635_ _09046_ _09055_ VGND VGND VPWR VPWR _09057_ sky130_fd_sc_hd__nand2_1
X_15847_ _05989_ _05978_ VGND VGND VPWR VPWR _05990_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18566_ _08970_ _08980_ VGND VGND VPWR VPWR _08981_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15778_ net473 net196 _05895_ VGND VGND VPWR VPWR _05914_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17517_ _07825_ _07826_ VGND VGND VPWR VPWR _07827_ sky130_fd_sc_hd__and2b_1
XFILLER_0_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14729_ net413 net186 _04565_ VGND VGND VPWR VPWR _04760_ sky130_fd_sc_hd__and3_1
XFILLER_0_157_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18497_ _06266_ _08860_ VGND VGND VPWR VPWR _08905_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17448_ _07747_ _07749_ VGND VGND VPWR VPWR _07751_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17379_ _07589_ _07590_ VGND VGND VPWR VPWR _07675_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19118_ net503 net555 net494 VGND VGND VPWR VPWR _09549_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19049_ net522 _09485_ _09464_ VGND VGND VPWR VPWR _09504_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_151_Right_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09704_ net48 _03870_ _03903_ net337 VGND VGND VPWR VPWR _00065_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09635_ _03380_ VGND VGND VPWR VPWR _03391_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_43_Left_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10410_ _00273_ _00314_ _00348_ VGND VGND VPWR VPWR _00349_ sky130_fd_sc_hd__o21a_1
X_11390_ _01325_ _01326_ _01327_ _01328_ VGND VGND VPWR VPWR _01329_ sky130_fd_sc_hd__or4b_1
XFILLER_0_6_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10341_ net372 _05424_ VGND VGND VPWR VPWR _00280_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_52_Left_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13060_ net266 _01806_ _02997_ _02999_ VGND VGND VPWR VPWR _03000_ sky130_fd_sc_hd__a31o_1
X_10272_ _00207_ _00208_ _00210_ VGND VGND VPWR VPWR _00211_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_29_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12011_ _01948_ _01949_ VGND VGND VPWR VPWR _01950_ sky130_fd_sc_hd__nor2_1
Xfanout460 prev_d_error\[6\] VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__buf_2
Xfanout471 net472 VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__buf_2
X_16750_ _06981_ _06982_ VGND VGND VPWR VPWR _06983_ sky130_fd_sc_hd__nor2_1
Xfanout482 prev_d_error\[1\] VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__clkbuf_2
X_13962_ net421 net138 _03931_ _03932_ VGND VGND VPWR VPWR _03934_ sky130_fd_sc_hd__o2bb2a_1
Xfanout493 net497 VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__dlymetal6s2s_1
X_15701_ _05796_ _05828_ VGND VGND VPWR VPWR _05829_ sky130_fd_sc_hd__xnor2_1
X_12913_ _02850_ _02851_ VGND VGND VPWR VPWR _02852_ sky130_fd_sc_hd__nor2_1
X_16681_ _06872_ _06906_ VGND VGND VPWR VPWR _06907_ sky130_fd_sc_hd__or2_1
X_13893_ _03339_ _03857_ _03268_ _03858_ VGND VGND VPWR VPWR _03860_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_69_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18420_ _08810_ _08815_ _08818_ _08819_ VGND VGND VPWR VPWR _08820_ sky130_fd_sc_hd__o2bb2a_1
X_15632_ _05691_ _05693_ VGND VGND VPWR VPWR _05753_ sky130_fd_sc_hd__or2_1
X_12844_ net261 net255 _01806_ _01812_ VGND VGND VPWR VPWR _02783_ sky130_fd_sc_hd__and4_1
XFILLER_0_152_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18351_ _08617_ _08741_ _08743_ VGND VGND VPWR VPWR _08744_ sky130_fd_sc_hd__a21o_1
XFILLER_0_139_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15563_ _05652_ _05656_ VGND VGND VPWR VPWR _05678_ sky130_fd_sc_hd__or2_1
X_12775_ _02620_ _02622_ VGND VGND VPWR VPWR _02714_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17302_ net288 _07095_ VGND VGND VPWR VPWR _07590_ sky130_fd_sc_hd__nand2_2
X_14514_ _04518_ _04520_ _04523_ VGND VGND VPWR VPWR _04524_ sky130_fd_sc_hd__o21a_1
XFILLER_0_139_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11726_ _01508_ _01662_ _01664_ VGND VGND VPWR VPWR _01665_ sky130_fd_sc_hd__o21ai_1
X_18282_ _08653_ _08667_ VGND VGND VPWR VPWR _08668_ sky130_fd_sc_hd__xor2_1
X_15494_ _05585_ _05568_ _05583_ VGND VGND VPWR VPWR _05602_ sky130_fd_sc_hd__nand3_1
XFILLER_0_44_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17233_ _07499_ _07512_ _07513_ VGND VGND VPWR VPWR _07515_ sky130_fd_sc_hd__nor3_4
XFILLER_0_153_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14445_ _04353_ _04447_ VGND VGND VPWR VPWR _04448_ sky130_fd_sc_hd__nor2_1
X_11657_ net399 _00798_ _01556_ _01557_ VGND VGND VPWR VPWR _01596_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17164_ _07436_ _07438_ VGND VGND VPWR VPWR _07439_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10608_ _00531_ _00546_ VGND VGND VPWR VPWR _00547_ sky130_fd_sc_hd__xor2_1
X_14376_ _04342_ _04318_ _04341_ VGND VGND VPWR VPWR _04372_ sky130_fd_sc_hd__nand3_1
X_11588_ _01492_ _01491_ _01483_ VGND VGND VPWR VPWR _01527_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16115_ _02406_ _06283_ _06284_ VGND VGND VPWR VPWR _06285_ sky130_fd_sc_hd__a21o_2
X_13327_ _03279_ _03182_ VGND VGND VPWR VPWR _03280_ sky130_fd_sc_hd__xnor2_1
X_17095_ _07358_ _07362_ VGND VGND VPWR VPWR _07363_ sky130_fd_sc_hd__xnor2_2
X_10539_ net376 _05413_ _00477_ VGND VGND VPWR VPWR _00478_ sky130_fd_sc_hd__and3_1
XFILLER_0_150_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16046_ _06200_ _06208_ VGND VGND VPWR VPWR _06209_ sky130_fd_sc_hd__xnor2_1
X_13258_ _03207_ _03210_ _03208_ VGND VGND VPWR VPWR _03211_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12209_ net218 net215 _01772_ VGND VGND VPWR VPWR _02148_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13189_ _03019_ _03020_ VGND VGND VPWR VPWR _03142_ sky130_fd_sc_hd__xnor2_2
X_17997_ _08352_ _08353_ _08354_ VGND VGND VPWR VPWR _08355_ sky130_fd_sc_hd__o21ba_1
X_16948_ net297 _06721_ VGND VGND VPWR VPWR _07201_ sky130_fd_sc_hd__nand2_1
X_16879_ _07123_ _07124_ VGND VGND VPWR VPWR _07125_ sky130_fd_sc_hd__or2b_1
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18618_ _09037_ _08853_ _08882_ VGND VGND VPWR VPWR _09038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18549_ _08885_ _08730_ VGND VGND VPWR VPWR _08962_ sky130_fd_sc_hd__nand2_2
XFILLER_0_75_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09618_ net56 _03102_ _03135_ net165 VGND VGND VPWR VPWR _00035_ sky130_fd_sc_hd__a22o_1
X_10890_ _00723_ _00744_ VGND VGND VPWR VPWR _00829_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_156_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12560_ _02497_ _02498_ VGND VGND VPWR VPWR _02499_ sky130_fd_sc_hd__or2b_1
XFILLER_0_109_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11511_ _01431_ _01449_ VGND VGND VPWR VPWR _01450_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12491_ _02429_ VGND VGND VPWR VPWR _02430_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14230_ _04209_ _04210_ VGND VGND VPWR VPWR _04211_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11442_ _01375_ _01380_ VGND VGND VPWR VPWR _01381_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14161_ net422 net123 _04133_ VGND VGND VPWR VPWR _04135_ sky130_fd_sc_hd__a21oi_1
X_11373_ _01299_ _01310_ _01311_ VGND VGND VPWR VPWR _01312_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_150_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13112_ net216 _02639_ VGND VGND VPWR VPWR _03057_ sky130_fd_sc_hd__nand2_1
X_10324_ _00187_ _00258_ _00262_ VGND VGND VPWR VPWR _00263_ sky130_fd_sc_hd__o21ba_1
X_14092_ _04062_ _04063_ VGND VGND VPWR VPWR _04064_ sky130_fd_sc_hd__or2_1
X_10255_ _05556_ net539 _09186_ VGND VGND VPWR VPWR _00194_ sky130_fd_sc_hd__a21o_1
X_13043_ _02975_ _02980_ _02981_ VGND VGND VPWR VPWR _02982_ sky130_fd_sc_hd__a21oi_1
X_17920_ _08227_ _08225_ VGND VGND VPWR VPWR _08270_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17851_ net307 _07568_ VGND VGND VPWR VPWR _08194_ sky130_fd_sc_hd__nand2_1
X_10186_ _09362_ _09384_ VGND VGND VPWR VPWR _09395_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16802_ _07037_ _07039_ VGND VGND VPWR VPWR _07040_ sky130_fd_sc_hd__or2b_1
X_17782_ _08116_ _08115_ _08099_ _08082_ VGND VGND VPWR VPWR _08118_ sky130_fd_sc_hd__o211a_1
X_14994_ _05016_ _05012_ VGND VGND VPWR VPWR _05052_ sky130_fd_sc_hd__or2b_1
Xfanout290 ki\[12\] VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__clkbuf_4
X_16733_ net293 _06438_ _06962_ _06963_ VGND VGND VPWR VPWR _06965_ sky130_fd_sc_hd__a31o_1
X_13945_ net481 net117 VGND VGND VPWR VPWR _03917_ sky130_fd_sc_hd__nand2_2
XFILLER_0_88_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16664_ _02328_ _06285_ VGND VGND VPWR VPWR _06889_ sky130_fd_sc_hd__xor2_4
X_13876_ _03719_ _03750_ VGND VGND VPWR VPWR _03842_ sky130_fd_sc_hd__xnor2_1
X_15615_ _05725_ _05726_ _05717_ VGND VGND VPWR VPWR _05735_ sky130_fd_sc_hd__a21o_1
X_18403_ _06149_ _06152_ VGND VGND VPWR VPWR _08802_ sky130_fd_sc_hd__and2_1
X_12827_ _02660_ _02732_ _02733_ _02765_ VGND VGND VPWR VPWR _02766_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_9_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16595_ net272 _06724_ VGND VGND VPWR VPWR _06813_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18334_ _08715_ _08725_ VGND VGND VPWR VPWR _08726_ sky130_fd_sc_hd__xnor2_1
X_15546_ _05651_ _05657_ _05582_ _05658_ VGND VGND VPWR VPWR _05659_ sky130_fd_sc_hd__a211o_1
X_12758_ _02696_ VGND VGND VPWR VPWR _02697_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11709_ _01606_ _01613_ _01632_ _01647_ VGND VGND VPWR VPWR _01648_ sky130_fd_sc_hd__o31a_1
X_18265_ _08648_ _08649_ VGND VGND VPWR VPWR _08650_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15477_ _05582_ VGND VGND VPWR VPWR _05583_ sky130_fd_sc_hd__inv_2
X_12689_ _02576_ _02607_ _02627_ VGND VGND VPWR VPWR _02628_ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17216_ _07489_ _07495_ VGND VGND VPWR VPWR _07496_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14428_ _04428_ VGND VGND VPWR VPWR _04429_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18196_ _08572_ _08494_ _08573_ VGND VGND VPWR VPWR _08574_ sky130_fd_sc_hd__nand3_1
X_17147_ _07409_ _07419_ VGND VGND VPWR VPWR _07420_ sky130_fd_sc_hd__xor2_2
X_14359_ _04351_ _04352_ net407 net170 VGND VGND VPWR VPWR _04353_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_40_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout9 net404 VGND VGND VPWR VPWR net564 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17078_ _07332_ _07333_ _07343_ VGND VGND VPWR VPWR _07344_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16029_ _06179_ _06189_ VGND VGND VPWR VPWR _06190_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_9_Left_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10040_ _05589_ _05677_ _05556_ VGND VGND VPWR VPWR _07789_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold43 i_error\[15\] VGND VGND VPWR VPWR net550 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 i_error\[4\] VGND VGND VPWR VPWR net561 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11991_ _01779_ VGND VGND VPWR VPWR _01930_ sky130_fd_sc_hd__buf_2
X_13730_ _03691_ _03694_ VGND VGND VPWR VPWR _03696_ sky130_fd_sc_hd__or2_1
X_10942_ net371 _08207_ _00879_ _00880_ VGND VGND VPWR VPWR _00881_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_79_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13661_ net240 _02913_ _02745_ net243 VGND VGND VPWR VPWR _03623_ sky130_fd_sc_hd__a22o_1
X_10873_ _00811_ VGND VGND VPWR VPWR _00812_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_156_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15400_ _05495_ _05496_ _05497_ VGND VGND VPWR VPWR _05498_ sky130_fd_sc_hd__o21ba_1
X_12612_ _02534_ _02537_ _02539_ VGND VGND VPWR VPWR _02551_ sky130_fd_sc_hd__or3_1
XFILLER_0_39_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16380_ _06574_ _06575_ VGND VGND VPWR VPWR _06576_ sky130_fd_sc_hd__nor2_1
X_13592_ _03549_ _03550_ VGND VGND VPWR VPWR _03551_ sky130_fd_sc_hd__nor2_1
X_15331_ _05420_ _05421_ net437 net193 VGND VGND VPWR VPWR _05422_ sky130_fd_sc_hd__and4bb_1
X_12543_ _02480_ _02481_ VGND VGND VPWR VPWR _02482_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18050_ _08411_ _08412_ _08348_ _08373_ VGND VGND VPWR VPWR _08413_ sky130_fd_sc_hd__or4_1
X_15262_ net423 net197 VGND VGND VPWR VPWR _05346_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12474_ _02325_ _02404_ _02412_ VGND VGND VPWR VPWR _02413_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17001_ _07186_ _07258_ VGND VGND VPWR VPWR _07259_ sky130_fd_sc_hd__nor2_1
X_14213_ net422 net119 _04190_ VGND VGND VPWR VPWR _04193_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11425_ _01360_ _01363_ VGND VGND VPWR VPWR _01364_ sky130_fd_sc_hd__xor2_2
X_15193_ _05268_ _05269_ VGND VGND VPWR VPWR _05271_ sky130_fd_sc_hd__or2_1
XANTENNA_7 net540 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14144_ _04114_ _04116_ VGND VGND VPWR VPWR _04117_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11356_ _01290_ _01294_ VGND VGND VPWR VPWR _01295_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10307_ net342 _09583_ _09540_ VGND VGND VPWR VPWR _00246_ sky130_fd_sc_hd__a21o_1
X_14075_ _03937_ _03952_ VGND VGND VPWR VPWR _04047_ sky130_fd_sc_hd__or2b_1
X_18952_ _09270_ _09404_ VGND VGND VPWR VPWR _09405_ sky130_fd_sc_hd__xnor2_1
X_11287_ _01220_ _01225_ VGND VGND VPWR VPWR _01226_ sky130_fd_sc_hd__and2_1
X_13026_ _02961_ _02963_ _02964_ VGND VGND VPWR VPWR _02965_ sky130_fd_sc_hd__nand3_2
X_17903_ _08248_ _08250_ VGND VGND VPWR VPWR _08252_ sky130_fd_sc_hd__xnor2_1
X_10238_ _00174_ _00176_ VGND VGND VPWR VPWR _00177_ sky130_fd_sc_hd__and2b_1
X_18883_ _09280_ _09328_ VGND VGND VPWR VPWR _09330_ sky130_fd_sc_hd__xnor2_1
X_10169_ _05545_ _09153_ VGND VGND VPWR VPWR _09208_ sky130_fd_sc_hd__xnor2_1
X_17834_ _08175_ _08060_ VGND VGND VPWR VPWR _08176_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14977_ _05020_ _05026_ _05032_ VGND VGND VPWR VPWR _05033_ sky130_fd_sc_hd__nand3_1
X_17765_ _08072_ _08074_ VGND VGND VPWR VPWR _08100_ sky130_fd_sc_hd__or2_1
Xrebuffer19 _09203_ VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13928_ net451 net456 net116 VGND VGND VPWR VPWR _03898_ sky130_fd_sc_hd__o21ai_1
X_16716_ _06845_ _06945_ VGND VGND VPWR VPWR _06946_ sky130_fd_sc_hd__xnor2_1
X_17696_ _08022_ _08023_ VGND VGND VPWR VPWR _08024_ sky130_fd_sc_hd__or2b_1
X_16647_ _06867_ _06869_ VGND VGND VPWR VPWR _06870_ sky130_fd_sc_hd__nor2_1
X_13859_ _03818_ _03824_ VGND VGND VPWR VPWR _03825_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16578_ _06734_ _06793_ VGND VGND VPWR VPWR _06794_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15529_ _05552_ _05639_ VGND VGND VPWR VPWR _05640_ sky130_fd_sc_hd__nor2_1
X_18317_ _08690_ _08706_ VGND VGND VPWR VPWR _08707_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19297_ clknet_4_8_0_clock _00055_ VGND VGND VPWR VPWR ki\[8\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_155_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18248_ net273 _06346_ _06517_ _06516_ VGND VGND VPWR VPWR _08631_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18179_ net570 _08434_ _08553_ _08049_ VGND VGND VPWR VPWR _08555_ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09952_ net353 _04896_ _05006_ net357 VGND VGND VPWR VPWR _06821_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09883_ _06051_ VGND VGND VPWR VPWR _06062_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_73_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11210_ _01143_ _01139_ VGND VGND VPWR VPWR _01149_ sky130_fd_sc_hd__xnor2_1
X_12190_ net206 _01810_ VGND VGND VPWR VPWR _02129_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11141_ _00975_ _00987_ _00986_ VGND VGND VPWR VPWR _01080_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11072_ _00998_ _01010_ VGND VGND VPWR VPWR _01011_ sky130_fd_sc_hd__xor2_1
XFILLER_0_37_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput88 net88 VGND VGND VPWR VPWR out_clocked[17] sky130_fd_sc_hd__clkbuf_4
X_10023_ _06447_ _06766_ VGND VGND VPWR VPWR _07602_ sky130_fd_sc_hd__nand2_1
X_14900_ _04016_ net194 VGND VGND VPWR VPWR _04948_ sky130_fd_sc_hd__nor2_1
X_15880_ _05995_ _06025_ VGND VGND VPWR VPWR _06026_ sky130_fd_sc_hd__nor2_1
X_14831_ _04864_ _04867_ VGND VGND VPWR VPWR _04872_ sky130_fd_sc_hd__xor2_1
XFILLER_0_99_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17550_ _07832_ _07835_ VGND VGND VPWR VPWR _07863_ sky130_fd_sc_hd__xnor2_1
X_14762_ net470 net135 net130 net475 VGND VGND VPWR VPWR _04796_ sky130_fd_sc_hd__a22o_1
X_11974_ net205 _01854_ _01912_ VGND VGND VPWR VPWR _01913_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_98_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16501_ _06707_ _06708_ VGND VGND VPWR VPWR _06709_ sky130_fd_sc_hd__and2_1
X_13713_ _03673_ _03676_ _03678_ VGND VGND VPWR VPWR _03679_ sky130_fd_sc_hd__o21a_1
X_10925_ _00760_ _00863_ VGND VGND VPWR VPWR _00864_ sky130_fd_sc_hd__or2_2
X_17481_ _07740_ _07742_ _07744_ VGND VGND VPWR VPWR _07787_ sky130_fd_sc_hd__a21oi_1
X_14693_ _04681_ _04719_ VGND VGND VPWR VPWR _04721_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16432_ _06474_ _06472_ VGND VGND VPWR VPWR _06633_ sky130_fd_sc_hd__or2_1
X_19220_ clknet_4_4_0_clock _00102_ VGND VGND VPWR VPWR prev_error\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13644_ _03602_ _03604_ VGND VGND VPWR VPWR _03605_ sky130_fd_sc_hd__or2_1
X_10856_ _00700_ _00794_ VGND VGND VPWR VPWR _00795_ sky130_fd_sc_hd__xor2_4
XFILLER_0_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19151_ net505 net560 net495 _09569_ VGND VGND VPWR VPWR _00130_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16363_ _06555_ _06556_ VGND VGND VPWR VPWR _06558_ sky130_fd_sc_hd__or2_1
X_13575_ _03529_ _03533_ VGND VGND VPWR VPWR _03534_ sky130_fd_sc_hd__xor2_1
XFILLER_0_66_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10787_ _00642_ _00636_ _00641_ VGND VGND VPWR VPWR _00726_ sky130_fd_sc_hd__and3_1
XFILLER_0_143_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18102_ _08467_ _08468_ _08457_ _08469_ VGND VGND VPWR VPWR _08470_ sky130_fd_sc_hd__o211ai_2
X_15314_ _05318_ _05403_ VGND VGND VPWR VPWR _05404_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12526_ _02356_ _02463_ VGND VGND VPWR VPWR _02465_ sky130_fd_sc_hd__nor2_1
X_19082_ _09523_ _00615_ _09526_ net487 VGND VGND VPWR VPWR _00097_ sky130_fd_sc_hd__o211a_1
X_16294_ _06462_ _06478_ _06481_ VGND VGND VPWR VPWR _06482_ sky130_fd_sc_hd__o21a_1
XFILLER_0_26_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18033_ net326 net540 VGND VGND VPWR VPWR _08395_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15245_ net454 net172 net167 net459 VGND VGND VPWR VPWR _05328_ sky130_fd_sc_hd__a22oi_1
X_12457_ _02377_ _02392_ _02394_ VGND VGND VPWR VPWR _02396_ sky130_fd_sc_hd__or3_1
XFILLER_0_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11408_ _01312_ _01346_ VGND VGND VPWR VPWR _01347_ sky130_fd_sc_hd__or2_1
X_15176_ _05250_ _05251_ VGND VGND VPWR VPWR _05252_ sky130_fd_sc_hd__and2_1
X_12388_ _01726_ VGND VGND VPWR VPWR _02327_ sky130_fd_sc_hd__inv_2
X_14127_ _03988_ net113 _04095_ _04096_ VGND VGND VPWR VPWR _04099_ sky130_fd_sc_hd__o211ai_1
X_11339_ _01244_ _01276_ _01277_ VGND VGND VPWR VPWR _01278_ sky130_fd_sc_hd__a21bo_2
X_14058_ _03931_ _03933_ _04028_ VGND VGND VPWR VPWR _04030_ sky130_fd_sc_hd__or3_1
X_18935_ _09385_ _09386_ VGND VGND VPWR VPWR _09387_ sky130_fd_sc_hd__and2_1
X_13009_ net256 _01834_ VGND VGND VPWR VPWR _02948_ sky130_fd_sc_hd__nand2_2
X_18866_ _09310_ VGND VGND VPWR VPWR _09311_ sky130_fd_sc_hd__buf_1
X_17817_ _08154_ _08155_ _08148_ _08149_ VGND VGND VPWR VPWR _08157_ sky130_fd_sc_hd__o211ai_4
X_18797_ _09233_ _09234_ VGND VGND VPWR VPWR _09235_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17748_ _08076_ _08080_ VGND VGND VPWR VPWR _08081_ sky130_fd_sc_hd__xnor2_2
X_17679_ _08004_ _07911_ VGND VGND VPWR VPWR _08005_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_147_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_99_Left_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09935_ _06623_ VGND VGND VPWR VPWR _06634_ sky130_fd_sc_hd__buf_2
X_09866_ _05479_ _05853_ _05864_ VGND VGND VPWR VPWR _05875_ sky130_fd_sc_hd__a21o_1
X_09797_ _04907_ _05105_ VGND VGND VPWR VPWR _05116_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_9_0_clock clknet_0_clock VGND VGND VPWR VPWR clknet_4_9_0_clock sky130_fd_sc_hd__clkbuf_8
X_10710_ _00629_ _00647_ _00648_ VGND VGND VPWR VPWR _00649_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_49_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11690_ _01626_ _01628_ VGND VGND VPWR VPWR _01629_ sky130_fd_sc_hd__and2b_1
XFILLER_0_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10641_ _00577_ _00578_ VGND VGND VPWR VPWR _00580_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13360_ _03307_ _03310_ _03312_ VGND VGND VPWR VPWR _03313_ sky130_fd_sc_hd__o21a_1
X_10572_ _00510_ VGND VGND VPWR VPWR _00511_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12311_ _02246_ _02249_ VGND VGND VPWR VPWR _02250_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13291_ _03242_ _03243_ VGND VGND VPWR VPWR _03244_ sky130_fd_sc_hd__and2b_1
X_15030_ _05064_ _05090_ VGND VGND VPWR VPWR _05091_ sky130_fd_sc_hd__nand2_1
X_12242_ _01768_ _02180_ VGND VGND VPWR VPWR _02181_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12173_ _02073_ _02111_ VGND VGND VPWR VPWR _02112_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11124_ net370 _00244_ VGND VGND VPWR VPWR _01063_ sky130_fd_sc_hd__nand2_1
X_16981_ _07235_ _07194_ _07198_ VGND VGND VPWR VPWR _07237_ sky130_fd_sc_hd__or3_1
X_18720_ _09148_ _09149_ VGND VGND VPWR VPWR _09150_ sky130_fd_sc_hd__or2b_1
X_15932_ _05946_ _03851_ _06081_ _06082_ VGND VGND VPWR VPWR _06083_ sky130_fd_sc_hd__or4_1
X_11055_ _00802_ _00892_ VGND VGND VPWR VPWR _00994_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10006_ _07393_ _07404_ VGND VGND VPWR VPWR _07415_ sky130_fd_sc_hd__or2_1
X_15863_ _03891_ _06006_ VGND VGND VPWR VPWR _06008_ sky130_fd_sc_hd__xor2_1
X_18651_ _06108_ _09073_ VGND VGND VPWR VPWR _09074_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14814_ _04791_ _04853_ VGND VGND VPWR VPWR _04854_ sky130_fd_sc_hd__nor2_1
X_17602_ _07905_ _07919_ VGND VGND VPWR VPWR _07920_ sky130_fd_sc_hd__nand2b_1
X_15794_ _05782_ _05823_ _05889_ VGND VGND VPWR VPWR _05932_ sky130_fd_sc_hd__o21ai_1
X_18582_ _08994_ _08997_ VGND VGND VPWR VPWR _08998_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14745_ _04658_ _04660_ VGND VGND VPWR VPWR _04778_ sky130_fd_sc_hd__and2_1
X_17533_ net328 _06437_ _07842_ _07843_ VGND VGND VPWR VPWR _07845_ sky130_fd_sc_hd__a31o_1
XFILLER_0_157_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11957_ _01878_ _01868_ VGND VGND VPWR VPWR _01896_ sky130_fd_sc_hd__xor2_1
XFILLER_0_98_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17464_ _07711_ _07730_ VGND VGND VPWR VPWR _07769_ sky130_fd_sc_hd__nor2_1
X_10908_ _00728_ _00846_ VGND VGND VPWR VPWR _00847_ sky130_fd_sc_hd__xnor2_2
X_14676_ net458 net139 VGND VGND VPWR VPWR _04702_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11888_ _01800_ _01826_ VGND VGND VPWR VPWR _01827_ sky130_fd_sc_hd__nor2_1
X_19203_ clknet_4_12_0_clock _00085_ VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16415_ _06614_ _06484_ VGND VGND VPWR VPWR _06615_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_13_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13627_ _03585_ VGND VGND VPWR VPWR _03586_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10839_ _00777_ _00687_ VGND VGND VPWR VPWR _00778_ sky130_fd_sc_hd__xor2_1
X_17395_ _07632_ VGND VGND VPWR VPWR _07693_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19134_ net503 i_error\[8\] VGND VGND VPWR VPWR _09560_ sky130_fd_sc_hd__or2_1
X_16346_ net319 VGND VGND VPWR VPWR _06539_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13558_ _03453_ _03516_ VGND VGND VPWR VPWR _03517_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_132_Right_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12509_ _02391_ _02390_ VGND VGND VPWR VPWR _02448_ sky130_fd_sc_hd__and2b_1
X_19065_ _09515_ _09516_ VGND VGND VPWR VPWR _00089_ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16277_ _06432_ _06433_ VGND VGND VPWR VPWR _06463_ sky130_fd_sc_hd__nand2_2
X_13489_ net229 _02914_ _02746_ net232 VGND VGND VPWR VPWR _03448_ sky130_fd_sc_hd__a22o_1
X_15228_ _05304_ _05306_ _05308_ VGND VGND VPWR VPWR _05309_ sky130_fd_sc_hd__o21ai_1
X_18016_ _08352_ _08375_ VGND VGND VPWR VPWR _08376_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15159_ _05232_ _05130_ VGND VGND VPWR VPWR _05233_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout119 net120 VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__buf_2
X_09720_ _04236_ _04247_ _04258_ VGND VGND VPWR VPWR _04269_ sky130_fd_sc_hd__a21oi_4
X_18918_ _09283_ _09302_ _09304_ VGND VGND VPWR VPWR _09368_ sky130_fd_sc_hd__a21oi_1
X_09651_ net46 _03347_ _03380_ net206 VGND VGND VPWR VPWR _00006_ sky130_fd_sc_hd__a22o_1
X_18849_ _09288_ _09291_ VGND VGND VPWR VPWR _09292_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09918_ _05875_ _06436_ VGND VGND VPWR VPWR _06447_ sky130_fd_sc_hd__xnor2_1
X_09849_ _04907_ _05094_ _05677_ _05083_ VGND VGND VPWR VPWR _05688_ sky130_fd_sc_hd__a2bb2o_1
X_12860_ net247 _01860_ VGND VGND VPWR VPWR _02799_ sky130_fd_sc_hd__nand2_2
XFILLER_0_69_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11811_ _01703_ _01748_ _01749_ VGND VGND VPWR VPWR _01750_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_96_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12791_ _02711_ _02728_ _02729_ VGND VGND VPWR VPWR _02730_ sky130_fd_sc_hd__nand3_2
XFILLER_0_68_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14530_ net413 net175 net170 net417 VGND VGND VPWR VPWR _04541_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_96_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11742_ _01210_ _01281_ _01680_ VGND VGND VPWR VPWR _01681_ sky130_fd_sc_hd__and3_2
XFILLER_0_96_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14461_ _04437_ _04464_ VGND VGND VPWR VPWR _04465_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11673_ _01591_ _01608_ VGND VGND VPWR VPWR _01612_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16200_ _06325_ _06328_ _06377_ VGND VGND VPWR VPWR _06378_ sky130_fd_sc_hd__and3b_1
X_13412_ _03354_ _03365_ _03367_ VGND VGND VPWR VPWR _03368_ sky130_fd_sc_hd__o21a_2
X_17180_ _07430_ _07441_ VGND VGND VPWR VPWR _07456_ sky130_fd_sc_hd__nand2_1
X_10624_ _00561_ _00562_ VGND VGND VPWR VPWR _00563_ sky130_fd_sc_hd__and2_2
X_14392_ net461 net120 _03910_ VGND VGND VPWR VPWR _04389_ sky130_fd_sc_hd__and3_1
XFILLER_0_52_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16131_ prev_error\[12\] _06051_ _06301_ _01741_ VGND VGND VPWR VPWR _06302_ sky130_fd_sc_hd__a31o_1
X_13343_ _03292_ _03288_ VGND VGND VPWR VPWR _03296_ sky130_fd_sc_hd__and2b_1
X_10555_ _00402_ _00493_ VGND VGND VPWR VPWR _00494_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16062_ _08504_ _00184_ VGND VGND VPWR VPWR _06226_ sky130_fd_sc_hd__nand2_1
X_13274_ _03137_ _03226_ VGND VGND VPWR VPWR _03227_ sky130_fd_sc_hd__and2_1
X_10486_ _00396_ _00424_ VGND VGND VPWR VPWR _00425_ sky130_fd_sc_hd__or2_2
X_15013_ _04942_ _05071_ VGND VGND VPWR VPWR _05073_ sky130_fd_sc_hd__nor2_1
X_12225_ _01971_ _02008_ _02006_ VGND VGND VPWR VPWR _02164_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12156_ _02092_ _02094_ VGND VGND VPWR VPWR _02095_ sky130_fd_sc_hd__or2b_1
X_11107_ _00963_ _00965_ net402 _05314_ VGND VGND VPWR VPWR _01046_ sky130_fd_sc_hd__a2bb2o_1
X_12087_ _02021_ _02025_ VGND VGND VPWR VPWR _02026_ sky130_fd_sc_hd__and2_1
X_16964_ net317 _06345_ VGND VGND VPWR VPWR _07219_ sky130_fd_sc_hd__and2_1
X_18703_ _06146_ _09129_ _09130_ VGND VGND VPWR VPWR _09132_ sky130_fd_sc_hd__a21o_1
X_15915_ _06061_ _06064_ VGND VGND VPWR VPWR _06065_ sky130_fd_sc_hd__nand2_1
X_11038_ net383 _06183_ _00970_ _00976_ VGND VGND VPWR VPWR _00977_ sky130_fd_sc_hd__a31o_1
X_16895_ _07117_ _07141_ _07142_ VGND VGND VPWR VPWR _07143_ sky130_fd_sc_hd__a21o_1
X_18634_ _09046_ _09055_ VGND VGND VPWR VPWR _09056_ sky130_fd_sc_hd__or2_1
X_15846_ _05987_ _05988_ VGND VGND VPWR VPWR _05989_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18565_ _08973_ _08976_ _08979_ VGND VGND VPWR VPWR _08980_ sky130_fd_sc_hd__o21a_1
X_15777_ _05868_ _05905_ _05910_ _05912_ VGND VGND VPWR VPWR _05913_ sky130_fd_sc_hd__o31a_1
X_12989_ prev_error\[0\] _00809_ VGND VGND VPWR VPWR _02928_ sky130_fd_sc_hd__nand2_4
XFILLER_0_75_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17516_ _07557_ _07560_ VGND VGND VPWR VPWR _07826_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14728_ _04754_ _04756_ _04758_ VGND VGND VPWR VPWR _04759_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18496_ _08750_ net100 _08901_ _08902_ _08903_ VGND VGND VPWR VPWR _08904_ sky130_fd_sc_hd__a2111oi_4
XFILLER_0_157_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14659_ prev_d_error\[18\] net470 net131 VGND VGND VPWR VPWR _04683_ sky130_fd_sc_hd__and3_1
X_17447_ _07747_ _07749_ VGND VGND VPWR VPWR _07750_ sky130_fd_sc_hd__and2_1
XFILLER_0_157_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17378_ _07577_ _07599_ VGND VGND VPWR VPWR _07674_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19117_ net503 net548 net494 _09548_ VGND VGND VPWR VPWR _00114_ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16329_ _06511_ _06518_ VGND VGND VPWR VPWR _06520_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19048_ _04126_ net97 VGND VGND VPWR VPWR _09503_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09703_ net47 _03870_ _03903_ net340 VGND VGND VPWR VPWR _00064_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09634_ _03369_ VGND VGND VPWR VPWR _03380_ sky130_fd_sc_hd__buf_2
XFILLER_0_93_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10340_ net380 net520 _05149_ VGND VGND VPWR VPWR _00279_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10271_ net364 _05413_ _00209_ VGND VGND VPWR VPWR _00210_ sky130_fd_sc_hd__and3_1
X_12010_ _01947_ _01929_ VGND VGND VPWR VPWR _01949_ sky130_fd_sc_hd__and2b_1
Xfanout450 prev_d_error\[8\] VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__clkbuf_4
Xfanout461 net464 VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__buf_2
Xfanout472 prev_d_error\[3\] VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__buf_2
X_13961_ _03931_ _03932_ net421 net138 VGND VGND VPWR VPWR _03933_ sky130_fd_sc_hd__and4bb_1
Xfanout483 net484 VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__buf_2
XFILLER_0_45_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout494 net496 VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__clkbuf_4
X_15700_ _05819_ _05818_ VGND VGND VPWR VPWR _05828_ sky130_fd_sc_hd__or2b_1
X_12912_ net211 _02546_ _02750_ VGND VGND VPWR VPWR _02851_ sky130_fd_sc_hd__a21oi_1
X_16680_ _06857_ _06871_ VGND VGND VPWR VPWR _06906_ sky130_fd_sc_hd__and2_1
X_13892_ _03177_ _03179_ _03267_ VGND VGND VPWR VPWR _03858_ sky130_fd_sc_hd__a21o_1
X_15631_ _05749_ _05751_ VGND VGND VPWR VPWR _05752_ sky130_fd_sc_hd__nand2_1
X_12843_ _02778_ _02781_ VGND VGND VPWR VPWR _02782_ sky130_fd_sc_hd__xor2_2
XFILLER_0_57_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15562_ _05616_ _05668_ VGND VGND VPWR VPWR _05676_ sky130_fd_sc_hd__xnor2_1
X_18350_ _08742_ VGND VGND VPWR VPWR _08743_ sky130_fd_sc_hd__buf_4
X_12774_ _02706_ _02702_ VGND VGND VPWR VPWR _02713_ sky130_fd_sc_hd__or2b_1
XFILLER_0_56_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14513_ _04507_ _04521_ VGND VGND VPWR VPWR _04523_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17301_ net287 _07157_ VGND VGND VPWR VPWR _07589_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11725_ _01503_ _01579_ _01583_ _01584_ _01521_ VGND VGND VPWR VPWR _01664_ sky130_fd_sc_hd__a32oi_1
X_15493_ _05598_ _05599_ VGND VGND VPWR VPWR _05601_ sky130_fd_sc_hd__nor2_1
X_18281_ _08654_ _08666_ VGND VGND VPWR VPWR _08667_ sky130_fd_sc_hd__xor2_1
XFILLER_0_126_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14444_ net410 net170 _04351_ _04352_ VGND VGND VPWR VPWR _04447_ sky130_fd_sc_hd__o2bb2a_1
X_17232_ _07478_ _07479_ _07498_ VGND VGND VPWR VPWR _07513_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11656_ _01590_ _01594_ VGND VGND VPWR VPWR _01595_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17163_ _07086_ _07109_ VGND VGND VPWR VPWR _07438_ sky130_fd_sc_hd__xor2_1
XFILLER_0_142_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10607_ _00532_ _00544_ _00545_ VGND VGND VPWR VPWR _00546_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14375_ _04367_ _04369_ _04360_ _04364_ VGND VGND VPWR VPWR _04371_ sky130_fd_sc_hd__a211o_1
XFILLER_0_101_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11587_ _01492_ _01483_ _01491_ VGND VGND VPWR VPWR _01526_ sky130_fd_sc_hd__nand3_1
XFILLER_0_10_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16114_ _01724_ _00397_ VGND VGND VPWR VPWR _06284_ sky130_fd_sc_hd__nor2_1
X_13326_ net239 _02331_ VGND VGND VPWR VPWR _03279_ sky130_fd_sc_hd__nand2_1
X_17094_ _07359_ _07361_ VGND VGND VPWR VPWR _07362_ sky130_fd_sc_hd__xor2_2
XFILLER_0_134_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10538_ net379 _05292_ _05303_ VGND VGND VPWR VPWR _00477_ sky130_fd_sc_hd__and3_1
X_16045_ _07393_ _06207_ VGND VGND VPWR VPWR _06208_ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13257_ _03208_ _03209_ VGND VGND VPWR VPWR _03210_ sky130_fd_sc_hd__nand2_1
X_10469_ _00406_ _00407_ VGND VGND VPWR VPWR _00408_ sky130_fd_sc_hd__and2_2
X_12208_ _01996_ _02146_ VGND VGND VPWR VPWR _02147_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13188_ _03075_ _03140_ VGND VGND VPWR VPWR _03141_ sky130_fd_sc_hd__or2_1
X_12139_ _02076_ _02077_ VGND VGND VPWR VPWR _02078_ sky130_fd_sc_hd__nor2_1
X_17996_ net322 net318 _02931_ _07568_ VGND VGND VPWR VPWR _08354_ sky130_fd_sc_hd__and4_1
X_16947_ _07198_ _07199_ VGND VGND VPWR VPWR _07200_ sky130_fd_sc_hd__or2_2
X_16878_ _07014_ _07020_ VGND VGND VPWR VPWR _07124_ sky130_fd_sc_hd__xnor2_2
X_18617_ _08851_ VGND VGND VPWR VPWR _09037_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15829_ _04463_ _04465_ VGND VGND VPWR VPWR _05970_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18548_ _08885_ _08730_ _08891_ _08960_ VGND VGND VPWR VPWR _08961_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_59_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18479_ _06261_ net101 _06175_ VGND VGND VPWR VPWR _08885_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_118_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09617_ net55 _03102_ _03135_ net170 VGND VGND VPWR VPWR _00034_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11510_ _01420_ _01428_ _01430_ VGND VGND VPWR VPWR _01449_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12490_ net264 _01759_ VGND VGND VPWR VPWR _02429_ sky130_fd_sc_hd__nand2_2
XFILLER_0_34_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11441_ _01377_ _01379_ VGND VGND VPWR VPWR _01380_ sky130_fd_sc_hd__and2_1
XFILLER_0_151_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14160_ net422 net123 _04133_ VGND VGND VPWR VPWR _04134_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11372_ _01237_ _01106_ VGND VGND VPWR VPWR _01311_ sky130_fd_sc_hd__nor2_1
X_13111_ net220 net216 _02543_ _02639_ VGND VGND VPWR VPWR _03056_ sky130_fd_sc_hd__and4_1
XFILLER_0_61_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10323_ _00259_ _00261_ VGND VGND VPWR VPWR _00262_ sky130_fd_sc_hd__and2b_1
X_14091_ _04017_ net150 _04061_ VGND VGND VPWR VPWR _04063_ sky130_fd_sc_hd__o21ba_1
X_13042_ _02869_ _02867_ VGND VGND VPWR VPWR _02981_ sky130_fd_sc_hd__xor2_1
X_10254_ net372 _05182_ _00191_ _00192_ VGND VGND VPWR VPWR _00193_ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17850_ _08189_ _08192_ VGND VGND VPWR VPWR _08193_ sky130_fd_sc_hd__xnor2_1
X_10185_ _08317_ _09373_ VGND VGND VPWR VPWR _09384_ sky130_fd_sc_hd__or2_1
X_16801_ _06902_ _06974_ _06976_ _07038_ VGND VGND VPWR VPWR _07039_ sky130_fd_sc_hd__o31ai_2
X_17781_ _08082_ _08099_ _08115_ _08116_ VGND VGND VPWR VPWR _08117_ sky130_fd_sc_hd__a211oi_2
X_14993_ _05009_ _05011_ VGND VGND VPWR VPWR _05051_ sky130_fd_sc_hd__or2b_1
Xfanout280 ki\[15\] VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__clkbuf_4
Xfanout291 net292 VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__clkbuf_4
X_16732_ _06861_ _06960_ VGND VGND VPWR VPWR _06963_ sky130_fd_sc_hd__nor2_1
X_13944_ _03909_ _03915_ VGND VGND VPWR VPWR _03916_ sky130_fd_sc_hd__nor2b_4
XFILLER_0_89_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16663_ net278 net274 _06723_ _06803_ VGND VGND VPWR VPWR _06888_ sky130_fd_sc_hd__and4_1
X_13875_ _03837_ _03838_ _03839_ _03840_ VGND VGND VPWR VPWR _03841_ sky130_fd_sc_hd__a31o_1
X_18402_ _08799_ VGND VGND VPWR VPWR _08800_ sky130_fd_sc_hd__inv_2
X_15614_ _05728_ _05729_ _05725_ _05727_ VGND VGND VPWR VPWR _05734_ sky130_fd_sc_hd__o211a_1
X_12826_ _02759_ _02735_ VGND VGND VPWR VPWR _02765_ sky130_fd_sc_hd__or2b_1
X_16594_ net283 _06470_ _06811_ _06808_ VGND VGND VPWR VPWR _06812_ sky130_fd_sc_hd__a31o_1
X_18333_ _08717_ _08723_ VGND VGND VPWR VPWR _08725_ sky130_fd_sc_hd__xnor2_1
X_12757_ _02681_ _02695_ VGND VGND VPWR VPWR _02696_ sky130_fd_sc_hd__or2b_1
X_15545_ _05568_ _05581_ _05580_ VGND VGND VPWR VPWR _05658_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11708_ _01634_ _01646_ VGND VGND VPWR VPWR _01647_ sky130_fd_sc_hd__nand2_1
X_15476_ _05568_ _05580_ _05581_ VGND VGND VPWR VPWR _05582_ sky130_fd_sc_hd__and3_1
X_18264_ _08628_ _08629_ _08646_ VGND VGND VPWR VPWR _08649_ sky130_fd_sc_hd__nor3_1
X_12688_ _02625_ _02626_ VGND VGND VPWR VPWR _02627_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14427_ _04425_ _04426_ _04417_ _04421_ VGND VGND VPWR VPWR _04428_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_21_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17215_ _07491_ _07494_ VGND VGND VPWR VPWR _07495_ sky130_fd_sc_hd__nor2_1
X_11639_ _01547_ _01577_ VGND VGND VPWR VPWR _01578_ sky130_fd_sc_hd__nor2_1
X_18195_ _07974_ _08440_ _08491_ VGND VGND VPWR VPWR _08573_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17146_ _07410_ _07418_ VGND VGND VPWR VPWR _07419_ sky130_fd_sc_hd__xor2_2
X_14358_ net412 net165 net160 net416 VGND VGND VPWR VPWR _04352_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13309_ _03167_ _03170_ _03169_ VGND VGND VPWR VPWR _03262_ sky130_fd_sc_hd__a21o_1
XFILLER_0_122_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17077_ _07334_ _07342_ VGND VGND VPWR VPWR _07343_ sky130_fd_sc_hd__xor2_1
X_14289_ _04273_ _04275_ VGND VGND VPWR VPWR _04276_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16028_ _06187_ _06188_ VGND VGND VPWR VPWR _06189_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_71_Left_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17979_ _08332_ _08322_ _08334_ VGND VGND VPWR VPWR _08335_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_80_Left_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold44 i_error\[7\] VGND VGND VPWR VPWR net551 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ _01928_ VGND VGND VPWR VPWR _01929_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_97_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10941_ net379 net375 _06623_ _06172_ VGND VGND VPWR VPWR _00880_ sky130_fd_sc_hd__and4_1
X_13660_ _03620_ _03621_ VGND VGND VPWR VPWR _03622_ sky130_fd_sc_hd__nand2_1
X_10872_ _00810_ VGND VGND VPWR VPWR _00811_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_119_Left_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12611_ net202 _02546_ _02548_ _02549_ VGND VGND VPWR VPWR _02550_ sky130_fd_sc_hd__a31o_1
XFILLER_0_38_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13591_ _03458_ _03494_ VGND VGND VPWR VPWR _03550_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15330_ net441 net190 net184 net446 VGND VGND VPWR VPWR _05421_ sky130_fd_sc_hd__a22oi_1
X_12542_ _02265_ _02372_ _02371_ VGND VGND VPWR VPWR _02481_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15261_ _05343_ _05341_ VGND VGND VPWR VPWR _05345_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12473_ net206 _02224_ _02332_ net204 VGND VGND VPWR VPWR _02412_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17000_ net271 _07183_ _07185_ VGND VGND VPWR VPWR _07258_ sky130_fd_sc_hd__a21oi_1
X_14212_ net422 net119 _04190_ VGND VGND VPWR VPWR _04191_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11424_ _01361_ _01362_ VGND VGND VPWR VPWR _01363_ sky130_fd_sc_hd__nor2_1
X_15192_ _05256_ _05258_ _05267_ VGND VGND VPWR VPWR _05269_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_8 kd_1\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14143_ _04049_ _04051_ _04113_ VGND VGND VPWR VPWR _04116_ sky130_fd_sc_hd__or3_1
X_11355_ _01291_ _01292_ _01293_ VGND VGND VPWR VPWR _01294_ sky130_fd_sc_hd__a21boi_1
XPHY_EDGE_ROW_128_Left_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10306_ _00244_ VGND VGND VPWR VPWR _00245_ sky130_fd_sc_hd__buf_2
X_18951_ net422 net117 _04189_ _04131_ VGND VGND VPWR VPWR _09404_ sky130_fd_sc_hd__a31o_1
X_14074_ _04023_ _04037_ VGND VGND VPWR VPWR _04046_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11286_ _01217_ _01219_ VGND VGND VPWR VPWR _01225_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13025_ _02960_ _02955_ _02959_ VGND VGND VPWR VPWR _02964_ sky130_fd_sc_hd__nand3_1
X_17902_ _08194_ _08249_ VGND VGND VPWR VPWR _08250_ sky130_fd_sc_hd__nor2_1
X_10237_ _08427_ _00175_ VGND VGND VPWR VPWR _00176_ sky130_fd_sc_hd__nor2_1
X_18882_ _09326_ _09327_ VGND VGND VPWR VPWR _09328_ sky130_fd_sc_hd__nor2_1
X_17833_ net326 _06801_ VGND VGND VPWR VPWR _08175_ sky130_fd_sc_hd__nand2_1
X_10168_ _09175_ _09186_ _05556_ _05006_ VGND VGND VPWR VPWR _09197_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_83_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17764_ _08083_ _08098_ VGND VGND VPWR VPWR _08099_ sky130_fd_sc_hd__or2_1
X_10099_ _07767_ _08064_ _08427_ VGND VGND VPWR VPWR _08438_ sky130_fd_sc_hd__a21oi_1
X_14976_ _05029_ _05031_ VGND VGND VPWR VPWR _05032_ sky130_fd_sc_hd__nand2_1
X_16715_ _06848_ _06846_ VGND VGND VPWR VPWR _06945_ sky130_fd_sc_hd__nor2_1
X_13927_ net451 net456 net116 VGND VGND VPWR VPWR _03897_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_137_Left_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17695_ _08016_ _08021_ VGND VGND VPWR VPWR _08023_ sky130_fd_sc_hd__xor2_1
XFILLER_0_107_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16646_ _06868_ _06811_ VGND VGND VPWR VPWR _06869_ sky130_fd_sc_hd__xor2_1
X_13858_ _03817_ _03813_ _03815_ VGND VGND VPWR VPWR _03824_ sky130_fd_sc_hd__nor3_1
XFILLER_0_147_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12809_ _02640_ VGND VGND VPWR VPWR _02748_ sky130_fd_sc_hd__inv_2
X_16577_ _06399_ _06621_ _06732_ VGND VGND VPWR VPWR _06793_ sky130_fd_sc_hd__o21ba_1
X_13789_ _03753_ _03754_ VGND VGND VPWR VPWR _03755_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18316_ _08698_ _08705_ VGND VGND VPWR VPWR _08706_ sky130_fd_sc_hd__xnor2_1
X_15528_ net479 net164 _05550_ _05551_ VGND VGND VPWR VPWR _05639_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_127_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19296_ clknet_4_8_0_clock _00054_ VGND VGND VPWR VPWR ki\[7\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_143_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18247_ _06399_ _06346_ VGND VGND VPWR VPWR _08630_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15459_ _05555_ _05562_ VGND VGND VPWR VPWR _05563_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18178_ _08049_ _08553_ _08434_ _08432_ VGND VGND VPWR VPWR _08554_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_40_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17129_ _07373_ _07394_ _07399_ VGND VGND VPWR VPWR _07400_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09951_ _05688_ _06799_ _05820_ VGND VGND VPWR VPWR _06810_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_111_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09882_ _06040_ VGND VGND VPWR VPWR _06051_ sky130_fd_sc_hd__buf_4
XFILLER_0_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_146_Right_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11140_ _00975_ _00986_ _00987_ VGND VGND VPWR VPWR _01079_ sky130_fd_sc_hd__and3_1
Xclkbuf_4_5_0_clock clknet_0_clock VGND VGND VPWR VPWR clknet_4_5_0_clock sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11071_ _01000_ _01005_ _01009_ VGND VGND VPWR VPWR _01010_ sky130_fd_sc_hd__a21boi_1
Xoutput89 net89 VGND VGND VPWR VPWR out_clocked[18] sky130_fd_sc_hd__clkbuf_4
X_10022_ _07250_ _07580_ VGND VGND VPWR VPWR _07591_ sky130_fd_sc_hd__xnor2_1
X_14830_ net414 net190 _04869_ _04870_ VGND VGND VPWR VPWR _04871_ sky130_fd_sc_hd__a31o_1
XFILLER_0_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14761_ net470 net475 net134 net130 VGND VGND VPWR VPWR _04795_ sky130_fd_sc_hd__and4_1
X_11973_ net203 _01875_ VGND VGND VPWR VPWR _01912_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16500_ _06682_ _06704_ _06706_ VGND VGND VPWR VPWR _06708_ sky130_fd_sc_hd__nand3_1
X_13712_ _03641_ _03677_ VGND VGND VPWR VPWR _03678_ sky130_fd_sc_hd__nor2_1
X_10924_ _00761_ _00858_ _00862_ VGND VGND VPWR VPWR _00863_ sky130_fd_sc_hd__o21a_1
X_14692_ _04700_ _04718_ VGND VGND VPWR VPWR _04719_ sky130_fd_sc_hd__and2_1
X_17480_ _07270_ _07785_ VGND VGND VPWR VPWR _07786_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_113_Right_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16431_ _06629_ _06631_ VGND VGND VPWR VPWR _06632_ sky130_fd_sc_hd__or2b_1
XFILLER_0_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13643_ _03545_ _03601_ _03596_ _03600_ VGND VGND VPWR VPWR _03604_ sky130_fd_sc_hd__a211oi_1
X_10855_ _00718_ _00717_ VGND VGND VPWR VPWR _00794_ sky130_fd_sc_hd__and2b_1
XFILLER_0_85_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19150_ net505 _08965_ VGND VGND VPWR VPWR _09569_ sky130_fd_sc_hd__nand2_1
X_13574_ net262 net258 _02223_ _02332_ _03532_ VGND VGND VPWR VPWR _03533_ sky130_fd_sc_hd__a41o_1
X_16362_ _06488_ _06504_ VGND VGND VPWR VPWR _06556_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10786_ _00672_ _00677_ VGND VGND VPWR VPWR _00725_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_26_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18101_ _08454_ _08455_ _08456_ VGND VGND VPWR VPWR _08469_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12525_ _02356_ _02463_ VGND VGND VPWR VPWR _02464_ sky130_fd_sc_hd__and2_1
X_15313_ _05315_ _05317_ VGND VGND VPWR VPWR _05403_ sky130_fd_sc_hd__or2_1
X_19081_ net498 prev_error\[2\] VGND VGND VPWR VPWR _09526_ sky130_fd_sc_hd__or2_1
X_16293_ _06444_ _06479_ VGND VGND VPWR VPWR _06481_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18032_ _08381_ _08392_ VGND VGND VPWR VPWR _08393_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12456_ _02377_ _02392_ _02394_ VGND VGND VPWR VPWR _02395_ sky130_fd_sc_hd__o21ai_1
X_15244_ net449 net177 VGND VGND VPWR VPWR _05327_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11407_ _01282_ _01344_ VGND VGND VPWR VPWR _01346_ sky130_fd_sc_hd__xnor2_4
X_15175_ _05246_ _05244_ VGND VGND VPWR VPWR _05251_ sky130_fd_sc_hd__xnor2_1
X_12387_ _01723_ _01725_ _01727_ VGND VGND VPWR VPWR _02326_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14126_ _04039_ VGND VGND VPWR VPWR _04098_ sky130_fd_sc_hd__inv_2
X_11338_ _01272_ _01275_ _01202_ _01245_ VGND VGND VPWR VPWR _01277_ sky130_fd_sc_hd__o211ai_2
X_14057_ _03931_ _03933_ _04028_ VGND VGND VPWR VPWR _04029_ sky130_fd_sc_hd__o21ai_1
X_18934_ _04017_ net132 net122 net411 VGND VGND VPWR VPWR _09386_ sky130_fd_sc_hd__o211ai_1
X_11269_ _01136_ _01206_ _01207_ VGND VGND VPWR VPWR _01208_ sky130_fd_sc_hd__a21oi_1
X_13008_ _02804_ _02805_ VGND VGND VPWR VPWR _02947_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_118_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18865_ _02148_ _09309_ VGND VGND VPWR VPWR _09310_ sky130_fd_sc_hd__or2_1
X_17816_ _08148_ _08149_ _08154_ _08155_ VGND VGND VPWR VPWR _08156_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_145_Left_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18796_ net412 net418 net126 net119 VGND VGND VPWR VPWR _09234_ sky130_fd_sc_hd__and4_1
X_17747_ _08077_ _08079_ VGND VGND VPWR VPWR _08080_ sky130_fd_sc_hd__xor2_2
X_14959_ net449 net163 VGND VGND VPWR VPWR _05013_ sky130_fd_sc_hd__nand2_1
X_17678_ net301 _07095_ VGND VGND VPWR VPWR _08004_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16629_ _06842_ _06841_ VGND VGND VPWR VPWR _06850_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_154_Left_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19279_ clknet_4_6_0_clock _00075_ VGND VGND VPWR VPWR kp\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09934_ _06612_ VGND VGND VPWR VPWR _06623_ sky130_fd_sc_hd__buf_2
X_09865_ _05666_ _05842_ VGND VGND VPWR VPWR _05864_ sky130_fd_sc_hd__nor2_1
X_09796_ _05006_ _05083_ _05094_ VGND VGND VPWR VPWR _05105_ sky130_fd_sc_hd__a21o_1
XFILLER_0_84_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10640_ _00577_ _00578_ VGND VGND VPWR VPWR _00579_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10571_ _00508_ _00509_ VGND VGND VPWR VPWR _00510_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12310_ _02248_ VGND VGND VPWR VPWR _02249_ sky130_fd_sc_hd__inv_2
X_13290_ _03236_ _03240_ VGND VGND VPWR VPWR _03243_ sky130_fd_sc_hd__xor2_2
XFILLER_0_90_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12241_ _02036_ _02179_ VGND VGND VPWR VPWR _02180_ sky130_fd_sc_hd__xor2_1
XFILLER_0_32_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12172_ _02073_ _02109_ _02110_ VGND VGND VPWR VPWR _02111_ sky130_fd_sc_hd__nor3_2
XFILLER_0_48_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11123_ _01045_ _01060_ VGND VGND VPWR VPWR _01062_ sky130_fd_sc_hd__xor2_4
X_16980_ _07194_ _07198_ _07235_ VGND VGND VPWR VPWR _07236_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15931_ _03609_ _03848_ _03850_ VGND VGND VPWR VPWR _06082_ sky130_fd_sc_hd__and3_1
X_11054_ _00985_ _00981_ VGND VGND VPWR VPWR _00993_ sky130_fd_sc_hd__and2b_1
X_10005_ _06810_ _06975_ VGND VGND VPWR VPWR _07404_ sky130_fd_sc_hd__xnor2_1
X_18650_ _06107_ _06060_ _06105_ VGND VGND VPWR VPWR _09073_ sky130_fd_sc_hd__nand3_1
X_15862_ _04158_ _06005_ VGND VGND VPWR VPWR _06006_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17601_ _07905_ _07906_ _07918_ VGND VGND VPWR VPWR _07919_ sky130_fd_sc_hd__or3_1
X_14813_ _04828_ _04851_ VGND VGND VPWR VPWR _04853_ sky130_fd_sc_hd__nor2_1
X_18581_ _06133_ _08993_ VGND VGND VPWR VPWR _08997_ sky130_fd_sc_hd__or2_1
X_15793_ _05929_ _05865_ VGND VGND VPWR VPWR _05931_ sky130_fd_sc_hd__or2b_1
X_17532_ net323 _06618_ _07480_ VGND VGND VPWR VPWR _07843_ sky130_fd_sc_hd__and3_1
X_14744_ _04773_ _04776_ VGND VGND VPWR VPWR _04777_ sky130_fd_sc_hd__nor2_1
X_11956_ _01848_ _01875_ VGND VGND VPWR VPWR _01895_ sky130_fd_sc_hd__or2_1
XFILLER_0_157_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17463_ _07732_ _07758_ VGND VGND VPWR VPWR _07768_ sky130_fd_sc_hd__nand2_1
X_10907_ _00731_ _00737_ VGND VGND VPWR VPWR _00846_ sky130_fd_sc_hd__xnor2_1
X_11887_ net221 _01810_ _01793_ _01794_ VGND VGND VPWR VPWR _01826_ sky130_fd_sc_hd__o2bb2a_1
X_14675_ net449 net148 VGND VGND VPWR VPWR _04701_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19202_ clknet_4_12_0_clock _00084_ VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dfxtp_1
X_16414_ _06399_ _06438_ VGND VGND VPWR VPWR _06614_ sky130_fd_sc_hd__or2_1
X_13626_ _03582_ _03584_ VGND VGND VPWR VPWR _03585_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10838_ net363 _08196_ VGND VGND VPWR VPWR _00777_ sky130_fd_sc_hd__nand2_1
X_17394_ _07655_ _07656_ _07691_ VGND VGND VPWR VPWR _07692_ sky130_fd_sc_hd__nor3_1
XFILLER_0_144_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19133_ _04137_ VGND VGND VPWR VPWR _09559_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16345_ net324 VGND VGND VPWR VPWR _06538_ sky130_fd_sc_hd__inv_2
X_13557_ net220 _03220_ _03452_ VGND VGND VPWR VPWR _03516_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10769_ _00618_ _00616_ VGND VGND VPWR VPWR _00708_ sky130_fd_sc_hd__and2b_1
XFILLER_0_81_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12508_ _02440_ _02445_ _02446_ VGND VGND VPWR VPWR _02447_ sky130_fd_sc_hd__o21ai_1
X_19064_ net505 net541 net495 VGND VGND VPWR VPWR _09516_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_113_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13488_ _03397_ _03446_ VGND VGND VPWR VPWR _03447_ sky130_fd_sc_hd__nor2_1
X_16276_ _06454_ _06459_ _06461_ VGND VGND VPWR VPWR _06462_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_152_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18015_ _08354_ _08353_ VGND VGND VPWR VPWR _08375_ sky130_fd_sc_hd__nor2_1
X_12439_ net221 _01861_ _02287_ VGND VGND VPWR VPWR _02378_ sky130_fd_sc_hd__a21oi_1
X_15227_ _05210_ _05307_ VGND VGND VPWR VPWR _05308_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15158_ _05131_ _05129_ VGND VGND VPWR VPWR _05232_ sky130_fd_sc_hd__nor2_1
X_14109_ _04080_ VGND VGND VPWR VPWR _04081_ sky130_fd_sc_hd__inv_2
X_15089_ _05045_ _05048_ VGND VGND VPWR VPWR _05156_ sky130_fd_sc_hd__nor2_1
X_18917_ _09366_ _09338_ _09335_ VGND VGND VPWR VPWR _09367_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09650_ net45 _03347_ _03380_ net210 VGND VGND VPWR VPWR _00005_ sky130_fd_sc_hd__a22o_1
X_18848_ _02129_ _09289_ _09290_ VGND VGND VPWR VPWR _09291_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_0_clock clock VGND VGND VPWR VPWR clknet_0_clock sky130_fd_sc_hd__clkbuf_16
X_18779_ _09214_ _09211_ VGND VGND VPWR VPWR _09215_ sky130_fd_sc_hd__or2_4
XFILLER_0_89_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09917_ _05941_ _06425_ VGND VGND VPWR VPWR _06436_ sky130_fd_sc_hd__xnor2_1
X_09848_ _05006_ VGND VGND VPWR VPWR _05677_ sky130_fd_sc_hd__buf_2
X_09779_ _04159_ _04797_ _04786_ _04808_ VGND VGND VPWR VPWR _04918_ sky130_fd_sc_hd__a31o_1
X_11810_ net520 _05149_ prev_error\[15\] VGND VGND VPWR VPWR _01749_ sky130_fd_sc_hd__a21bo_1
X_12790_ _02606_ _02710_ _02697_ _02709_ VGND VGND VPWR VPWR _02729_ sky130_fd_sc_hd__a211o_1
XFILLER_0_157_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11741_ _01350_ _01677_ _01678_ _01679_ _01280_ VGND VGND VPWR VPWR _01680_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_84_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14460_ _04436_ _04409_ _04433_ VGND VGND VPWR VPWR _04464_ sky130_fd_sc_hd__nand3_1
XFILLER_0_55_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11672_ _01587_ _01610_ VGND VGND VPWR VPWR _01611_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13411_ _03318_ _03366_ VGND VGND VPWR VPWR _03367_ sky130_fd_sc_hd__nor2_1
X_10623_ _00559_ _00560_ VGND VGND VPWR VPWR _00562_ sky130_fd_sc_hd__or2_1
X_14391_ _04386_ _04387_ net448 net133 VGND VGND VPWR VPWR _04388_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13342_ _03294_ _03222_ VGND VGND VPWR VPWR _03295_ sky130_fd_sc_hd__xnor2_1
X_16130_ prev_error\[13\] _05314_ VGND VGND VPWR VPWR _06301_ sky130_fd_sc_hd__or2_1
X_10554_ net350 _09583_ _00401_ VGND VGND VPWR VPWR _00493_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16061_ _06223_ _06224_ VGND VGND VPWR VPWR _06225_ sky130_fd_sc_hd__nor2_1
X_13273_ _03130_ _03133_ _03136_ VGND VGND VPWR VPWR _03226_ sky130_fd_sc_hd__nand3_1
XFILLER_0_122_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10485_ _00421_ _00423_ VGND VGND VPWR VPWR _00424_ sky130_fd_sc_hd__and2b_1
X_12224_ _02145_ _02162_ VGND VGND VPWR VPWR _02163_ sky130_fd_sc_hd__xnor2_1
X_15012_ net410 kd_2\[0\] _04939_ _05070_ VGND VGND VPWR VPWR _05071_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_60_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12155_ _02084_ _02093_ VGND VGND VPWR VPWR _02094_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11106_ _00968_ _00972_ VGND VGND VPWR VPWR _01045_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_75_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16963_ _07211_ _07216_ VGND VGND VPWR VPWR _07218_ sky130_fd_sc_hd__xor2_1
X_12086_ _02022_ _02024_ VGND VGND VPWR VPWR _02025_ sky130_fd_sc_hd__nand2_1
X_18702_ _08930_ _08964_ _09127_ _09124_ VGND VGND VPWR VPWR _09130_ sky130_fd_sc_hd__o211a_1
X_15914_ _03860_ _06063_ VGND VGND VPWR VPWR _06064_ sky130_fd_sc_hd__and2_1
X_11037_ net388 _05996_ _00567_ VGND VGND VPWR VPWR _00976_ sky130_fd_sc_hd__and3_1
X_16894_ _07138_ _07139_ VGND VGND VPWR VPWR _07142_ sky130_fd_sc_hd__nor2_1
X_18633_ _09048_ _09051_ _09053_ VGND VGND VPWR VPWR _09055_ sky130_fd_sc_hd__o21ba_1
X_15845_ _05986_ _05972_ _05983_ VGND VGND VPWR VPWR _05988_ sky130_fd_sc_hd__nor3_1
XFILLER_0_59_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18564_ _06131_ _08978_ VGND VGND VPWR VPWR _08979_ sky130_fd_sc_hd__nand2_1
X_15776_ _05889_ _05911_ VGND VGND VPWR VPWR _05912_ sky130_fd_sc_hd__nand2_1
X_12988_ _02924_ _02926_ VGND VGND VPWR VPWR _02927_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17515_ _07556_ _07821_ _07824_ VGND VGND VPWR VPWR _07825_ sky130_fd_sc_hd__o21ba_1
X_14727_ _04569_ _04757_ VGND VGND VPWR VPWR _04758_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11939_ _01869_ _01870_ _01877_ VGND VGND VPWR VPWR _01878_ sky130_fd_sc_hd__o21ai_1
X_18495_ _08899_ _08764_ VGND VGND VPWR VPWR _08903_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17446_ _07683_ _07748_ VGND VGND VPWR VPWR _07749_ sky130_fd_sc_hd__nand2_1
X_14658_ _04614_ _04616_ _03917_ VGND VGND VPWR VPWR _04682_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13609_ net243 net240 _02640_ _02746_ VGND VGND VPWR VPWR _03568_ sky130_fd_sc_hd__and4_1
XFILLER_0_28_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17377_ _07664_ _07672_ VGND VGND VPWR VPWR _07673_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14589_ _03913_ _04603_ _04605_ VGND VGND VPWR VPWR _04606_ sky130_fd_sc_hd__o21a_1
XFILLER_0_144_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19116_ net503 _09128_ VGND VGND VPWR VPWR _09548_ sky130_fd_sc_hd__nand2_1
X_16328_ _06511_ _06518_ VGND VGND VPWR VPWR _06519_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19047_ _09501_ _09502_ net492 VGND VGND VPWR VPWR _00083_ sky130_fd_sc_hd__o21a_1
XFILLER_0_152_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16259_ _06427_ _06429_ VGND VGND VPWR VPWR _06443_ sky130_fd_sc_hd__xor2_1
XFILLER_0_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09702_ net46 _03870_ _03903_ net343 VGND VGND VPWR VPWR _00063_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09633_ _03069_ _03336_ net487 VGND VGND VPWR VPWR _03369_ sky130_fd_sc_hd__o21a_1
XFILLER_0_65_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10270_ net368 _05292_ _05303_ VGND VGND VPWR VPWR _00209_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout440 net442 VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__clkbuf_4
Xfanout451 net452 VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__buf_2
Xfanout462 net464 VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__buf_2
Xfanout473 net474 VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__buf_2
X_13960_ net426 net133 net128 net567 VGND VGND VPWR VPWR _03932_ sky130_fd_sc_hd__a22oi_1
Xfanout484 net485 VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__buf_2
Xfanout495 net496 VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__clkbuf_4
X_12911_ net211 _02545_ _02750_ VGND VGND VPWR VPWR _02850_ sky130_fd_sc_hd__and3_1
X_13891_ _03423_ _03855_ _03856_ VGND VGND VPWR VPWR _03857_ sky130_fd_sc_hd__a21oi_2
X_15630_ _05744_ _05750_ VGND VGND VPWR VPWR _05751_ sky130_fd_sc_hd__and2_1
X_12842_ _02779_ _02780_ VGND VGND VPWR VPWR _02781_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_100_Left_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15561_ _05548_ _05674_ VGND VGND VPWR VPWR _05675_ sky130_fd_sc_hd__xor2_1
X_12773_ _02700_ _02701_ VGND VGND VPWR VPWR _02712_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17300_ _07586_ _07587_ VGND VGND VPWR VPWR _07588_ sky130_fd_sc_hd__xnor2_1
X_14512_ net435 net152 _04505_ _04506_ VGND VGND VPWR VPWR _04521_ sky130_fd_sc_hd__o2bb2a_1
X_11724_ _01508_ _01662_ VGND VGND VPWR VPWR _01663_ sky130_fd_sc_hd__nand2_1
X_18280_ _06555_ _08665_ VGND VGND VPWR VPWR _08666_ sky130_fd_sc_hd__xor2_1
X_15492_ _05593_ _05597_ VGND VGND VPWR VPWR _05599_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17231_ _07504_ _07511_ VGND VGND VPWR VPWR _07512_ sky130_fd_sc_hd__xnor2_1
X_14443_ _04443_ _04444_ net420 net161 VGND VGND VPWR VPWR _04446_ sky130_fd_sc_hd__and4bb_1
X_11655_ net381 _00810_ _01588_ _01589_ VGND VGND VPWR VPWR _01594_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17162_ _07396_ _07398_ _07400_ VGND VGND VPWR VPWR _07436_ sky130_fd_sc_hd__a21bo_1
X_10606_ _00533_ _00543_ VGND VGND VPWR VPWR _00545_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14374_ _04360_ _04364_ _04367_ _04369_ VGND VGND VPWR VPWR _04370_ sky130_fd_sc_hd__o211ai_2
X_11586_ _01497_ _01524_ VGND VGND VPWR VPWR _01525_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16113_ _06274_ _06280_ _06281_ VGND VGND VPWR VPWR _06283_ sky130_fd_sc_hd__a21o_2
X_13325_ _03276_ _03277_ VGND VGND VPWR VPWR _03278_ sky130_fd_sc_hd__nand2_1
X_10537_ net375 _05314_ _05413_ net379 VGND VGND VPWR VPWR _00476_ sky130_fd_sc_hd__a22oi_1
X_17093_ _07058_ _07059_ VGND VGND VPWR VPWR _07361_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_10_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16044_ _06201_ _06206_ VGND VGND VPWR VPWR _06207_ sky130_fd_sc_hd__xnor2_1
X_13256_ net228 _02545_ _02409_ net232 VGND VGND VPWR VPWR _03209_ sky130_fd_sc_hd__a22o_1
X_10468_ _04280_ _00238_ _04335_ VGND VGND VPWR VPWR _00407_ sky130_fd_sc_hd__a21o_1
XFILLER_0_150_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12207_ kd_1\[11\] _01789_ VGND VGND VPWR VPWR _02146_ sky130_fd_sc_hd__nand2_1
X_13187_ _03073_ _03074_ VGND VGND VPWR VPWR _03140_ sky130_fd_sc_hd__nor2_1
X_10399_ _00336_ _00337_ VGND VGND VPWR VPWR _00338_ sky130_fd_sc_hd__nor2_1
X_12138_ net213 _01861_ _01835_ net217 VGND VGND VPWR VPWR _02077_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_19_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17995_ net318 _02931_ _07568_ net322 VGND VGND VPWR VPWR _08353_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_19_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16946_ net294 _06724_ _07197_ VGND VGND VPWR VPWR _07199_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12069_ _02006_ _02007_ VGND VGND VPWR VPWR _02008_ sky130_fd_sc_hd__nor2_1
X_16877_ _07120_ _07122_ VGND VGND VPWR VPWR _07123_ sky130_fd_sc_hd__nand2_1
X_18616_ _06113_ _09035_ VGND VGND VPWR VPWR _09036_ sky130_fd_sc_hd__xnor2_2
X_15828_ _04670_ _04671_ VGND VGND VPWR VPWR _05969_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18547_ _08954_ _08958_ _08959_ VGND VGND VPWR VPWR _08960_ sky130_fd_sc_hd__a21o_1
X_15759_ _05891_ _05892_ VGND VGND VPWR VPWR _05893_ sky130_fd_sc_hd__or2_1
X_18478_ _08883_ VGND VGND VPWR VPWR _08884_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17429_ _07711_ _07713_ _07729_ VGND VGND VPWR VPWR _07730_ sky130_fd_sc_hd__nor3_1
XFILLER_0_62_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09616_ net54 _03102_ _03135_ net175 VGND VGND VPWR VPWR _00033_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11440_ net400 _08185_ _01377_ _01378_ VGND VGND VPWR VPWR _01379_ sky130_fd_sc_hd__nand4_1
XFILLER_0_18_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11371_ _01300_ _01309_ VGND VGND VPWR VPWR _01310_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13110_ _02939_ _03054_ VGND VGND VPWR VPWR _03055_ sky130_fd_sc_hd__or2_1
X_10322_ _00223_ _00224_ _00260_ VGND VGND VPWR VPWR _00261_ sky130_fd_sc_hd__a21bo_2
X_14090_ net150 _04061_ prev_d_error\[18\] VGND VGND VPWR VPWR _04062_ sky130_fd_sc_hd__and3b_1
XFILLER_0_104_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13041_ _02977_ _02979_ VGND VGND VPWR VPWR _02980_ sky130_fd_sc_hd__nand2_1
X_10253_ net379 _04984_ _00190_ VGND VGND VPWR VPWR _00192_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10184_ net348 _06007_ _08306_ VGND VGND VPWR VPWR _09373_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16800_ _07005_ _06978_ VGND VGND VPWR VPWR _07038_ sky130_fd_sc_hd__or2b_1
X_17780_ _08104_ _08105_ _08114_ VGND VGND VPWR VPWR _08116_ sky130_fd_sc_hd__nor3_1
X_14992_ _05045_ _05048_ VGND VGND VPWR VPWR _05049_ sky130_fd_sc_hd__and2_1
Xfanout270 ki\[18\] VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__buf_4
Xfanout281 ki\[14\] VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__clkbuf_4
X_16731_ _06861_ _06960_ _06961_ VGND VGND VPWR VPWR _06962_ sky130_fd_sc_hd__o21a_1
Xfanout292 ki\[11\] VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__clkbuf_4
X_13943_ _03911_ _03913_ VGND VGND VPWR VPWR _03915_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_88_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16662_ _06884_ _06885_ VGND VGND VPWR VPWR _06886_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13874_ _03807_ _03808_ _03786_ VGND VGND VPWR VPWR _03840_ sky130_fd_sc_hd__o21a_1
X_18401_ _08798_ _08564_ VGND VGND VPWR VPWR _08799_ sky130_fd_sc_hd__xnor2_2
X_15613_ _05676_ _05731_ VGND VGND VPWR VPWR _05733_ sky130_fd_sc_hd__or2_1
X_12825_ _02678_ _02763_ VGND VGND VPWR VPWR _02764_ sky130_fd_sc_hd__xnor2_1
X_16593_ _06808_ _06809_ VGND VGND VPWR VPWR _06811_ sky130_fd_sc_hd__nor2_1
X_18332_ _08718_ _08722_ VGND VGND VPWR VPWR _08723_ sky130_fd_sc_hd__xnor2_1
X_15544_ _05652_ _05656_ VGND VGND VPWR VPWR _05657_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12756_ _02683_ _02688_ _02694_ VGND VGND VPWR VPWR _02695_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11707_ _01643_ _01644_ _01645_ VGND VGND VPWR VPWR _01646_ sky130_fd_sc_hd__and3b_1
X_18263_ _08628_ _08629_ _08646_ VGND VGND VPWR VPWR _08648_ sky130_fd_sc_hd__o21a_1
X_15475_ _05566_ _05555_ _05564_ VGND VGND VPWR VPWR _05581_ sky130_fd_sc_hd__nand3_1
X_12687_ _02576_ _02607_ VGND VGND VPWR VPWR _02626_ sky130_fd_sc_hd__xor2_1
XFILLER_0_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17214_ net332 _06344_ _07493_ VGND VGND VPWR VPWR _07494_ sky130_fd_sc_hd__a21boi_1
X_14426_ _04417_ _04421_ _04425_ _04426_ VGND VGND VPWR VPWR _04427_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_127_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11638_ _01573_ _01576_ VGND VGND VPWR VPWR _01577_ sky130_fd_sc_hd__and2b_1
X_18194_ _08484_ _08490_ VGND VGND VPWR VPWR _08572_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17145_ _07416_ _07417_ VGND VGND VPWR VPWR _07418_ sky130_fd_sc_hd__nor2_1
X_14357_ net412 net416 net165 net160 VGND VGND VPWR VPWR _04351_ sky130_fd_sc_hd__and4_1
X_11569_ _01479_ _01505_ VGND VGND VPWR VPWR _01508_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13308_ _03259_ _03260_ VGND VGND VPWR VPWR _03261_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17076_ _07335_ _07341_ VGND VGND VPWR VPWR _07342_ sky130_fd_sc_hd__xor2_1
X_14288_ _04272_ _04263_ _04270_ VGND VGND VPWR VPWR _04275_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16027_ _06186_ _06185_ VGND VGND VPWR VPWR _06188_ sky130_fd_sc_hd__and2b_1
X_13239_ _03101_ _03100_ VGND VGND VPWR VPWR _03192_ sky130_fd_sc_hd__and2b_1
XFILLER_0_122_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17978_ _08331_ _08333_ VGND VGND VPWR VPWR _08334_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_127_Right_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16929_ net274 _07157_ VGND VGND VPWR VPWR _07180_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold34 net84 VGND VGND VPWR VPWR net541 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 i_error\[6\] VGND VGND VPWR VPWR net552 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10940_ net375 _06623_ _06172_ net379 VGND VGND VPWR VPWR _00879_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10871_ _00809_ VGND VGND VPWR VPWR _00810_ sky130_fd_sc_hd__buf_2
Xclkbuf_4_1_0_clock clknet_0_clock VGND VGND VPWR VPWR clknet_4_1_0_clock sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12610_ _02404_ _02547_ VGND VGND VPWR VPWR _02549_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13590_ _03501_ _03548_ VGND VGND VPWR VPWR _03549_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12541_ net235 _01807_ VGND VGND VPWR VPWR _02480_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15260_ _05341_ _05343_ VGND VGND VPWR VPWR _05344_ sky130_fd_sc_hd__and2b_1
XFILLER_0_152_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12472_ net202 _02410_ VGND VGND VPWR VPWR _02411_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14211_ _04131_ _04189_ net117 VGND VGND VPWR VPWR _04190_ sky130_fd_sc_hd__and3b_1
X_11423_ _01293_ _01292_ _01291_ VGND VGND VPWR VPWR _01362_ sky130_fd_sc_hd__a21oi_1
X_15191_ _05256_ _05258_ _05267_ VGND VGND VPWR VPWR _05268_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_9 ki\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14142_ _04049_ _04051_ _04113_ VGND VGND VPWR VPWR _04114_ sky130_fd_sc_hd__o21ai_2
X_11354_ net377 net374 _00798_ _01001_ VGND VGND VPWR VPWR _01293_ sky130_fd_sc_hd__nand4_1
XFILLER_0_132_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10305_ _00243_ VGND VGND VPWR VPWR _00244_ sky130_fd_sc_hd__clkbuf_4
X_18950_ _09379_ _09402_ VGND VGND VPWR VPWR _09403_ sky130_fd_sc_hd__xnor2_1
X_14073_ _04041_ _04042_ _04044_ VGND VGND VPWR VPWR _04045_ sky130_fd_sc_hd__nor3_1
X_11285_ _01221_ _01222_ _01223_ VGND VGND VPWR VPWR _01224_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_120_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10236_ _08405_ _08416_ VGND VGND VPWR VPWR _00175_ sky130_fd_sc_hd__nor2_1
X_13024_ _02891_ _02962_ VGND VGND VPWR VPWR _02963_ sky130_fd_sc_hd__and2_1
X_17901_ net310 _02931_ VGND VGND VPWR VPWR _08249_ sky130_fd_sc_hd__nand2_1
X_18881_ _09324_ _09325_ VGND VGND VPWR VPWR _09327_ sky130_fd_sc_hd__and2_1
X_17832_ _08171_ _08172_ VGND VGND VPWR VPWR _08173_ sky130_fd_sc_hd__xor2_1
X_10167_ net380 _05072_ net539 net376 VGND VGND VPWR VPWR _09186_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_83_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17763_ _08089_ _08096_ VGND VGND VPWR VPWR _08098_ sky130_fd_sc_hd__xnor2_2
X_10098_ _08405_ _08416_ VGND VGND VPWR VPWR _08427_ sky130_fd_sc_hd__and2_1
X_14975_ _05030_ _05025_ VGND VGND VPWR VPWR _05031_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16714_ _06938_ _06941_ _06943_ VGND VGND VPWR VPWR _06944_ sky130_fd_sc_hd__o21ai_2
X_13926_ _03893_ _03894_ _03895_ VGND VGND VPWR VPWR _03896_ sky130_fd_sc_hd__o21ba_2
X_17694_ net290 _02933_ VGND VGND VPWR VPWR _08022_ sky130_fd_sc_hd__nand2_1
X_16645_ net283 _06470_ VGND VGND VPWR VPWR _06868_ sky130_fd_sc_hd__nand2_1
X_13857_ _03808_ _03822_ VGND VGND VPWR VPWR _03823_ sky130_fd_sc_hd__xnor2_1
X_12808_ _02746_ VGND VGND VPWR VPWR _02747_ sky130_fd_sc_hd__clkbuf_4
X_16576_ _06770_ _06782_ _06791_ VGND VGND VPWR VPWR _06792_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13788_ net251 _02913_ _02407_ net267 VGND VGND VPWR VPWR _03754_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18315_ _08699_ _08704_ VGND VGND VPWR VPWR _08705_ sky130_fd_sc_hd__xnor2_1
X_15527_ _05636_ _05637_ net479 net166 VGND VGND VPWR VPWR _05638_ sky130_fd_sc_hd__and4bb_1
X_12739_ _02666_ _02677_ VGND VGND VPWR VPWR _02678_ sky130_fd_sc_hd__nand2_1
X_19295_ clknet_4_8_0_clock _00053_ VGND VGND VPWR VPWR ki\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18246_ _06571_ _06560_ VGND VGND VPWR VPWR _08629_ sky130_fd_sc_hd__and2b_1
XFILLER_0_155_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15458_ _05554_ _05550_ _05552_ VGND VGND VPWR VPWR _05562_ sky130_fd_sc_hd__or3_1
XFILLER_0_60_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14409_ _04398_ _04407_ _04405_ VGND VGND VPWR VPWR _04408_ sky130_fd_sc_hd__a21o_1
X_18177_ _07969_ _07977_ _08048_ VGND VGND VPWR VPWR _08553_ sky130_fd_sc_hd__and3_1
X_15389_ _05412_ _05415_ VGND VGND VPWR VPWR _05486_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17128_ _07396_ _07398_ VGND VGND VPWR VPWR _07399_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09950_ _05732_ VGND VGND VPWR VPWR _06799_ sky130_fd_sc_hd__inv_2
X_17059_ net334 _01755_ _06314_ _07322_ VGND VGND VPWR VPWR _07323_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09881_ _04709_ _06029_ VGND VGND VPWR VPWR _06040_ sky130_fd_sc_hd__and2_1
XFILLER_0_148_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11070_ _01006_ _01008_ VGND VGND VPWR VPWR _01009_ sky130_fd_sc_hd__nand2_1
X_10021_ _07558_ _07569_ VGND VGND VPWR VPWR _07580_ sky130_fd_sc_hd__nor2_1
X_14760_ _04685_ _04793_ VGND VGND VPWR VPWR _04794_ sky130_fd_sc_hd__nor2_1
X_11972_ _01870_ _01904_ VGND VGND VPWR VPWR _01911_ sky130_fd_sc_hd__or2_1
X_13711_ net263 _02330_ _03640_ VGND VGND VPWR VPWR _03677_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10923_ _00859_ _00861_ VGND VGND VPWR VPWR _00862_ sky130_fd_sc_hd__or2b_1
X_14691_ _04715_ _04717_ VGND VGND VPWR VPWR _04718_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16430_ _06628_ _06630_ VGND VGND VPWR VPWR _06631_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13642_ _03596_ _03600_ _03545_ _03601_ VGND VGND VPWR VPWR _03602_ sky130_fd_sc_hd__o211a_1
X_10854_ _00776_ _00792_ VGND VGND VPWR VPWR _00793_ sky130_fd_sc_hd__nand2_2
XFILLER_0_156_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16361_ _06549_ _06554_ VGND VGND VPWR VPWR _06555_ sky130_fd_sc_hd__nand2_2
XFILLER_0_39_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13573_ net265 _02090_ _03530_ _03531_ VGND VGND VPWR VPWR _03532_ sky130_fd_sc_hd__and4_1
XFILLER_0_67_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10785_ _00632_ _00644_ VGND VGND VPWR VPWR _00724_ sky130_fd_sc_hd__xor2_4
XFILLER_0_94_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18100_ _07781_ _07794_ VGND VGND VPWR VPWR _08468_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15312_ _05396_ _05400_ VGND VGND VPWR VPWR _05401_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12524_ _02358_ _02462_ VGND VGND VPWR VPWR _02463_ sky130_fd_sc_hd__nor2_1
X_19080_ _09523_ _00818_ _09525_ net487 VGND VGND VPWR VPWR _00096_ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16292_ _06442_ _06443_ VGND VGND VPWR VPWR _06479_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18031_ _08380_ _08391_ VGND VGND VPWR VPWR _08392_ sky130_fd_sc_hd__or2b_1
XFILLER_0_109_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15243_ _05322_ _05324_ VGND VGND VPWR VPWR _05326_ sky130_fd_sc_hd__xnor2_1
X_12455_ _02393_ _02338_ VGND VGND VPWR VPWR _02394_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11406_ _01282_ _01344_ VGND VGND VPWR VPWR _01345_ sky130_fd_sc_hd__or2_1
X_15174_ _05174_ _05249_ VGND VGND VPWR VPWR _05250_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_111_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12386_ net204 _02224_ VGND VGND VPWR VPWR _02325_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14125_ _03988_ net113 _04095_ _04096_ VGND VGND VPWR VPWR _04097_ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11337_ _01202_ _01245_ _01272_ _01275_ VGND VGND VPWR VPWR _01276_ sky130_fd_sc_hd__a211o_1
X_14056_ _04026_ _04027_ VGND VGND VPWR VPWR _04028_ sky130_fd_sc_hd__nor2_1
X_18933_ net411 net122 net132 _04017_ VGND VGND VPWR VPWR _09385_ sky130_fd_sc_hd__a211o_1
X_11268_ _01205_ _01137_ VGND VGND VPWR VPWR _01207_ sky130_fd_sc_hd__and2b_1
XFILLER_0_120_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13007_ _02808_ _02832_ _02831_ VGND VGND VPWR VPWR _02946_ sky130_fd_sc_hd__a21oi_1
X_10219_ _00156_ _09533_ _00154_ VGND VGND VPWR VPWR _00158_ sky130_fd_sc_hd__or3_1
X_18864_ net218 net215 _01772_ VGND VGND VPWR VPWR _09309_ sky130_fd_sc_hd__o21ai_1
X_11199_ _01065_ _00982_ _01064_ VGND VGND VPWR VPWR _01138_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17815_ _08033_ _08153_ _08151_ _08150_ VGND VGND VPWR VPWR _08155_ sky130_fd_sc_hd__o211a_1
X_18795_ net412 net126 net119 net418 VGND VGND VPWR VPWR _09233_ sky130_fd_sc_hd__a22oi_1
X_17746_ _07490_ _08078_ VGND VGND VPWR VPWR _08079_ sky130_fd_sc_hd__xor2_2
X_14958_ _05009_ _05011_ VGND VGND VPWR VPWR _05012_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13909_ _02570_ _02672_ VGND VGND VPWR VPWR _03877_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17677_ _07986_ _07989_ _08002_ VGND VGND VPWR VPWR _08003_ sky130_fd_sc_hd__o21bai_1
X_14889_ _04870_ _04869_ VGND VGND VPWR VPWR _04936_ sky130_fd_sc_hd__and2b_1
XFILLER_0_89_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16628_ _06845_ _06846_ _06848_ VGND VGND VPWR VPWR _06849_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_58_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16559_ net300 _06352_ _06345_ net296 VGND VGND VPWR VPWR _06773_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19278_ clknet_4_6_0_clock _00074_ VGND VGND VPWR VPWR kp\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18229_ i_error\[14\] _08533_ VGND VGND VPWR VPWR _08610_ sky130_fd_sc_hd__xor2_2
XFILLER_0_32_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09933_ _06590_ _06601_ VGND VGND VPWR VPWR _06612_ sky130_fd_sc_hd__nand2_4
X_09864_ _05666_ _05842_ VGND VGND VPWR VPWR _05853_ sky130_fd_sc_hd__xor2_2
X_09795_ net369 _05072_ _05006_ net365 VGND VGND VPWR VPWR _05094_ sky130_fd_sc_hd__a22oi_2
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10570_ _00412_ _00411_ VGND VGND VPWR VPWR _00509_ sky130_fd_sc_hd__or2b_1
XFILLER_0_119_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12240_ _02038_ _02037_ VGND VGND VPWR VPWR _02179_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12171_ _02019_ _02072_ _02045_ _02071_ VGND VGND VPWR VPWR _02110_ sky130_fd_sc_hd__a211oi_2
X_11122_ _01045_ _01060_ VGND VGND VPWR VPWR _01061_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15930_ _05673_ _05943_ _05945_ VGND VGND VPWR VPWR _06081_ sky130_fd_sc_hd__nor3_2
X_11053_ _00980_ _00977_ VGND VGND VPWR VPWR _00992_ sky130_fd_sc_hd__and2b_1
X_10004_ _07360_ _07382_ VGND VGND VPWR VPWR _07393_ sky130_fd_sc_hd__nand2_4
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15861_ _04216_ _06004_ VGND VGND VPWR VPWR _06005_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17600_ _07916_ _07917_ VGND VGND VPWR VPWR _07918_ sky130_fd_sc_hd__nand2_1
X_14812_ _04847_ _04848_ _04850_ VGND VGND VPWR VPWR _04851_ sky130_fd_sc_hd__and3_1
X_18580_ _08985_ _08995_ VGND VGND VPWR VPWR _08996_ sky130_fd_sc_hd__nand2_1
X_15792_ _05825_ _05928_ VGND VGND VPWR VPWR _05929_ sky130_fd_sc_hd__and2_1
X_17531_ net323 _06618_ _07480_ _07841_ VGND VGND VPWR VPWR _07842_ sky130_fd_sc_hd__a31oi_2
X_14743_ _04747_ _04774_ VGND VGND VPWR VPWR _04776_ sky130_fd_sc_hd__or2_1
X_11955_ _01825_ _01846_ _01893_ VGND VGND VPWR VPWR _01894_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17462_ _07736_ _07753_ _07765_ VGND VGND VPWR VPWR _07766_ sky130_fd_sc_hd__a21bo_1
X_10906_ _00840_ _00844_ VGND VGND VPWR VPWR _00845_ sky130_fd_sc_hd__and2_1
X_14674_ _04688_ _04696_ _04699_ VGND VGND VPWR VPWR _04700_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11886_ _01824_ VGND VGND VPWR VPWR _01825_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19201_ clknet_4_12_0_clock _00083_ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dfxtp_1
X_16413_ _06594_ _06611_ VGND VGND VPWR VPWR _06613_ sky130_fd_sc_hd__nand2_1
X_13625_ _03579_ _03583_ VGND VGND VPWR VPWR _03584_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_157_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10837_ _00768_ _00774_ _00775_ VGND VGND VPWR VPWR _00776_ sky130_fd_sc_hd__o21ai_1
X_17393_ _07673_ _07689_ VGND VGND VPWR VPWR _07691_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19132_ net503 net551 net494 _09557_ VGND VGND VPWR VPWR _00121_ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16344_ net329 VGND VGND VPWR VPWR _06537_ sky130_fd_sc_hd__inv_2
X_13556_ _03511_ _03514_ _03509_ VGND VGND VPWR VPWR _03515_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_81_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10768_ kp\[17\] _00615_ VGND VGND VPWR VPWR _00707_ sky130_fd_sc_hd__nand2_1
X_12507_ _02269_ _02277_ VGND VGND VPWR VPWR _02446_ sky130_fd_sc_hd__xor2_1
X_19063_ _04126_ _09446_ VGND VGND VPWR VPWR _09515_ sky130_fd_sc_hd__nor2_4
XFILLER_0_70_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16275_ _06460_ _06441_ VGND VGND VPWR VPWR _06461_ sky130_fd_sc_hd__xor2_1
X_13487_ net224 _02915_ _03396_ VGND VGND VPWR VPWR _03446_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10699_ net393 _05138_ _05149_ net568 VGND VGND VPWR VPWR _00638_ sky130_fd_sc_hd__a31o_1
X_18014_ _08362_ _08363_ VGND VGND VPWR VPWR _08374_ sky130_fd_sc_hd__nor2_1
X_15226_ net479 net145 _05208_ _05209_ VGND VGND VPWR VPWR _05307_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_140_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12438_ _02361_ _02376_ VGND VGND VPWR VPWR _02377_ sky130_fd_sc_hd__and2b_1
XFILLER_0_140_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15157_ _05214_ _04801_ _05218_ _05216_ VGND VGND VPWR VPWR _05231_ sky130_fd_sc_hd__o22a_1
X_12369_ _01848_ _02091_ VGND VGND VPWR VPWR _02308_ sky130_fd_sc_hd__or2_1
X_14108_ _04075_ _04079_ VGND VGND VPWR VPWR _04080_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15088_ _05132_ _05128_ VGND VGND VPWR VPWR _05155_ sky130_fd_sc_hd__or2b_1
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14039_ _04009_ _04010_ VGND VGND VPWR VPWR _04011_ sky130_fd_sc_hd__and2_1
X_18916_ _02168_ _02169_ _09334_ VGND VGND VPWR VPWR _09366_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_38_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18847_ net206 _01787_ _01810_ net204 VGND VGND VPWR VPWR _09290_ sky130_fd_sc_hd__a22o_1
X_18778_ _09022_ net526 _09008_ VGND VGND VPWR VPWR _09214_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_145_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17729_ _08054_ _08059_ VGND VGND VPWR VPWR _08060_ sky130_fd_sc_hd__xor2_1
XFILLER_0_89_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09916_ _06403_ _06414_ VGND VGND VPWR VPWR _06425_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09847_ _05633_ _05655_ VGND VGND VPWR VPWR _05666_ sky130_fd_sc_hd__nor2_4
XPHY_EDGE_ROW_13_Left_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09778_ net360 _04896_ VGND VGND VPWR VPWR _04907_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11740_ _01212_ _01278_ VGND VGND VPWR VPWR _01679_ sky130_fd_sc_hd__and2_1
XFILLER_0_96_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11671_ _01591_ _01608_ _01609_ VGND VGND VPWR VPWR _01610_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13410_ _03315_ _03317_ VGND VGND VPWR VPWR _03366_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10622_ _00559_ _00560_ VGND VGND VPWR VPWR _00561_ sky130_fd_sc_hd__nand2_1
X_14390_ net451 net128 net125 net456 VGND VGND VPWR VPWR _04387_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_119_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_22_Left_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13341_ net212 _02935_ VGND VGND VPWR VPWR _03294_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10553_ _00490_ _00491_ VGND VGND VPWR VPWR _00492_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16060_ _09098_ _06222_ VGND VGND VPWR VPWR _06224_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13272_ net207 _03220_ _03224_ VGND VGND VPWR VPWR _03225_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10484_ _00396_ _00422_ VGND VGND VPWR VPWR _00423_ sky130_fd_sc_hd__nor2_1
X_15011_ _04941_ VGND VGND VPWR VPWR _05070_ sky130_fd_sc_hd__inv_2
X_12223_ _02160_ _02161_ VGND VGND VPWR VPWR _02162_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12154_ net203 _01910_ _01875_ net205 VGND VGND VPWR VPWR _02093_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11105_ _01042_ _01043_ VGND VGND VPWR VPWR _01044_ sky130_fd_sc_hd__nor2_2
X_16962_ _07214_ _07215_ VGND VGND VPWR VPWR _07216_ sky130_fd_sc_hd__and2b_1
X_12085_ _02023_ _02020_ VGND VGND VPWR VPWR _02024_ sky130_fd_sc_hd__xnor2_1
X_18701_ _09124_ _09128_ VGND VGND VPWR VPWR _09129_ sky130_fd_sc_hd__xnor2_2
X_15913_ _03268_ _03858_ _03339_ _03857_ VGND VGND VPWR VPWR _06063_ sky130_fd_sc_hd__a211o_1
X_11036_ _00935_ _00960_ _00974_ VGND VGND VPWR VPWR _00975_ sky130_fd_sc_hd__nand3_4
X_16893_ _07138_ _07139_ VGND VGND VPWR VPWR _07141_ sky130_fd_sc_hd__xor2_1
X_15844_ _05972_ _05983_ _05986_ VGND VGND VPWR VPWR _05987_ sky130_fd_sc_hd__o21a_1
X_18632_ _06135_ _09052_ VGND VGND VPWR VPWR _09053_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15775_ _05866_ _05888_ VGND VGND VPWR VPWR _05911_ sky130_fd_sc_hd__nand2_1
X_18563_ _08973_ _08976_ VGND VGND VPWR VPWR _08978_ sky130_fd_sc_hd__xor2_1
X_12987_ net207 _02914_ VGND VGND VPWR VPWR _02926_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14726_ net409 net186 _04567_ _04568_ VGND VGND VPWR VPWR _04757_ sky130_fd_sc_hd__o2bb2a_1
X_17514_ net291 _07182_ _07823_ VGND VGND VPWR VPWR _07824_ sky130_fd_sc_hd__and3_1
X_11938_ net200 _01875_ _01876_ VGND VGND VPWR VPWR _01877_ sky130_fd_sc_hd__nand3_1
X_18494_ _08754_ _08755_ _08898_ VGND VGND VPWR VPWR _08902_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17445_ _07667_ _07682_ VGND VGND VPWR VPWR _07748_ sky130_fd_sc_hd__nand2_1
X_14657_ _04613_ _04631_ VGND VGND VPWR VPWR _04681_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11869_ _01807_ VGND VGND VPWR VPWR _01808_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13608_ net243 _02640_ _03566_ VGND VGND VPWR VPWR _03567_ sky130_fd_sc_hd__a21bo_1
X_17376_ _07670_ _07671_ VGND VGND VPWR VPWR _07672_ sky130_fd_sc_hd__and2_1
XFILLER_0_144_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14588_ _04403_ _04604_ VGND VGND VPWR VPWR _04605_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16327_ _06512_ _06517_ VGND VGND VPWR VPWR _06518_ sky130_fd_sc_hd__xnor2_1
X_19115_ _09536_ _05600_ _09547_ net489 VGND VGND VPWR VPWR _00113_ sky130_fd_sc_hd__o211a_1
X_13539_ _03497_ _03418_ VGND VGND VPWR VPWR _03498_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19046_ net522 _09485_ _09456_ VGND VGND VPWR VPWR _09502_ sky130_fd_sc_hd__a21oi_1
X_16258_ net272 _06438_ _06441_ _06439_ VGND VGND VPWR VPWR _06442_ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15209_ _05286_ _05287_ VGND VGND VPWR VPWR _05288_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16189_ net309 net306 _06324_ VGND VGND VPWR VPWR _06366_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09701_ net45 _03870_ _03903_ net347 VGND VGND VPWR VPWR _00062_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09632_ _03347_ VGND VGND VPWR VPWR _03358_ sky130_fd_sc_hd__buf_2
XFILLER_0_148_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout430 net567 VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__buf_2
Xfanout441 net442 VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__clkbuf_4
Xfanout452 net455 VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__clkbuf_4
Xfanout463 net464 VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__clkbuf_2
Xfanout474 net475 VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__clkbuf_2
Xfanout485 net486 VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__clkbuf_4
X_12910_ _02845_ _02848_ VGND VGND VPWR VPWR _02849_ sky130_fd_sc_hd__nand2_1
Xfanout496 net497 VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__clkbuf_4
X_13890_ _03270_ _03338_ VGND VGND VPWR VPWR _03856_ sky130_fd_sc_hd__xnor2_1
X_12841_ net264 _01785_ VGND VGND VPWR VPWR _02780_ sky130_fd_sc_hd__nand2_1
X_15560_ _05612_ _05672_ VGND VGND VPWR VPWR _05674_ sky130_fd_sc_hd__nand2_1
X_12772_ _02697_ _02709_ _02606_ _02710_ VGND VGND VPWR VPWR _02711_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_69_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14511_ _04518_ _04519_ net436 net155 VGND VGND VPWR VPWR _04520_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_68_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11723_ _01578_ _01585_ _01661_ VGND VGND VPWR VPWR _01662_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15491_ _05593_ _05597_ VGND VGND VPWR VPWR _05598_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17230_ _07505_ _07510_ VGND VGND VPWR VPWR _07511_ sky130_fd_sc_hd__xor2_1
X_14442_ net425 net155 net152 net430 VGND VGND VPWR VPWR _04444_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_83_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11654_ _01553_ _01560_ VGND VGND VPWR VPWR _01593_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17161_ _07410_ _07418_ _07416_ VGND VGND VPWR VPWR _07435_ sky130_fd_sc_hd__a21oi_1
X_10605_ _00533_ _00543_ VGND VGND VPWR VPWR _00544_ sky130_fd_sc_hd__xor2_4
X_14373_ _04334_ _04365_ _04366_ VGND VGND VPWR VPWR _04369_ sky130_fd_sc_hd__nand3_1
X_11585_ _01494_ _01496_ _01495_ VGND VGND VPWR VPWR _01524_ sky130_fd_sc_hd__o21a_1
XFILLER_0_52_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16112_ prev_error\[4\] _00406_ _00407_ VGND VGND VPWR VPWR _06281_ sky130_fd_sc_hd__and3_1
X_13324_ _03181_ _03185_ VGND VGND VPWR VPWR _03277_ sky130_fd_sc_hd__xor2_1
XFILLER_0_107_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10536_ net372 _06062_ VGND VGND VPWR VPWR _00475_ sky130_fd_sc_hd__nand2_1
X_17092_ net312 _06353_ _07324_ _07323_ VGND VGND VPWR VPWR _07359_ sky130_fd_sc_hd__a31o_1
XFILLER_0_101_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16043_ _05666_ _06204_ VGND VGND VPWR VPWR _06206_ sky130_fd_sc_hd__xor2_1
X_13255_ net232 net228 _02545_ _02409_ VGND VGND VPWR VPWR _03208_ sky130_fd_sc_hd__nand4_1
XPHY_EDGE_ROW_108_Right_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10467_ _04280_ _00238_ _04335_ VGND VGND VPWR VPWR _00406_ sky130_fd_sc_hd__nand3_2
X_12206_ _02142_ _02144_ VGND VGND VPWR VPWR _02145_ sky130_fd_sc_hd__xnor2_1
X_13186_ _03123_ _03126_ _03138_ VGND VGND VPWR VPWR _03139_ sky130_fd_sc_hd__a21bo_1
X_10398_ _00335_ _00331_ VGND VGND VPWR VPWR _00337_ sky130_fd_sc_hd__and2b_1
XFILLER_0_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12137_ net217 net213 _01861_ _01835_ VGND VGND VPWR VPWR _02076_ sky130_fd_sc_hd__and4_1
X_17994_ net327 _07182_ VGND VGND VPWR VPWR _08352_ sky130_fd_sc_hd__nand2_1
X_16945_ net294 _06723_ _07197_ VGND VGND VPWR VPWR _07198_ sky130_fd_sc_hd__and3_1
X_12068_ _01979_ _02005_ _01987_ VGND VGND VPWR VPWR _02007_ sky130_fd_sc_hd__nor3_1
X_11019_ _00867_ _00956_ VGND VGND VPWR VPWR _00958_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16876_ net329 _06324_ _07120_ _07121_ VGND VGND VPWR VPWR _07122_ sky130_fd_sc_hd__nand4_1
XFILLER_0_35_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18615_ _06046_ _06112_ VGND VGND VPWR VPWR _09035_ sky130_fd_sc_hd__and2_1
X_15827_ _04667_ _04668_ _04664_ VGND VGND VPWR VPWR _05968_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15758_ _05890_ _05865_ _05889_ VGND VGND VPWR VPWR _05892_ sky130_fd_sc_hd__and3_1
X_18546_ _08886_ _08890_ _08615_ _06268_ VGND VGND VPWR VPWR _08959_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14709_ _04728_ _04733_ _04736_ _04737_ VGND VGND VPWR VPWR _04738_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_75_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15689_ _05815_ VGND VGND VPWR VPWR _05816_ sky130_fd_sc_hd__inv_2
X_18477_ _08615_ _08623_ _08882_ VGND VGND VPWR VPWR _08883_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17428_ _07715_ _07728_ VGND VGND VPWR VPWR _07729_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17359_ _07632_ _07633_ _07652_ VGND VGND VPWR VPWR _07653_ sky130_fd_sc_hd__or3_4
XFILLER_0_27_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19029_ _09487_ _09488_ net492 VGND VGND VPWR VPWR _00077_ sky130_fd_sc_hd__o21a_1
XFILLER_0_141_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09615_ net53 _03102_ _03135_ net182 VGND VGND VPWR VPWR _00032_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11370_ _01237_ _01307_ _01308_ VGND VGND VPWR VPWR _01309_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_104_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10321_ _00225_ _00254_ VGND VGND VPWR VPWR _00260_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13040_ _02975_ _02978_ VGND VGND VPWR VPWR _02979_ sky130_fd_sc_hd__and2_1
X_10252_ net379 _04984_ _00190_ VGND VGND VPWR VPWR _00191_ sky130_fd_sc_hd__a21o_1
X_10183_ _09351_ _09329_ VGND VGND VPWR VPWR _09362_ sky130_fd_sc_hd__xor2_1
X_14991_ _04933_ _05047_ VGND VGND VPWR VPWR _05048_ sky130_fd_sc_hd__nor2_1
Xfanout260 net261 VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__buf_2
Xfanout271 ki\[17\] VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__buf_2
Xfanout282 net284 VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__buf_2
X_16730_ net300 _06409_ _06402_ net296 VGND VGND VPWR VPWR _06961_ sky130_fd_sc_hd__a22o_1
X_13942_ net481 _03912_ VGND VGND VPWR VPWR _03913_ sky130_fd_sc_hd__and2_2
Xfanout293 net294 VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__clkbuf_4
X_16661_ _06805_ _06804_ VGND VGND VPWR VPWR _06885_ sky130_fd_sc_hd__and2b_1
X_13873_ _03823_ _03835_ VGND VGND VPWR VPWR _03839_ sky130_fd_sc_hd__or2_1
X_15612_ _05730_ VGND VGND VPWR VPWR _05731_ sky130_fd_sc_hd__inv_2
X_18400_ _08565_ _08556_ VGND VGND VPWR VPWR _08798_ sky130_fd_sc_hd__and2b_1
X_12824_ _02680_ _02731_ _02762_ VGND VGND VPWR VPWR _02763_ sky130_fd_sc_hd__o21a_1
X_16592_ net289 _06402_ _06438_ net286 VGND VGND VPWR VPWR _06809_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_97_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15543_ _05654_ VGND VGND VPWR VPWR _05656_ sky130_fd_sc_hd__inv_2
X_18331_ _08719_ _08721_ VGND VGND VPWR VPWR _08722_ sky130_fd_sc_hd__xnor2_1
X_12755_ _02692_ _02693_ VGND VGND VPWR VPWR _02694_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11706_ _01614_ _01631_ VGND VGND VPWR VPWR _01645_ sky130_fd_sc_hd__xor2_1
X_18262_ _08630_ _08645_ VGND VGND VPWR VPWR _08646_ sky130_fd_sc_hd__xor2_1
X_15474_ _05577_ _05579_ VGND VGND VPWR VPWR _05580_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12686_ _02610_ _02624_ VGND VGND VPWR VPWR _02625_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14425_ _04393_ _04396_ _04424_ VGND VGND VPWR VPWR _04426_ sky130_fd_sc_hd__nand3_1
XFILLER_0_53_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17213_ net315 _06467_ VGND VGND VPWR VPWR _07493_ sky130_fd_sc_hd__nand2_1
X_11637_ _01574_ _01573_ _01575_ VGND VGND VPWR VPWR _01576_ sky130_fd_sc_hd__or3_1
X_18193_ i_error\[5\] _08543_ _08549_ _08568_ _08569_ VGND VGND VPWR VPWR _08571_
+ sky130_fd_sc_hd__a221oi_2
XFILLER_0_126_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17144_ _07414_ _07411_ _07412_ VGND VGND VPWR VPWR _07417_ sky130_fd_sc_hd__and3_1
XFILLER_0_80_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14356_ _04344_ _04347_ _04349_ VGND VGND VPWR VPWR _04350_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_135_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11568_ _01479_ _01505_ _01506_ VGND VGND VPWR VPWR _01507_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13307_ _03231_ _03256_ VGND VGND VPWR VPWR _03260_ sky130_fd_sc_hd__xor2_1
X_17075_ _07339_ _07340_ VGND VGND VPWR VPWR _07341_ sky130_fd_sc_hd__nor2_1
X_10519_ _00429_ _00457_ _00455_ VGND VGND VPWR VPWR _00458_ sky130_fd_sc_hd__a21o_1
X_14287_ _04017_ net160 VGND VGND VPWR VPWR _04274_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11499_ net382 _00410_ _01413_ _01414_ VGND VGND VPWR VPWR _01438_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16026_ _06185_ _06186_ VGND VGND VPWR VPWR _06187_ sky130_fd_sc_hd__and2b_1
X_13238_ net248 _01908_ _03190_ VGND VGND VPWR VPWR _03191_ sky130_fd_sc_hd__nand3_1
XFILLER_0_21_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13169_ _03099_ _03105_ _03107_ VGND VGND VPWR VPWR _03120_ sky130_fd_sc_hd__and3_1
X_17977_ _08330_ _08324_ _08327_ VGND VGND VPWR VPWR _08333_ sky130_fd_sc_hd__nor3_1
X_16928_ _07159_ _07161_ VGND VGND VPWR VPWR _07179_ sky130_fd_sc_hd__xnor2_1
X_16859_ _07092_ _07102_ VGND VGND VPWR VPWR _07103_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18529_ _08927_ _08934_ _08939_ _08926_ VGND VGND VPWR VPWR _08940_ sky130_fd_sc_hd__or4b_1
XFILLER_0_146_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold35 net89 VGND VGND VPWR VPWR net542 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 kd_2\[18\] VGND VGND VPWR VPWR net553 sky130_fd_sc_hd__dlygate4sd3_1
X_10870_ _04236_ _00808_ VGND VGND VPWR VPWR _00809_ sky130_fd_sc_hd__nand2_2
XFILLER_0_79_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12540_ net246 _01799_ _02478_ _02477_ VGND VGND VPWR VPWR _02479_ sky130_fd_sc_hd__a31o_1
XFILLER_0_81_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12471_ _02409_ VGND VGND VPWR VPWR _02410_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_136_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14210_ net428 net433 VGND VGND VPWR VPWR _04189_ sky130_fd_sc_hd__or2_1
X_11422_ _01293_ _01291_ _01292_ VGND VGND VPWR VPWR _01361_ sky130_fd_sc_hd__and3_1
XFILLER_0_124_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15190_ _05169_ _05266_ VGND VGND VPWR VPWR _05267_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14141_ _04106_ _04112_ VGND VGND VPWR VPWR _04113_ sky130_fd_sc_hd__xnor2_1
X_11353_ net374 _00798_ _01001_ net377 VGND VGND VPWR VPWR _01292_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10304_ _00242_ VGND VGND VPWR VPWR _00243_ sky130_fd_sc_hd__clkbuf_4
X_14072_ _03988_ _04043_ VGND VGND VPWR VPWR _04044_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11284_ net377 _00322_ _01145_ VGND VGND VPWR VPWR _01223_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13023_ _02885_ _02890_ VGND VGND VPWR VPWR _02962_ sky130_fd_sc_hd__or2_1
X_17900_ _08245_ _08247_ VGND VGND VPWR VPWR _08248_ sky130_fd_sc_hd__xor2_1
X_10235_ _00161_ _00173_ _00171_ VGND VGND VPWR VPWR _00174_ sky130_fd_sc_hd__o21ba_1
X_18880_ _09324_ _09325_ VGND VGND VPWR VPWR _09326_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_5_Left_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17831_ net313 _07156_ VGND VGND VPWR VPWR _08172_ sky130_fd_sc_hd__nand2_1
X_10166_ net371 _04885_ VGND VGND VPWR VPWR _09175_ sky130_fd_sc_hd__nand2_1
X_17762_ _08090_ _08095_ VGND VGND VPWR VPWR _08096_ sky130_fd_sc_hd__xor2_2
X_10097_ _07767_ _08064_ VGND VGND VPWR VPWR _08416_ sky130_fd_sc_hd__xor2_1
X_14974_ _04965_ _05021_ VGND VGND VPWR VPWR _05030_ sky130_fd_sc_hd__nor2_1
X_16713_ _06364_ _06320_ VGND VGND VPWR VPWR _06943_ sky130_fd_sc_hd__nand2_1
X_13925_ net465 net485 net116 VGND VGND VPWR VPWR _03895_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17693_ net291 _02932_ _08017_ _08019_ VGND VGND VPWR VPWR _08021_ sky130_fd_sc_hd__a31o_1
XFILLER_0_16_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16644_ _06860_ _06866_ VGND VGND VPWR VPWR _06867_ sky130_fd_sc_hd__xnor2_1
X_13856_ _03820_ _03821_ _03807_ VGND VGND VPWR VPWR _03822_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12807_ _02745_ VGND VGND VPWR VPWR _02746_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16575_ _06767_ _06769_ VGND VGND VPWR VPWR _06791_ sky130_fd_sc_hd__nor2_1
X_13787_ net267 net251 _02913_ _02408_ VGND VGND VPWR VPWR _03753_ sky130_fd_sc_hd__nand4_1
XFILLER_0_57_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10999_ _00844_ _00925_ _00936_ VGND VGND VPWR VPWR _00938_ sky130_fd_sc_hd__nand3_1
XFILLER_0_85_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18314_ net279 _06316_ _06318_ _08701_ _08703_ VGND VGND VPWR VPWR _08704_ sky130_fd_sc_hd__a41o_1
X_15526_ net471 net176 net171 net476 VGND VGND VPWR VPWR _05637_ sky130_fd_sc_hd__a22oi_1
X_12738_ _02664_ _02665_ VGND VGND VPWR VPWR _02677_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19294_ clknet_4_8_0_clock _00052_ VGND VGND VPWR VPWR ki\[5\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15457_ _05559_ _05560_ VGND VGND VPWR VPWR _05561_ sky130_fd_sc_hd__xnor2_1
X_18245_ _06376_ _06570_ VGND VGND VPWR VPWR _08628_ sky130_fd_sc_hd__nor2_1
X_12669_ _02597_ _02603_ _02595_ VGND VGND VPWR VPWR _02608_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_115_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14408_ _04405_ _04406_ VGND VGND VPWR VPWR _04407_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15388_ _05482_ _05484_ VGND VGND VPWR VPWR _05485_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18176_ _08550_ _08551_ i_error\[3\] VGND VGND VPWR VPWR _08552_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17127_ _07077_ _07397_ VGND VGND VPWR VPWR _07398_ sky130_fd_sc_hd__and2_1
X_14339_ _03896_ _04311_ VGND VGND VPWR VPWR _04331_ sky130_fd_sc_hd__or2b_1
XFILLER_0_40_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17058_ net317 _06334_ VGND VGND VPWR VPWR _07322_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16009_ _00464_ _06167_ VGND VGND VPWR VPWR _06168_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_111_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09880_ net562 _04687_ _04698_ VGND VGND VPWR VPWR _06029_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10020_ _07360_ _07547_ _07415_ VGND VGND VPWR VPWR _07569_ sky130_fd_sc_hd__and3_1
XFILLER_0_99_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11971_ _01909_ VGND VGND VPWR VPWR _01910_ sky130_fd_sc_hd__buf_2
X_13710_ net263 _02408_ _03675_ VGND VGND VPWR VPWR _03676_ sky130_fd_sc_hd__and3_1
XFILLER_0_98_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10922_ _00793_ _00795_ _00860_ VGND VGND VPWR VPWR _00861_ sky130_fd_sc_hd__a21o_1
X_14690_ _04700_ _04716_ VGND VGND VPWR VPWR _04717_ sky130_fd_sc_hd__nand2_1
X_13641_ _03541_ _03544_ _03543_ VGND VGND VPWR VPWR _03601_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10853_ _00789_ _00791_ VGND VGND VPWR VPWR _00792_ sky130_fd_sc_hd__or2b_1
XFILLER_0_156_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16360_ _06536_ _06553_ VGND VGND VPWR VPWR _06554_ sky130_fd_sc_hd__nand2_1
X_13572_ net262 _02222_ _02330_ net258 VGND VGND VPWR VPWR _03531_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10784_ _00695_ _00722_ VGND VGND VPWR VPWR _00723_ sky130_fd_sc_hd__nor2_2
XFILLER_0_66_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15311_ _05397_ _05398_ _05399_ VGND VGND VPWR VPWR _05400_ sky130_fd_sc_hd__o21ba_1
X_12523_ _02360_ _02458_ _02461_ VGND VGND VPWR VPWR _02462_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_137_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16291_ _06475_ _06477_ VGND VGND VPWR VPWR _06478_ sky130_fd_sc_hd__and2b_1
XFILLER_0_152_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15242_ _05230_ _05323_ VGND VGND VPWR VPWR _05324_ sky130_fd_sc_hd__nor2_1
X_18030_ _08364_ _08374_ VGND VGND VPWR VPWR _08391_ sky130_fd_sc_hd__or2_1
X_12454_ _01848_ _02224_ VGND VGND VPWR VPWR _02393_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11405_ _01314_ _01342_ _01343_ VGND VGND VPWR VPWR _01344_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_152_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15173_ net423 net193 VGND VGND VPWR VPWR _05249_ sky130_fd_sc_hd__nand2_1
X_12385_ net205 _02091_ VGND VGND VPWR VPWR _02324_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14124_ _04067_ _04068_ _04094_ VGND VGND VPWR VPWR _04096_ sky130_fd_sc_hd__o21ai_1
X_11336_ _01273_ _01274_ VGND VGND VPWR VPWR _01275_ sky130_fd_sc_hd__and2b_1
X_14055_ net408 net150 _04024_ _04025_ VGND VGND VPWR VPWR _04027_ sky130_fd_sc_hd__o2bb2a_1
X_18932_ _09311_ _09382_ VGND VGND VPWR VPWR _09383_ sky130_fd_sc_hd__xnor2_1
X_11267_ _01137_ _01205_ VGND VGND VPWR VPWR _01206_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_120_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13006_ _02912_ _02944_ VGND VGND VPWR VPWR _02945_ sky130_fd_sc_hd__xnor2_1
X_10218_ _09533_ _00154_ _00156_ VGND VGND VPWR VPWR _00157_ sky130_fd_sc_hd__o21ai_1
X_18863_ _02152_ _02153_ _02146_ VGND VGND VPWR VPWR _09308_ sky130_fd_sc_hd__a21boi_1
X_11198_ _01126_ _01127_ VGND VGND VPWR VPWR _01137_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_27_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17814_ _08150_ _08151_ _08153_ _08033_ VGND VGND VPWR VPWR _08154_ sky130_fd_sc_hd__a211oi_4
X_10149_ _08834_ _07525_ _08977_ VGND VGND VPWR VPWR _08988_ sky130_fd_sc_hd__o21a_1
X_18794_ net408 net130 VGND VGND VPWR VPWR _09232_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17745_ net314 _06889_ VGND VGND VPWR VPWR _08078_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14957_ _04903_ _05010_ VGND VGND VPWR VPWR _05011_ sky130_fd_sc_hd__xnor2_1
X_13908_ _02873_ _03873_ _03875_ VGND VGND VPWR VPWR _03876_ sky130_fd_sc_hd__a21o_1
X_17676_ net315 _06802_ _07462_ VGND VGND VPWR VPWR _08002_ sky130_fd_sc_hd__and3_1
X_14888_ net413 net190 VGND VGND VPWR VPWR _04935_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_59_Left_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16627_ net306 _06310_ _06847_ VGND VGND VPWR VPWR _06848_ sky130_fd_sc_hd__and3_1
X_13839_ _03798_ _03804_ VGND VGND VPWR VPWR _03805_ sky130_fd_sc_hd__or2b_1
XFILLER_0_58_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16558_ _06771_ _06688_ VGND VGND VPWR VPWR _06772_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15509_ net467 net178 net157 net484 VGND VGND VPWR VPWR _05618_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19277_ clknet_4_6_0_clock _00073_ VGND VGND VPWR VPWR kp\[7\] sky130_fd_sc_hd__dfxtp_2
X_16489_ _06684_ _06695_ VGND VGND VPWR VPWR _06696_ sky130_fd_sc_hd__xor2_2
X_18228_ i_error\[13\] _08535_ _08606_ i_error\[12\] VGND VGND VPWR VPWR _08609_ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18159_ _08531_ _08532_ VGND VGND VPWR VPWR _08533_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_102_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_68_Left_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09932_ _04621_ _06579_ _04533_ VGND VGND VPWR VPWR _06601_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_111_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09863_ _05820_ _05831_ VGND VGND VPWR VPWR _05842_ sky130_fd_sc_hd__nand2_1
X_09794_ net368 net365 _05072_ VGND VGND VPWR VPWR _05083_ sky130_fd_sc_hd__and3_1
XFILLER_0_84_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_77_Left_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_86_Left_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12170_ _02107_ _02108_ VGND VGND VPWR VPWR _02109_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11121_ _01052_ _01059_ VGND VGND VPWR VPWR _01060_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11052_ _00975_ _00988_ _00989_ _00990_ VGND VGND VPWR VPWR _00991_ sky130_fd_sc_hd__a211oi_2
X_10003_ _07371_ _07316_ _07272_ VGND VGND VPWR VPWR _07382_ sky130_fd_sc_hd__or3b_4
X_15860_ _04299_ _06003_ VGND VGND VPWR VPWR _06004_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_95_Left_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14811_ _04828_ _04849_ VGND VGND VPWR VPWR _04850_ sky130_fd_sc_hd__nor2_1
X_15791_ _05822_ _05824_ VGND VGND VPWR VPWR _05928_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17530_ net323 _06463_ _06465_ _06618_ net319 VGND VGND VPWR VPWR _07841_ sky130_fd_sc_hd__a32oi_2
X_11954_ _01855_ _01892_ VGND VGND VPWR VPWR _01893_ sky130_fd_sc_hd__xnor2_1
X_14742_ _04746_ _04721_ _04744_ VGND VGND VPWR VPWR _04774_ sky130_fd_sc_hd__and3_1
XFILLER_0_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10905_ _00841_ _00842_ _00843_ VGND VGND VPWR VPWR _00844_ sky130_fd_sc_hd__nand3_1
X_14673_ _04626_ _04697_ VGND VGND VPWR VPWR _04699_ sky130_fd_sc_hd__or2_1
X_17461_ _07670_ _07684_ _07754_ VGND VGND VPWR VPWR _07765_ sky130_fd_sc_hd__or3_1
X_11885_ _01783_ _01823_ VGND VGND VPWR VPWR _01824_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19200_ clknet_4_14_0_clock _00082_ VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dfxtp_1
X_13624_ _03574_ _03577_ VGND VGND VPWR VPWR _03583_ sky130_fd_sc_hd__nor2_1
X_16412_ _06608_ _06610_ VGND VGND VPWR VPWR _06611_ sky130_fd_sc_hd__or2b_1
XFILLER_0_39_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10836_ _00689_ _00691_ VGND VGND VPWR VPWR _00775_ sky130_fd_sc_hd__xnor2_1
X_17392_ _07687_ _07688_ VGND VGND VPWR VPWR _07689_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19131_ _09080_ _09081_ net563 VGND VGND VPWR VPWR _09557_ sky130_fd_sc_hd__a21o_1
X_13555_ net237 _02747_ _03512_ _03513_ VGND VGND VPWR VPWR _03514_ sky130_fd_sc_hd__a31o_1
X_16343_ _06373_ _06374_ VGND VGND VPWR VPWR _06536_ sky130_fd_sc_hd__xnor2_1
X_10767_ net359 _00245_ _00503_ _00705_ VGND VGND VPWR VPWR _00706_ sky130_fd_sc_hd__a31o_1
X_12506_ _02442_ _02444_ VGND VGND VPWR VPWR _02445_ sky130_fd_sc_hd__nor2_1
X_19062_ _09218_ _09512_ _09513_ VGND VGND VPWR VPWR _00088_ sky130_fd_sc_hd__a21oi_1
X_16274_ net272 _06438_ VGND VGND VPWR VPWR _06460_ sky130_fd_sc_hd__nand2_1
X_13486_ _03442_ _03443_ VGND VGND VPWR VPWR _03445_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10698_ net401 _05061_ _00537_ _00538_ VGND VGND VPWR VPWR _00637_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15225_ _05304_ _05305_ net482 net149 VGND VGND VPWR VPWR _05306_ sky130_fd_sc_hd__and4bb_1
X_18013_ _08351_ _08371_ VGND VGND VPWR VPWR _08373_ sky130_fd_sc_hd__or2b_1
X_12437_ _02366_ _02369_ _02375_ VGND VGND VPWR VPWR _02376_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_152_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15156_ _05228_ _05229_ net450 net172 VGND VGND VPWR VPWR _05230_ sky130_fd_sc_hd__and4bb_1
X_12368_ _02280_ _02282_ _02299_ VGND VGND VPWR VPWR _02307_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_50_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14107_ net435 _03940_ _04078_ VGND VGND VPWR VPWR _04079_ sky130_fd_sc_hd__o21ai_1
X_11319_ _06590_ _06601_ _01257_ _00440_ VGND VGND VPWR VPWR _01258_ sky130_fd_sc_hd__a211o_1
X_15087_ _05124_ _05126_ VGND VGND VPWR VPWR _05154_ sky130_fd_sc_hd__or2b_1
X_12299_ _02189_ _02201_ _02236_ VGND VGND VPWR VPWR _02238_ sky130_fd_sc_hd__and3_1
X_14038_ _03972_ _03974_ _04008_ VGND VGND VPWR VPWR _04010_ sky130_fd_sc_hd__or3_1
X_18915_ _09361_ _09364_ VGND VGND VPWR VPWR _09365_ sky130_fd_sc_hd__xnor2_2
X_18846_ net203 _01787_ VGND VGND VPWR VPWR _09289_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18777_ _09210_ _09212_ VGND VGND VPWR VPWR _09213_ sky130_fd_sc_hd__xnor2_1
X_15989_ _01671_ _01673_ VGND VGND VPWR VPWR _06146_ sky130_fd_sc_hd__xor2_4
X_17728_ net318 _06991_ VGND VGND VPWR VPWR _08059_ sky130_fd_sc_hd__nand2_1
X_17659_ net328 _06467_ _07886_ _07887_ VGND VGND VPWR VPWR _07983_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19329_ clknet_4_2_0_clock _00030_ VGND VGND VPWR VPWR kd_2\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09915_ _06392_ _06128_ _06271_ VGND VGND VPWR VPWR _06414_ sky130_fd_sc_hd__nor3_1
X_09846_ _05556_ _05589_ _05644_ VGND VGND VPWR VPWR _05655_ sky130_fd_sc_hd__o21a_1
X_09777_ _04885_ VGND VGND VPWR VPWR _04896_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11670_ _01592_ _01607_ VGND VGND VPWR VPWR _01609_ sky130_fd_sc_hd__and2b_1
XFILLER_0_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10621_ _00359_ _00461_ VGND VGND VPWR VPWR _00560_ sky130_fd_sc_hd__xor2_1
XFILLER_0_154_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13340_ _03288_ _03292_ VGND VGND VPWR VPWR _03293_ sky130_fd_sc_hd__xnor2_1
X_10552_ _00489_ _00485_ VGND VGND VPWR VPWR _00491_ sky130_fd_sc_hd__or2b_1
XFILLER_0_63_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13271_ net212 _03220_ _03222_ _03223_ VGND VGND VPWR VPWR _03224_ sky130_fd_sc_hd__a31o_1
X_10483_ _00378_ _00393_ _00395_ VGND VGND VPWR VPWR _00422_ sky130_fd_sc_hd__and3_1
X_15010_ net423 net189 _05067_ _05068_ VGND VGND VPWR VPWR _05069_ sky130_fd_sc_hd__a31o_1
X_12222_ _01979_ _02159_ _02003_ VGND VGND VPWR VPWR _02161_ sky130_fd_sc_hd__nor3_1
X_12153_ net200 _02091_ VGND VGND VPWR VPWR _02092_ sky130_fd_sc_hd__nand2_1
X_11104_ _01039_ _01041_ _01040_ VGND VGND VPWR VPWR _01043_ sky130_fd_sc_hd__a21oi_1
X_16961_ _07212_ _07213_ VGND VGND VPWR VPWR _07215_ sky130_fd_sc_hd__nand2_1
X_12084_ _01987_ _02010_ VGND VGND VPWR VPWR _02023_ sky130_fd_sc_hd__or2_1
X_18700_ _08930_ _08963_ _09127_ VGND VGND VPWR VPWR _09128_ sky130_fd_sc_hd__o21ai_2
X_15912_ _05295_ _05954_ VGND VGND VPWR VPWR _06061_ sky130_fd_sc_hd__xor2_2
X_11035_ _00968_ _00972_ _00973_ VGND VGND VPWR VPWR _00974_ sky130_fd_sc_hd__a21o_1
X_16892_ _07013_ _07027_ VGND VGND VPWR VPWR _07139_ sky130_fd_sc_hd__xnor2_1
X_18631_ _09048_ _09051_ VGND VGND VPWR VPWR _09052_ sky130_fd_sc_hd__xor2_1
X_15843_ _04474_ _05984_ VGND VGND VPWR VPWR _05986_ sky130_fd_sc_hd__nor2_1
X_18562_ _08893_ _08975_ _08964_ VGND VGND VPWR VPWR _08976_ sky130_fd_sc_hd__mux2_2
X_15774_ _05907_ _05909_ VGND VGND VPWR VPWR _05910_ sky130_fd_sc_hd__nand2_1
X_12986_ _02924_ _02852_ VGND VGND VPWR VPWR _02925_ sky130_fd_sc_hd__xnor2_1
X_17513_ _07556_ _07821_ VGND VGND VPWR VPWR _07823_ sky130_fd_sc_hd__xor2_1
X_14725_ _04754_ _04755_ net421 net175 VGND VGND VPWR VPWR _04756_ sky130_fd_sc_hd__and4bb_1
X_11937_ _01869_ _01870_ VGND VGND VPWR VPWR _01876_ sky130_fd_sc_hd__xor2_1
X_18493_ _08898_ _08754_ _08755_ _08764_ _08899_ VGND VGND VPWR VPWR _08901_ sky130_fd_sc_hd__a32o_2
XFILLER_0_24_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17444_ _07744_ _07746_ VGND VGND VPWR VPWR _07747_ sky130_fd_sc_hd__nor2_1
X_11868_ _01806_ VGND VGND VPWR VPWR _01807_ sky130_fd_sc_hd__buf_2
XFILLER_0_28_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14656_ _04581_ _04679_ VGND VGND VPWR VPWR _04680_ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13607_ net240 _02745_ VGND VGND VPWR VPWR _03566_ sky130_fd_sc_hd__nand2_1
X_10819_ _00755_ _00756_ VGND VGND VPWR VPWR _00758_ sky130_fd_sc_hd__or2_1
X_17375_ _07565_ _07572_ _07669_ VGND VGND VPWR VPWR _07671_ sky130_fd_sc_hd__nand3_1
X_14587_ _04399_ _04402_ VGND VGND VPWR VPWR _04604_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11799_ prev_error\[12\] VGND VGND VPWR VPWR _01738_ sky130_fd_sc_hd__inv_2
X_19114_ net500 prev_error\[18\] VGND VGND VPWR VPWR _09547_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16326_ _06515_ _06516_ VGND VGND VPWR VPWR _06517_ sky130_fd_sc_hd__nor2_1
X_13538_ _03411_ _03413_ VGND VGND VPWR VPWR _03497_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19045_ _04126_ net96 VGND VGND VPWR VPWR _09501_ sky130_fd_sc_hd__and2_1
X_13469_ net236 _02546_ VGND VGND VPWR VPWR _03428_ sky130_fd_sc_hd__nand2_1
X_16257_ _06439_ _06440_ VGND VGND VPWR VPWR _06441_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15208_ net112 _05285_ _05265_ _05284_ VGND VGND VPWR VPWR _05287_ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16188_ net312 _06328_ _06362_ _06364_ VGND VGND VPWR VPWR _06365_ sky130_fd_sc_hd__a31o_2
XFILLER_0_140_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15139_ net479 net139 _05106_ _05107_ VGND VGND VPWR VPWR _05211_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09700_ net44 _03870_ _03903_ net351 VGND VGND VPWR VPWR _00061_ sky130_fd_sc_hd__a22o_1
X_09631_ _03069_ _03336_ VGND VGND VPWR VPWR _03347_ sky130_fd_sc_hd__nor2_4
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18829_ _04209_ _09226_ _09269_ VGND VGND VPWR VPWR _09270_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout420 net421 VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__clkbuf_2
Xfanout431 prev_d_error\[12\] VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__buf_1
Xfanout442 prev_d_error\[10\] VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__buf_2
Xfanout453 net454 VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__clkbuf_4
Xfanout464 prev_d_error\[5\] VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__buf_2
Xfanout475 net477 VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__buf_2
Xfanout486 prev_d_error\[0\] VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__clkbuf_4
X_09829_ _05270_ _05457_ VGND VGND VPWR VPWR _05468_ sky130_fd_sc_hd__or2_1
Xfanout497 net59 VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__clkbuf_4
X_12840_ net268 net111 VGND VGND VPWR VPWR _02779_ sky130_fd_sc_hd__nand2_1
X_12771_ _02591_ _02605_ _02604_ VGND VGND VPWR VPWR _02710_ sky130_fd_sc_hd__a21o_1
X_14510_ net439 net152 net147 net445 VGND VGND VPWR VPWR _04519_ sky130_fd_sc_hd__a22oi_1
X_11722_ _01611_ _01659_ _01585_ _01660_ VGND VGND VPWR VPWR _01661_ sky130_fd_sc_hd__o211a_1
X_15490_ _05595_ _05596_ VGND VGND VPWR VPWR _05597_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14441_ net425 net430 net155 net152 VGND VGND VPWR VPWR _04443_ sky130_fd_sc_hd__and4_1
X_11653_ _01568_ _01570_ VGND VGND VPWR VPWR _01592_ sky130_fd_sc_hd__xor2_1
XFILLER_0_126_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10604_ _00535_ _00541_ _00542_ VGND VGND VPWR VPWR _00543_ sky130_fd_sc_hd__a21oi_2
X_17160_ _07432_ _07433_ VGND VGND VPWR VPWR _07434_ sky130_fd_sc_hd__xor2_1
X_14372_ _04334_ _04365_ _04366_ VGND VGND VPWR VPWR _04367_ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11584_ _01521_ _01522_ VGND VGND VPWR VPWR _01523_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13323_ net252 _01908_ _02880_ _03275_ VGND VGND VPWR VPWR _03276_ sky130_fd_sc_hd__a31o_1
X_16111_ _02637_ _06278_ _06279_ VGND VGND VPWR VPWR _06280_ sky130_fd_sc_hd__a21o_2
XFILLER_0_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10535_ _00470_ _00473_ VGND VGND VPWR VPWR _00474_ sky130_fd_sc_hd__xor2_4
X_17091_ _07057_ _07212_ _07339_ VGND VGND VPWR VPWR _07358_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_150_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16042_ _06920_ _06203_ VGND VGND VPWR VPWR _06204_ sky130_fd_sc_hd__xor2_2
X_13254_ net224 _02641_ VGND VGND VPWR VPWR _03207_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10466_ _00399_ _00402_ _00404_ VGND VGND VPWR VPWR _00405_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12205_ _01953_ _01965_ _02143_ VGND VGND VPWR VPWR _02144_ sky130_fd_sc_hd__a21oi_1
X_13185_ _03127_ _03128_ _03137_ VGND VGND VPWR VPWR _03138_ sky130_fd_sc_hd__or3_1
XFILLER_0_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10397_ _00331_ _00335_ VGND VGND VPWR VPWR _00336_ sky130_fd_sc_hd__and2b_1
XFILLER_0_103_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12136_ _01918_ _02074_ VGND VGND VPWR VPWR _02075_ sky130_fd_sc_hd__nand2_1
X_17993_ _08343_ _08349_ VGND VGND VPWR VPWR _08351_ sky130_fd_sc_hd__nand2_1
X_16944_ _07194_ _07196_ VGND VGND VPWR VPWR _07197_ sky130_fd_sc_hd__nor2_1
X_12067_ _01979_ _01987_ _02005_ VGND VGND VPWR VPWR _02006_ sky130_fd_sc_hd__o21a_1
X_11018_ _00867_ _00956_ VGND VGND VPWR VPWR _00957_ sky130_fd_sc_hd__nand2_1
X_16875_ net324 _06314_ _06318_ _06309_ net320 VGND VGND VPWR VPWR _07121_ sky130_fd_sc_hd__a32o_1
XFILLER_0_35_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18614_ _06134_ _09030_ VGND VGND VPWR VPWR _09034_ sky130_fd_sc_hd__xor2_1
X_15826_ _05960_ _05964_ _05966_ VGND VGND VPWR VPWR _05967_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18545_ _08917_ _08957_ _06268_ _08615_ VGND VGND VPWR VPWR _08958_ sky130_fd_sc_hd__o2bb2a_4
X_15757_ _05865_ _05889_ _05890_ VGND VGND VPWR VPWR _05891_ sky130_fd_sc_hd__a21oi_1
X_12969_ _02905_ _02907_ VGND VGND VPWR VPWR _02908_ sky130_fd_sc_hd__and2b_1
XFILLER_0_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14708_ _04710_ _04713_ _04735_ VGND VGND VPWR VPWR _04737_ sky130_fd_sc_hd__nand3_1
X_18476_ _08881_ VGND VGND VPWR VPWR _08882_ sky130_fd_sc_hd__buf_4
XFILLER_0_28_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15688_ _05814_ _05811_ VGND VGND VPWR VPWR _05815_ sky130_fd_sc_hd__xor2_2
XFILLER_0_142_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17427_ _07717_ _07727_ VGND VGND VPWR VPWR _07728_ sky130_fd_sc_hd__xor2_2
XFILLER_0_118_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14639_ _04658_ _04660_ VGND VGND VPWR VPWR _04661_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17358_ _07636_ _07651_ VGND VGND VPWR VPWR _07652_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16309_ _06496_ _06497_ VGND VGND VPWR VPWR _06498_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17289_ _07574_ _07575_ VGND VGND VPWR VPWR _07576_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19028_ _09448_ _09485_ _09475_ VGND VGND VPWR VPWR _09488_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_141_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_41_Left_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09614_ net52 _03102_ _03135_ net186 VGND VGND VPWR VPWR _00031_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10320_ _00187_ _00258_ VGND VGND VPWR VPWR _00259_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_61_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10251_ net375 _04841_ _04852_ VGND VGND VPWR VPWR _00190_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10182_ _07899_ _09285_ VGND VGND VPWR VPWR _09351_ sky130_fd_sc_hd__or2_1
Xfanout250 net253 VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__clkbuf_4
X_14990_ net422 net186 _04931_ _05046_ VGND VGND VPWR VPWR _05047_ sky130_fd_sc_hd__o2bb2a_1
Xfanout261 kd_1\[2\] VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__buf_2
Xfanout272 ki\[17\] VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__buf_2
X_13941_ net470 net475 net116 VGND VGND VPWR VPWR _03912_ sky130_fd_sc_hd__and3_1
Xfanout283 net284 VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__clkbuf_4
Xfanout294 ki\[11\] VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__clkbuf_4
X_16660_ net271 _06803_ VGND VGND VPWR VPWR _06884_ sky130_fd_sc_hd__nand2_1
X_13872_ _03808_ _03820_ _03821_ VGND VGND VPWR VPWR _03838_ sky130_fd_sc_hd__or3_1
XFILLER_0_97_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15611_ _05725_ _05727_ _05728_ _05729_ VGND VGND VPWR VPWR _05730_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_97_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12823_ _02760_ _02761_ VGND VGND VPWR VPWR _02762_ sky130_fd_sc_hd__nand2_1
X_16591_ net286 _06402_ _06807_ VGND VGND VPWR VPWR _06808_ sky130_fd_sc_hd__and3_1
X_18330_ _08654_ _08666_ _08720_ VGND VGND VPWR VPWR _08721_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_141_Right_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15542_ _05651_ _05653_ VGND VGND VPWR VPWR _05654_ sky130_fd_sc_hd__nand2_1
X_12754_ _02683_ _02687_ VGND VGND VPWR VPWR _02693_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11705_ _01623_ _01624_ VGND VGND VPWR VPWR _01644_ sky130_fd_sc_hd__xnor2_1
X_18261_ _08643_ _08644_ VGND VGND VPWR VPWR _08645_ sky130_fd_sc_hd__nor2_1
X_12685_ _02612_ _02619_ _02623_ VGND VGND VPWR VPWR _02624_ sky130_fd_sc_hd__a21oi_1
X_15473_ _05576_ _05572_ VGND VGND VPWR VPWR _05579_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17212_ net316 _06344_ _07490_ VGND VGND VPWR VPWR _07491_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14424_ _04393_ _04396_ _04424_ VGND VGND VPWR VPWR _04425_ sky130_fd_sc_hd__a21o_1
X_11636_ _01544_ _01572_ _01563_ _01571_ VGND VGND VPWR VPWR _01575_ sky130_fd_sc_hd__a211oi_1
X_18192_ i_error\[4\] _08547_ VGND VGND VPWR VPWR _08569_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17143_ _07411_ _07412_ _07414_ VGND VGND VPWR VPWR _07416_ sky130_fd_sc_hd__a21oi_1
X_14355_ _04266_ _04348_ VGND VGND VPWR VPWR _04349_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11567_ _01481_ _01504_ VGND VGND VPWR VPWR _01506_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13306_ _03229_ _03258_ VGND VGND VPWR VPWR _03259_ sky130_fd_sc_hd__nor2_1
X_10518_ _00455_ _00456_ VGND VGND VPWR VPWR _00457_ sky130_fd_sc_hd__nor2_1
X_17074_ net304 _06402_ _07337_ VGND VGND VPWR VPWR _07340_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14286_ _04263_ _04270_ _04272_ VGND VGND VPWR VPWR _04273_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_123_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11498_ _01379_ _01433_ _01436_ VGND VGND VPWR VPWR _01437_ sky130_fd_sc_hd__nand3_1
XFILLER_0_122_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16025_ net349 _05677_ _08889_ _07448_ VGND VGND VPWR VPWR _06186_ sky130_fd_sc_hd__a31o_1
X_13237_ _03187_ _03188_ VGND VGND VPWR VPWR _03190_ sky130_fd_sc_hd__xor2_1
X_10449_ _00386_ _00381_ VGND VGND VPWR VPWR _00388_ sky130_fd_sc_hd__or2b_1
XFILLER_0_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13168_ _03110_ _03114_ _03118_ VGND VGND VPWR VPWR _03119_ sky130_fd_sc_hd__a21oi_1
X_12119_ net221 _01814_ VGND VGND VPWR VPWR _02058_ sky130_fd_sc_hd__nand2_1
X_13099_ _03035_ _03042_ VGND VGND VPWR VPWR _03043_ sky130_fd_sc_hd__and2b_1
X_17976_ net313 _02931_ _08321_ VGND VGND VPWR VPWR _08332_ sky130_fd_sc_hd__a21o_1
X_16927_ _07165_ _07174_ _07177_ VGND VGND VPWR VPWR _07178_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16858_ _07090_ _07091_ VGND VGND VPWR VPWR _07102_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15809_ _05469_ _05470_ _05544_ VGND VGND VPWR VPWR _05948_ sky130_fd_sc_hd__nor3_1
XFILLER_0_149_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16789_ _06541_ _07023_ _07024_ VGND VGND VPWR VPWR _07026_ sky130_fd_sc_hd__nand3_1
XFILLER_0_88_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18528_ _08799_ _08935_ _08937_ _08938_ VGND VGND VPWR VPWR _08939_ sky130_fd_sc_hd__a211o_1
XFILLER_0_1_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18459_ _08858_ _08862_ VGND VGND VPWR VPWR _08863_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold36 net87 VGND VGND VPWR VPWR net543 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 i_error\[17\] VGND VGND VPWR VPWR net554 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12470_ _02408_ VGND VGND VPWR VPWR _02409_ sky130_fd_sc_hd__buf_2
XFILLER_0_53_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11421_ net381 _00324_ _01357_ _01359_ VGND VGND VPWR VPWR _01360_ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14140_ _04109_ _04111_ VGND VGND VPWR VPWR _04112_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11352_ net373 _00515_ VGND VGND VPWR VPWR _01291_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10303_ _09552_ _04478_ _00241_ VGND VGND VPWR VPWR _00242_ sky130_fd_sc_hd__and3_2
XFILLER_0_131_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14071_ _03954_ _03987_ VGND VGND VPWR VPWR _04043_ sky130_fd_sc_hd__nor2_1
X_11283_ net377 _00243_ _00323_ net374 VGND VGND VPWR VPWR _01222_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_104_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13022_ _02955_ _02959_ _02960_ VGND VGND VPWR VPWR _02961_ sky130_fd_sc_hd__a21o_1
X_10234_ _00171_ _00172_ VGND VGND VPWR VPWR _00173_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17830_ _07897_ _08170_ VGND VGND VPWR VPWR _08171_ sky130_fd_sc_hd__xor2_2
X_10165_ _09153_ _05545_ VGND VGND VPWR VPWR _09164_ sky130_fd_sc_hd__and2b_1
X_17761_ _08091_ _08094_ VGND VGND VPWR VPWR _08095_ sky130_fd_sc_hd__xnor2_2
X_10096_ _08130_ _08394_ VGND VGND VPWR VPWR _08405_ sky130_fd_sc_hd__xor2_1
X_14973_ _05027_ _05007_ VGND VGND VPWR VPWR _05029_ sky130_fd_sc_hd__xnor2_1
X_16712_ _06939_ _06940_ VGND VGND VPWR VPWR _06941_ sky130_fd_sc_hd__xnor2_2
X_13924_ net461 net116 VGND VGND VPWR VPWR _03894_ sky130_fd_sc_hd__nand2_1
X_17692_ _07926_ _08018_ VGND VGND VPWR VPWR _08019_ sky130_fd_sc_hd__nor2_1
X_16643_ net294 _06404_ _06864_ _06862_ VGND VGND VPWR VPWR _06866_ sky130_fd_sc_hd__a31o_1
X_13855_ _03788_ _03806_ VGND VGND VPWR VPWR _03821_ sky130_fd_sc_hd__xor2_2
XFILLER_0_57_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12806_ _01719_ _02744_ VGND VGND VPWR VPWR _02745_ sky130_fd_sc_hd__xnor2_4
X_16574_ _06783_ _06787_ _06789_ VGND VGND VPWR VPWR _06790_ sky130_fd_sc_hd__o21ba_1
X_13786_ _03749_ _03751_ VGND VGND VPWR VPWR _03752_ sky130_fd_sc_hd__or2_1
X_10998_ _00844_ _00925_ _00936_ VGND VGND VPWR VPWR _00937_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18313_ net279 _06379_ _08701_ VGND VGND VPWR VPWR _08703_ sky130_fd_sc_hd__a21oi_1
X_15525_ net471 net476 net176 net171 VGND VGND VPWR VPWR _05636_ sky130_fd_sc_hd__and4_1
XFILLER_0_155_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12737_ _02669_ _02668_ VGND VGND VPWR VPWR _02676_ sky130_fd_sc_hd__xor2_1
X_19293_ clknet_4_3_0_clock _00051_ VGND VGND VPWR VPWR ki\[4\] sky130_fd_sc_hd__dfxtp_2
XPHY_EDGE_ROW_106_Left_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18244_ _06506_ _06529_ _06532_ VGND VGND VPWR VPWR _08627_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_143_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15456_ net462 net176 VGND VGND VPWR VPWR _05560_ sky130_fd_sc_hd__nand2_1
X_12668_ _02591_ _02606_ VGND VGND VPWR VPWR _02607_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14407_ _03913_ _04403_ _04404_ VGND VGND VPWR VPWR _04406_ sky130_fd_sc_hd__nor3_1
X_11619_ net399 _00798_ _01556_ _01557_ VGND VGND VPWR VPWR _01558_ sky130_fd_sc_hd__nand4_1
X_18175_ _07972_ _07975_ _08437_ VGND VGND VPWR VPWR _08551_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_5_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15387_ _05476_ _05483_ VGND VGND VPWR VPWR _05484_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12599_ _02411_ _02413_ VGND VGND VPWR VPWR _02538_ sky130_fd_sc_hd__and2_1
XFILLER_0_108_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17126_ _07073_ _07076_ VGND VGND VPWR VPWR _07397_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14338_ _04327_ _04329_ VGND VGND VPWR VPWR _04330_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17057_ net312 _06353_ VGND VGND VPWR VPWR _07321_ sky130_fd_sc_hd__nand2_1
X_14269_ _04251_ _04253_ VGND VGND VPWR VPWR _04254_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16008_ _00563_ _01692_ _00561_ VGND VGND VPWR VPWR _06167_ sky130_fd_sc_hd__a21boi_2
XPHY_EDGE_ROW_115_Left_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17959_ _08303_ _08307_ _08312_ VGND VGND VPWR VPWR _08313_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_124_Left_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_133_Left_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11970_ _01908_ VGND VGND VPWR VPWR _01909_ sky130_fd_sc_hd__buf_2
X_10921_ _00827_ _00796_ VGND VGND VPWR VPWR _00860_ sky130_fd_sc_hd__and2b_1
X_13640_ _03596_ _03598_ _03599_ VGND VGND VPWR VPWR _03600_ sky130_fd_sc_hd__nor3_1
X_10852_ _00776_ _00790_ VGND VGND VPWR VPWR _00791_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13571_ net262 net258 _02222_ _02330_ VGND VGND VPWR VPWR _03530_ sky130_fd_sc_hd__nand4_1
X_10783_ _00694_ _00693_ VGND VGND VPWR VPWR _00722_ sky130_fd_sc_hd__and2b_1
XFILLER_0_26_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15310_ net453 net460 net177 net172 VGND VGND VPWR VPWR _05399_ sky130_fd_sc_hd__and4_1
XFILLER_0_54_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12522_ _02395_ _02459_ _02460_ VGND VGND VPWR VPWR _02461_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16290_ _06462_ _06476_ VGND VGND VPWR VPWR _06477_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15241_ net450 net171 _05228_ _05229_ VGND VGND VPWR VPWR _05323_ sky130_fd_sc_hd__o2bb2a_1
X_12453_ _02390_ _02391_ VGND VGND VPWR VPWR _02392_ sky130_fd_sc_hd__and2b_1
XFILLER_0_152_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11404_ _01337_ _01341_ _01315_ _01316_ VGND VGND VPWR VPWR _01343_ sky130_fd_sc_hd__a211o_1
X_12384_ _02321_ _02322_ VGND VGND VPWR VPWR _02323_ sky130_fd_sc_hd__or2_1
X_15172_ _05244_ _05246_ VGND VGND VPWR VPWR _05247_ sky130_fd_sc_hd__and2b_1
XFILLER_0_105_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14123_ _04067_ _04068_ _04094_ VGND VGND VPWR VPWR _04095_ sky130_fd_sc_hd__or3_2
X_11335_ _01243_ _01214_ VGND VGND VPWR VPWR _01274_ sky130_fd_sc_hd__xnor2_2
X_18931_ _01848_ _01817_ VGND VGND VPWR VPWR _09382_ sky130_fd_sc_hd__nor2_1
X_14054_ _04024_ _04025_ net408 net150 VGND VGND VPWR VPWR _04026_ sky130_fd_sc_hd__and4bb_1
X_11266_ _01169_ _01203_ _01204_ VGND VGND VPWR VPWR _01205_ sky130_fd_sc_hd__a21oi_2
X_13005_ _02916_ _02943_ _02941_ VGND VGND VPWR VPWR _02944_ sky130_fd_sc_hd__o21a_1
X_10217_ _08262_ _00155_ VGND VGND VPWR VPWR _00156_ sky130_fd_sc_hd__xnor2_1
X_18862_ _09304_ _09305_ VGND VGND VPWR VPWR _09306_ sky130_fd_sc_hd__nor2_1
X_11197_ _08097_ _00812_ VGND VGND VPWR VPWR _01136_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17813_ _08013_ _08014_ _08032_ VGND VGND VPWR VPWR _08153_ sky130_fd_sc_hd__o21a_1
X_10148_ _07393_ _08966_ VGND VGND VPWR VPWR _08977_ sky130_fd_sc_hd__xnor2_1
X_18793_ net410 net134 _04166_ _04165_ VGND VGND VPWR VPWR _09231_ sky130_fd_sc_hd__a31o_1
X_17744_ net313 _06992_ VGND VGND VPWR VPWR _08077_ sky130_fd_sc_hd__nand2_2
X_14956_ _04905_ _04904_ VGND VGND VPWR VPWR _05010_ sky130_fd_sc_hd__nor2_1
X_10079_ net338 _08207_ VGND VGND VPWR VPWR _08218_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13907_ _02770_ _03874_ VGND VGND VPWR VPWR _03875_ sky130_fd_sc_hd__nand2_1
X_17675_ net301 _07157_ _07997_ _08000_ VGND VGND VPWR VPWR _08001_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14887_ _04931_ _04933_ VGND VGND VPWR VPWR _04934_ sky130_fd_sc_hd__or2_1
X_16626_ net309 _06335_ VGND VGND VPWR VPWR _06847_ sky130_fd_sc_hd__and2_1
X_13838_ _03803_ _03802_ VGND VGND VPWR VPWR _03804_ sky130_fd_sc_hd__xnor2_1
X_19345_ clknet_4_0_0_clock _00028_ VGND VGND VPWR VPWR kd_2\[18\] sky130_fd_sc_hd__dfxtp_1
X_16557_ net293 _06345_ VGND VGND VPWR VPWR _06771_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13769_ _03734_ _03727_ VGND VGND VPWR VPWR _03735_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15508_ net466 net484 net178 net157 VGND VGND VPWR VPWR _05617_ sky130_fd_sc_hd__and4_1
X_19276_ clknet_4_6_0_clock _00072_ VGND VGND VPWR VPWR kp\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16488_ _06686_ _06691_ _06694_ VGND VGND VPWR VPWR _06695_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_45_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18227_ _08596_ _08600_ _08601_ _08607_ VGND VGND VPWR VPWR _08608_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_115_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15439_ _05539_ _05540_ VGND VGND VPWR VPWR _05541_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18158_ _07046_ _08520_ _07044_ VGND VGND VPWR VPWR _08532_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_13_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17109_ _07375_ _07377_ VGND VGND VPWR VPWR _07378_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_13_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18089_ _08446_ _08447_ VGND VGND VPWR VPWR _08456_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09931_ _04621_ _06579_ _04533_ VGND VGND VPWR VPWR _06590_ sky130_fd_sc_hd__or3_4
XFILLER_0_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09862_ _05743_ _05809_ VGND VGND VPWR VPWR _05831_ sky130_fd_sc_hd__nand2_1
X_09793_ _05061_ VGND VGND VPWR VPWR _05072_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11120_ _01057_ _01052_ _01058_ VGND VGND VPWR VPWR _01059_ sky130_fd_sc_hd__nand3_1
XFILLER_0_101_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11051_ _00938_ _00937_ _00924_ VGND VGND VPWR VPWR _00990_ sky130_fd_sc_hd__a21oi_1
X_10002_ net403 net398 kp\[3\] _05072_ VGND VGND VPWR VPWR _07371_ sky130_fd_sc_hd__o31a_1
X_14810_ _04718_ _04792_ _04827_ VGND VGND VPWR VPWR _04849_ sky130_fd_sc_hd__a21oi_1
X_15790_ _05893_ _05913_ _05925_ _05926_ VGND VGND VPWR VPWR _05927_ sky130_fd_sc_hd__and4bb_1
X_14741_ _04751_ _04772_ VGND VGND VPWR VPWR _04773_ sky130_fd_sc_hd__xnor2_1
X_11953_ _01890_ _01891_ VGND VGND VPWR VPWR _01892_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17460_ _07760_ _07763_ VGND VGND VPWR VPWR _07764_ sky130_fd_sc_hd__nand2_1
X_10904_ _00833_ _00839_ VGND VGND VPWR VPWR _00843_ sky130_fd_sc_hd__xnor2_1
X_14672_ _04623_ _04625_ VGND VGND VPWR VPWR _04697_ sky130_fd_sc_hd__nor2_1
X_11884_ _01821_ _01822_ VGND VGND VPWR VPWR _01823_ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16411_ _06594_ _06609_ VGND VGND VPWR VPWR _06610_ sky130_fd_sc_hd__and2_1
XFILLER_0_157_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13623_ _03559_ _03581_ VGND VGND VPWR VPWR _03582_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17391_ _07597_ _07674_ _07686_ VGND VGND VPWR VPWR _07688_ sky130_fd_sc_hd__nor3_1
X_10835_ _00772_ _00773_ VGND VGND VPWR VPWR _00774_ sky130_fd_sc_hd__and2b_1
XFILLER_0_104_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19130_ net506 net552 net496 _09556_ VGND VGND VPWR VPWR _00120_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16342_ _06532_ _06533_ VGND VGND VPWR VPWR _06534_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13554_ net244 net240 _02544_ _02640_ VGND VGND VPWR VPWR _03513_ sky130_fd_sc_hd__and4_1
X_10766_ _00702_ _00704_ VGND VGND VPWR VPWR _00705_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12505_ _02440_ _02443_ VGND VGND VPWR VPWR _02444_ sky130_fd_sc_hd__or2_1
X_19061_ net504 net549 net493 VGND VGND VPWR VPWR _09513_ sky130_fd_sc_hd__o21ai_1
X_16273_ _06455_ _06457_ VGND VGND VPWR VPWR _06459_ sky130_fd_sc_hd__or2b_1
X_13485_ _03442_ _03443_ VGND VGND VPWR VPWR _03444_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10697_ _00634_ _00635_ VGND VGND VPWR VPWR _00636_ sky130_fd_sc_hd__xnor2_2
X_18012_ _08368_ _08370_ VGND VGND VPWR VPWR _08371_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15224_ prev_d_error\[3\] net157 net153 net477 VGND VGND VPWR VPWR _05305_ sky130_fd_sc_hd__a22oi_1
X_12436_ _02370_ _02374_ VGND VGND VPWR VPWR _02375_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15155_ net453 net167 net162 net459 VGND VGND VPWR VPWR _05229_ sky130_fd_sc_hd__a22oi_1
X_12367_ _02279_ _02304_ _02206_ _02305_ VGND VGND VPWR VPWR _02306_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_105_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14106_ _04076_ _04077_ VGND VGND VPWR VPWR _04078_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11318_ _00439_ _06579_ _08163_ VGND VGND VPWR VPWR _01257_ sky130_fd_sc_hd__or3_1
X_12298_ _02189_ _02201_ _02236_ VGND VGND VPWR VPWR _02237_ sky130_fd_sc_hd__a21oi_1
X_15086_ _05148_ _05152_ VGND VGND VPWR VPWR _05153_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14037_ _03972_ _03974_ _04008_ VGND VGND VPWR VPWR _04009_ sky130_fd_sc_hd__o21ai_1
X_18914_ _01929_ _09363_ VGND VGND VPWR VPWR _09364_ sky130_fd_sc_hd__xnor2_1
X_11249_ _01059_ _01172_ _01186_ VGND VGND VPWR VPWR _01188_ sky130_fd_sc_hd__nand3_1
XFILLER_0_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18845_ net201 _01817_ VGND VGND VPWR VPWR _09288_ sky130_fd_sc_hd__nand2_1
X_18776_ _08998_ _09007_ _09211_ VGND VGND VPWR VPWR _09212_ sky130_fd_sc_hd__o21bai_1
X_15988_ _06142_ _06144_ VGND VGND VPWR VPWR _06145_ sky130_fd_sc_hd__xnor2_4
X_17727_ net327 _06720_ _08055_ _08056_ VGND VGND VPWR VPWR _08058_ sky130_fd_sc_hd__a22o_1
X_14939_ _04881_ _04882_ VGND VGND VPWR VPWR _04991_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17658_ net327 _06619_ _07980_ _07981_ VGND VGND VPWR VPWR _07982_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16609_ _06826_ _06827_ VGND VGND VPWR VPWR _06828_ sky130_fd_sc_hd__and2b_1
XFILLER_0_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17589_ _07852_ _07904_ _07903_ VGND VGND VPWR VPWR _07906_ sky130_fd_sc_hd__a21oi_1
X_19328_ clknet_4_3_0_clock _00029_ VGND VGND VPWR VPWR kd_2\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19259_ clknet_4_10_0_clock _00141_ VGND VGND VPWR VPWR prev_d_error\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09914_ _06128_ _06271_ _06392_ VGND VGND VPWR VPWR _06403_ sky130_fd_sc_hd__o21a_1
X_09845_ _05545_ _05622_ VGND VGND VPWR VPWR _05644_ sky130_fd_sc_hd__xor2_2
X_09776_ _04874_ VGND VGND VPWR VPWR _04885_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_68_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10620_ _00465_ _00558_ VGND VGND VPWR VPWR _00559_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10551_ _00485_ _00489_ VGND VGND VPWR VPWR _00490_ sky130_fd_sc_hd__or2b_1
XFILLER_0_134_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13270_ _03221_ _03129_ VGND VGND VPWR VPWR _03223_ sky130_fd_sc_hd__nor2_1
X_10482_ net336 _00397_ _00420_ _00418_ VGND VGND VPWR VPWR _00421_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_122_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12221_ _01979_ _02003_ _02159_ VGND VGND VPWR VPWR _02160_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12152_ _02090_ VGND VGND VPWR VPWR _02091_ sky130_fd_sc_hd__buf_2
XFILLER_0_102_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11103_ _01039_ _01040_ _01041_ VGND VGND VPWR VPWR _01042_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16960_ _07212_ _07213_ VGND VGND VPWR VPWR _07214_ sky130_fd_sc_hd__nor2_1
X_12083_ _01923_ _01921_ VGND VGND VPWR VPWR _02022_ sky130_fd_sc_hd__xnor2_1
X_15911_ _06057_ _06059_ VGND VGND VPWR VPWR _06060_ sky130_fd_sc_hd__nand2_1
X_11034_ _00967_ _00962_ VGND VGND VPWR VPWR _00973_ sky130_fd_sc_hd__and2b_1
X_16891_ _07133_ _07136_ _07137_ VGND VGND VPWR VPWR _07138_ sky130_fd_sc_hd__o21a_1
X_18630_ _08908_ _09050_ _08964_ VGND VGND VPWR VPWR _09051_ sky130_fd_sc_hd__mux2_1
X_15842_ _04473_ _04472_ VGND VGND VPWR VPWR _05984_ sky130_fd_sc_hd__and2b_1
X_18561_ _08974_ _08744_ _08882_ VGND VGND VPWR VPWR _08975_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15773_ _05887_ _05885_ VGND VGND VPWR VPWR _05909_ sky130_fd_sc_hd__xnor2_1
X_12985_ net204 _02747_ VGND VGND VPWR VPWR _02924_ sky130_fd_sc_hd__nand2_1
X_17512_ net295 _07156_ VGND VGND VPWR VPWR _07821_ sky130_fd_sc_hd__nand2_1
X_14724_ net426 net174 _04558_ VGND VGND VPWR VPWR _04755_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11936_ _01874_ VGND VGND VPWR VPWR _01875_ sky130_fd_sc_hd__buf_2
X_18492_ _06266_ _08761_ VGND VGND VPWR VPWR _08899_ sky130_fd_sc_hd__or2_2
XFILLER_0_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17443_ _07677_ _07738_ _07743_ VGND VGND VPWR VPWR _07746_ sky130_fd_sc_hd__and3_1
X_14655_ _04677_ _04678_ VGND VGND VPWR VPWR _04679_ sky130_fd_sc_hd__or2b_1
XFILLER_0_39_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11867_ _01745_ _01805_ VGND VGND VPWR VPWR _01806_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13606_ _03560_ _03563_ VGND VGND VPWR VPWR _03565_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17374_ _07565_ _07572_ _07669_ VGND VGND VPWR VPWR _07670_ sky130_fd_sc_hd__a21o_1
X_10818_ _00755_ _00756_ VGND VGND VPWR VPWR _00757_ sky130_fd_sc_hd__nand2_1
X_14586_ _04596_ _04602_ VGND VGND VPWR VPWR _04603_ sky130_fd_sc_hd__nor2_1
X_11798_ _01707_ _01734_ _01735_ _01736_ VGND VGND VPWR VPWR _01737_ sky130_fd_sc_hd__o211ai_2
X_19113_ _09536_ _05677_ _09545_ net488 VGND VGND VPWR VPWR _00112_ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16325_ _06419_ _06514_ VGND VGND VPWR VPWR _06516_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13537_ _03458_ _03494_ _03495_ VGND VGND VPWR VPWR _03496_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_153_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10749_ net365 _08207_ _00687_ _00685_ VGND VGND VPWR VPWR _00688_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19044_ _09498_ _09500_ net493 VGND VGND VPWR VPWR _00082_ sky130_fd_sc_hd__o21a_1
XFILLER_0_113_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16256_ net279 _06410_ _06404_ net275 VGND VGND VPWR VPWR _06440_ sky130_fd_sc_hd__a22oi_1
X_13468_ _03422_ _03426_ VGND VGND VPWR VPWR _03427_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15207_ _05265_ _05284_ net112 _05285_ VGND VGND VPWR VPWR _05286_ sky130_fd_sc_hd__a211oi_1
X_12419_ _02351_ _02357_ VGND VGND VPWR VPWR _02358_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16187_ _06363_ VGND VGND VPWR VPWR _06364_ sky130_fd_sc_hd__buf_2
XFILLER_0_23_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13399_ _03348_ _03353_ VGND VGND VPWR VPWR _03354_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15138_ _05208_ _05209_ net479 net143 VGND VGND VPWR VPWR _05210_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_49_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15069_ _05111_ _05120_ _05122_ VGND VGND VPWR VPWR _05134_ sky130_fd_sc_hd__nand3_1
XFILLER_0_49_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_155_Right_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09630_ net21 net33 net32 net79 VGND VGND VPWR VPWR _03336_ sky130_fd_sc_hd__or4_2
X_18828_ _09227_ _09268_ VGND VGND VPWR VPWR _09269_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_156_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18759_ _09072_ _09085_ VGND VGND VPWR VPWR _09193_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout410 prev_d_error\[17\] VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__clkbuf_4
Xfanout421 net424 VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout432 net433 VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__clkbuf_4
Xfanout443 net445 VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__buf_2
Xfanout454 net455 VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__clkbuf_4
Xfanout465 net468 VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__buf_2
Xfanout476 net477 VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__buf_2
X_09828_ _05347_ _05446_ VGND VGND VPWR VPWR _05457_ sky130_fd_sc_hd__xnor2_1
Xfanout487 net497 VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_122_Right_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout498 net1 VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__clkbuf_4
X_09759_ net63 net5 VGND VGND VPWR VPWR _04698_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_69_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12770_ _02696_ _02707_ _02708_ VGND VGND VPWR VPWR _02709_ sky130_fd_sc_hd__and3_2
XFILLER_0_68_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11721_ _01547_ _01577_ VGND VGND VPWR VPWR _01660_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14440_ _04016_ net170 VGND VGND VPWR VPWR _04442_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11652_ _01588_ _01590_ _01518_ VGND VGND VPWR VPWR _01591_ sky130_fd_sc_hd__a21oi_1
X_10603_ _00540_ _00536_ VGND VGND VPWR VPWR _00542_ sky130_fd_sc_hd__and2b_1
XFILLER_0_80_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14371_ _04274_ _04276_ VGND VGND VPWR VPWR _04366_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11583_ _01520_ _01516_ _01519_ VGND VGND VPWR VPWR _01522_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16110_ _01714_ _00600_ VGND VGND VPWR VPWR _06279_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13322_ net248 _02090_ _03274_ VGND VGND VPWR VPWR _03275_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10534_ _00471_ _00472_ VGND VGND VPWR VPWR _00473_ sky130_fd_sc_hd__xor2_4
X_17090_ _07354_ _07356_ VGND VGND VPWR VPWR _07357_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_10_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16041_ _06202_ net349 _08889_ VGND VGND VPWR VPWR _06203_ sky130_fd_sc_hd__mux2_1
X_13253_ _03204_ _03205_ VGND VGND VPWR VPWR _03206_ sky130_fd_sc_hd__xnor2_1
X_10465_ _00327_ _00403_ VGND VGND VPWR VPWR _00404_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12204_ _01962_ _01964_ VGND VGND VPWR VPWR _02143_ sky130_fd_sc_hd__and2b_1
XFILLER_0_110_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13184_ _03130_ _03133_ _03136_ VGND VGND VPWR VPWR _03137_ sky130_fd_sc_hd__a21o_1
X_10396_ _00332_ _00333_ _00334_ VGND VGND VPWR VPWR _00335_ sky130_fd_sc_hd__o21bai_1
X_12135_ _01915_ _01917_ VGND VGND VPWR VPWR _02074_ sky130_fd_sc_hd__or2_1
X_17992_ _08337_ _08342_ _08341_ VGND VGND VPWR VPWR _08349_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16943_ net297 _06620_ _07193_ VGND VGND VPWR VPWR _07196_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12066_ _02003_ _02004_ VGND VGND VPWR VPWR _02005_ sky130_fd_sc_hd__nor2_1
X_11017_ _00868_ _00955_ VGND VGND VPWR VPWR _00956_ sky130_fd_sc_hd__nor2_1
X_16874_ net320 _06316_ _06318_ _07119_ VGND VGND VPWR VPWR _07120_ sky130_fd_sc_hd__nand4_2
X_15825_ _04894_ _05965_ VGND VGND VPWR VPWR _05966_ sky130_fd_sc_hd__nand2_1
X_18613_ _09024_ _09031_ VGND VGND VPWR VPWR _09033_ sky130_fd_sc_hd__xor2_1
XFILLER_0_126_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15756_ _05788_ _05821_ VGND VGND VPWR VPWR _05890_ sky130_fd_sc_hd__xnor2_1
X_18544_ _08923_ _08931_ _08940_ _08956_ VGND VGND VPWR VPWR _08957_ sky130_fd_sc_hd__nor4_1
XFILLER_0_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12968_ _02893_ _02906_ VGND VGND VPWR VPWR _02907_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14707_ _04710_ _04713_ _04735_ VGND VGND VPWR VPWR _04736_ sky130_fd_sc_hd__a21o_1
XFILLER_0_157_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18475_ _08880_ VGND VGND VPWR VPWR _08881_ sky130_fd_sc_hd__buf_6
X_11919_ _01705_ _01737_ VGND VGND VPWR VPWR _01858_ sky130_fd_sc_hd__nand2_2
X_15687_ _05752_ _05799_ VGND VGND VPWR VPWR _05814_ sky130_fd_sc_hd__nand2_1
XFILLER_0_142_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12899_ kd_1\[18\] _02748_ _02757_ VGND VGND VPWR VPWR _02838_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17426_ _07724_ _07726_ VGND VGND VPWR VPWR _07727_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_157_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14638_ _04657_ _04659_ VGND VGND VPWR VPWR _04660_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17357_ _07638_ _07650_ VGND VGND VPWR VPWR _07651_ sky130_fd_sc_hd__xor2_1
X_14569_ _04583_ _04582_ VGND VGND VPWR VPWR _04584_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16308_ net289 _06389_ _06320_ VGND VGND VPWR VPWR _06497_ sky130_fd_sc_hd__nand3_1
XFILLER_0_126_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17288_ _07555_ _07562_ VGND VGND VPWR VPWR _07575_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19027_ net563 net90 VGND VGND VPWR VPWR _09487_ sky130_fd_sc_hd__and2_1
X_16239_ net280 _06386_ _06346_ net275 VGND VGND VPWR VPWR _06421_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09613_ net51 _03102_ _03135_ net190 VGND VGND VPWR VPWR _00030_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10250_ _07778_ _00163_ VGND VGND VPWR VPWR _00189_ sky130_fd_sc_hd__xnor2_1
X_10181_ _07899_ _09285_ _09329_ VGND VGND VPWR VPWR _09340_ sky130_fd_sc_hd__or3b_1
Xfanout240 net241 VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__buf_2
XFILLER_0_100_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout251 net253 VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__buf_2
Xfanout262 kd_1\[2\] VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__clkbuf_4
X_13940_ _03910_ _03894_ VGND VGND VPWR VPWR _03911_ sky130_fd_sc_hd__xor2_2
Xfanout273 ki\[17\] VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__clkbuf_4
Xfanout284 ki\[14\] VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__buf_2
Xfanout295 ki\[10\] VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__clkbuf_4
X_13871_ _03823_ _03835_ _03836_ VGND VGND VPWR VPWR _03837_ sky130_fd_sc_hd__a21o_1
X_15610_ _05667_ _05665_ _05634_ VGND VGND VPWR VPWR _05729_ sky130_fd_sc_hd__a21oi_1
X_12822_ _02680_ _02731_ VGND VGND VPWR VPWR _02761_ sky130_fd_sc_hd__xor2_1
X_16590_ net288 _06431_ _06434_ VGND VGND VPWR VPWR _06807_ sky130_fd_sc_hd__and3_2
X_15541_ _05650_ _05641_ _05648_ VGND VGND VPWR VPWR _05653_ sky130_fd_sc_hd__nand3_1
X_12753_ _02690_ _02691_ VGND VGND VPWR VPWR _02692_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11704_ _01636_ _01639_ _01642_ VGND VGND VPWR VPWR _01643_ sky130_fd_sc_hd__a21oi_1
X_18260_ _06519_ _06522_ _08642_ VGND VGND VPWR VPWR _08644_ sky130_fd_sc_hd__and3_1
X_15472_ _05572_ _05576_ VGND VGND VPWR VPWR _05577_ sky130_fd_sc_hd__and2b_1
X_12684_ _02620_ _02622_ VGND VGND VPWR VPWR _02623_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17211_ net332 _06463_ _06465_ VGND VGND VPWR VPWR _07490_ sky130_fd_sc_hd__and3_1
X_14423_ _04330_ _04422_ VGND VGND VPWR VPWR _04424_ sky130_fd_sc_hd__or2_1
X_11635_ _01565_ _01567_ VGND VGND VPWR VPWR _01574_ sky130_fd_sc_hd__nand2_1
X_18191_ _08552_ _08566_ _08567_ VGND VGND VPWR VPWR _08568_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17142_ _07104_ _07413_ VGND VGND VPWR VPWR _07414_ sky130_fd_sc_hd__nand2_1
X_14354_ net407 net165 _04264_ _04265_ VGND VGND VPWR VPWR _04348_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_64_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11566_ _01481_ _01504_ VGND VGND VPWR VPWR _01505_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13305_ _03219_ _03228_ VGND VGND VPWR VPWR _03258_ sky130_fd_sc_hd__and2_1
X_17073_ net304 _06402_ _07337_ VGND VGND VPWR VPWR _07339_ sky130_fd_sc_hd__and3_1
X_10517_ _00431_ _00454_ VGND VGND VPWR VPWR _00456_ sky130_fd_sc_hd__and2_1
X_14285_ _04003_ _04271_ VGND VGND VPWR VPWR _04272_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11497_ net400 _09577_ _01434_ _01435_ VGND VGND VPWR VPWR _01436_ sky130_fd_sc_hd__a31o_1
XFILLER_0_33_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16024_ _06180_ _06184_ VGND VGND VPWR VPWR _06185_ sky130_fd_sc_hd__xnor2_1
X_13236_ _03187_ _03188_ VGND VGND VPWR VPWR _03189_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10448_ _00381_ _00386_ VGND VGND VPWR VPWR _00387_ sky130_fd_sc_hd__or2b_1
XFILLER_0_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13167_ _03115_ _03117_ VGND VGND VPWR VPWR _03118_ sky130_fd_sc_hd__and2_1
X_10379_ _00315_ _00317_ VGND VGND VPWR VPWR _00318_ sky130_fd_sc_hd__xnor2_1
X_12118_ _02054_ _02056_ VGND VGND VPWR VPWR _02057_ sky130_fd_sc_hd__or2b_1
X_13098_ _03040_ _03041_ VGND VGND VPWR VPWR _03042_ sky130_fd_sc_hd__nor2_1
X_17975_ _08324_ _08327_ _08330_ VGND VGND VPWR VPWR _08331_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16926_ net282 _06993_ _07176_ VGND VGND VPWR VPWR _07177_ sky130_fd_sc_hd__nand3_1
X_12049_ net223 _01931_ VGND VGND VPWR VPWR _01988_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16857_ net271 _07095_ _07100_ _07098_ VGND VGND VPWR VPWR _07101_ sky130_fd_sc_hd__a31o_1
X_15808_ _05613_ _05544_ _05614_ _05946_ VGND VGND VPWR VPWR _05947_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16788_ _06541_ _07023_ _07024_ VGND VGND VPWR VPWR _07025_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15739_ net469 net196 net192 net473 VGND VGND VPWR VPWR _05871_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18527_ _08810_ _08936_ VGND VGND VPWR VPWR _08938_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18458_ _08861_ VGND VGND VPWR VPWR _08862_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17409_ _07699_ _07707_ VGND VGND VPWR VPWR _07708_ sky130_fd_sc_hd__xor2_1
XFILLER_0_8_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18389_ _06158_ _06141_ VGND VGND VPWR VPWR _08786_ sky130_fd_sc_hd__or2b_1
XFILLER_0_145_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold37 net86 VGND VGND VPWR VPWR net544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 i_error\[1\] VGND VGND VPWR VPWR net555 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11420_ _01053_ _01358_ VGND VGND VPWR VPWR _01359_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11351_ _01288_ _01284_ VGND VGND VPWR VPWR _01290_ sky130_fd_sc_hd__xor2_1
XFILLER_0_22_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10302_ _04280_ _00238_ _00239_ _00240_ VGND VGND VPWR VPWR _00241_ sky130_fd_sc_hd__a31o_1
X_14070_ _04039_ _04040_ _04015_ _04021_ VGND VGND VPWR VPWR _04042_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11282_ net370 _00798_ VGND VGND VPWR VPWR _01221_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13021_ _02782_ _02791_ VGND VGND VPWR VPWR _02960_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10233_ _08053_ _00170_ _00165_ _00169_ VGND VGND VPWR VPWR _00172_ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10164_ _05589_ _05006_ _09142_ VGND VGND VPWR VPWR _09153_ sky130_fd_sc_hd__a21o_1
XFILLER_0_100_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10095_ _08152_ _08361_ _08383_ VGND VGND VPWR VPWR _08394_ sky130_fd_sc_hd__o21a_1
X_14972_ _05005_ _05008_ VGND VGND VPWR VPWR _05027_ sky130_fd_sc_hd__nor2_1
X_17760_ _08092_ _08093_ VGND VGND VPWR VPWR _08094_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13923_ net465 net485 net116 VGND VGND VPWR VPWR _03893_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16711_ net317 _06316_ _06318_ VGND VGND VPWR VPWR _06940_ sky130_fd_sc_hd__and3_1
X_17691_ net298 _07570_ VGND VGND VPWR VPWR _08018_ sky130_fd_sc_hd__nand2_1
X_16642_ _06862_ _06863_ VGND VGND VPWR VPWR _06864_ sky130_fd_sc_hd__and2b_1
X_13854_ _03818_ _03819_ VGND VGND VPWR VPWR _03820_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12805_ prev_error\[2\] _00612_ VGND VGND VPWR VPWR _02744_ sky130_fd_sc_hd__xor2_4
X_16573_ _06784_ _06786_ VGND VGND VPWR VPWR _06789_ sky130_fd_sc_hd__and2b_1
X_13785_ _03746_ _03748_ _03747_ VGND VGND VPWR VPWR _03751_ sky130_fd_sc_hd__o21a_1
X_10997_ _00931_ _00935_ VGND VGND VPWR VPWR _00936_ sky130_fd_sc_hd__nand2_1
X_15524_ _05586_ _05602_ _05601_ VGND VGND VPWR VPWR _05635_ sky130_fd_sc_hd__a21o_1
X_18312_ net273 _06386_ _08635_ _08700_ VGND VGND VPWR VPWR _08701_ sky130_fd_sc_hd__a31o_1
X_12736_ _02672_ _02674_ VGND VGND VPWR VPWR _02675_ sky130_fd_sc_hd__nor2_1
X_19292_ clknet_4_8_0_clock _00050_ VGND VGND VPWR VPWR ki\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18243_ _06588_ _06487_ VGND VGND VPWR VPWR _08626_ sky130_fd_sc_hd__or2b_1
X_15455_ _05214_ _05557_ _05558_ VGND VGND VPWR VPWR _05559_ sky130_fd_sc_hd__a21oi_2
X_12667_ _02591_ _02604_ _02605_ VGND VGND VPWR VPWR _02606_ sky130_fd_sc_hd__nand3_2
XFILLER_0_72_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14406_ _03913_ _04403_ _04404_ VGND VGND VPWR VPWR _04405_ sky130_fd_sc_hd__o21a_1
X_11618_ net394 _00514_ _00612_ net390 VGND VGND VPWR VPWR _01557_ sky130_fd_sc_hd__a22o_1
X_18174_ _07972_ _07975_ _08437_ VGND VGND VPWR VPWR _08550_ sky130_fd_sc_hd__or3b_1
XFILLER_0_108_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15386_ _05475_ _05471_ _05473_ VGND VGND VPWR VPWR _05483_ sky130_fd_sc_hd__or3_1
X_12598_ net209 _02224_ _02536_ VGND VGND VPWR VPWR _02537_ sky130_fd_sc_hd__and3_1
XFILLER_0_80_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17125_ _07359_ _07361_ _07395_ VGND VGND VPWR VPWR _07396_ sky130_fd_sc_hd__a21bo_1
X_14337_ _04260_ _04328_ VGND VGND VPWR VPWR _04329_ sky130_fd_sc_hd__nor2_1
X_11549_ net394 _00406_ _00407_ VGND VGND VPWR VPWR _01488_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17056_ _07122_ _07318_ _07317_ VGND VGND VPWR VPWR _07320_ sky130_fd_sc_hd__a21oi_1
X_14268_ _04230_ _04252_ VGND VGND VPWR VPWR _04253_ sky130_fd_sc_hd__nand2_1
X_16007_ _06134_ _06163_ _06165_ VGND VGND VPWR VPWR _06166_ sky130_fd_sc_hd__or3_1
X_13219_ _03167_ _03171_ VGND VGND VPWR VPWR _03172_ sky130_fd_sc_hd__and2_1
X_14199_ _04175_ _04176_ VGND VGND VPWR VPWR _04177_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17958_ _08304_ _08305_ VGND VGND VPWR VPWR _08312_ sky130_fd_sc_hd__nor2_1
X_16909_ net278 _07095_ VGND VGND VPWR VPWR _07158_ sky130_fd_sc_hd__nand2_2
X_17889_ net331 _06801_ _07156_ net314 VGND VGND VPWR VPWR _08236_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10920_ _00761_ _00858_ VGND VGND VPWR VPWR _00859_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10851_ _00768_ _00774_ _00775_ VGND VGND VPWR VPWR _00790_ sky130_fd_sc_hd__or3_1
XFILLER_0_39_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13570_ _03468_ _03528_ VGND VGND VPWR VPWR _03529_ sky130_fd_sc_hd__nor2_1
X_10782_ _00629_ _00647_ VGND VGND VPWR VPWR _00721_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_136_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12521_ _02360_ _02458_ VGND VGND VPWR VPWR _02460_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15240_ _05310_ _05313_ _05311_ VGND VGND VPWR VPWR _05322_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_152_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12452_ _02376_ _02361_ VGND VGND VPWR VPWR _02391_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_136_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11403_ _01315_ _01316_ _01337_ _01341_ VGND VGND VPWR VPWR _01342_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_140_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15171_ _05245_ _05142_ VGND VGND VPWR VPWR _05246_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12383_ _02320_ _02315_ VGND VGND VPWR VPWR _02322_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14122_ _04092_ _04093_ VGND VGND VPWR VPWR _04094_ sky130_fd_sc_hd__or2_1
X_11334_ _01246_ _01271_ VGND VGND VPWR VPWR _01273_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_132_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14053_ net412 net144 net138 net418 VGND VGND VPWR VPWR _04025_ sky130_fd_sc_hd__a22oi_1
X_18930_ _09299_ _09380_ VGND VGND VPWR VPWR _09381_ sky130_fd_sc_hd__or2_1
X_11265_ _01198_ _01202_ net109 _01170_ VGND VGND VPWR VPWR _01204_ sky130_fd_sc_hd__a211oi_1
X_13004_ _02941_ _02942_ VGND VGND VPWR VPWR _02943_ sky130_fd_sc_hd__nand2_1
X_10216_ _08350_ _08339_ VGND VGND VPWR VPWR _00155_ sky130_fd_sc_hd__nor2_1
X_18861_ _09303_ _09281_ VGND VGND VPWR VPWR _09305_ sky130_fd_sc_hd__and2b_1
X_11196_ _01044_ _01129_ VGND VGND VPWR VPWR _01135_ sky130_fd_sc_hd__xnor2_1
X_17812_ _08137_ _08143_ VGND VGND VPWR VPWR _08151_ sky130_fd_sc_hd__or2_1
X_10147_ _08944_ _08955_ VGND VGND VPWR VPWR _08966_ sky130_fd_sc_hd__nor2_1
X_18792_ prev_d_error\[18\] _04961_ VGND VGND VPWR VPWR _09229_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14955_ _05005_ _05007_ _05008_ VGND VGND VPWR VPWR _05009_ sky130_fd_sc_hd__o21ba_1
X_17743_ _08072_ _08074_ VGND VGND VPWR VPWR _08076_ sky130_fd_sc_hd__xnor2_1
X_10078_ _08196_ VGND VGND VPWR VPWR _08207_ sky130_fd_sc_hd__clkbuf_4
X_13906_ _02675_ _02769_ VGND VGND VPWR VPWR _03874_ sky130_fd_sc_hd__or2_1
X_14886_ _04931_ _04932_ net422 net184 VGND VGND VPWR VPWR _04933_ sky130_fd_sc_hd__and4b_1
X_17674_ _07907_ _07999_ VGND VGND VPWR VPWR _08000_ sky130_fd_sc_hd__nor2_1
X_13837_ _03770_ _03789_ VGND VGND VPWR VPWR _03803_ sky130_fd_sc_hd__nor2_1
X_16625_ net306 _06335_ _06310_ net309 VGND VGND VPWR VPWR _06846_ sky130_fd_sc_hd__a22oi_2
X_16556_ _06767_ _06769_ VGND VGND VPWR VPWR _06770_ sky130_fd_sc_hd__xnor2_1
X_19344_ clknet_4_0_0_clock _00027_ VGND VGND VPWR VPWR kd_2\[17\] sky130_fd_sc_hd__dfxtp_1
X_13768_ _03676_ _03722_ VGND VGND VPWR VPWR _03734_ sky130_fd_sc_hd__nor2_1
X_12719_ _02657_ VGND VGND VPWR VPWR _02658_ sky130_fd_sc_hd__inv_2
X_15507_ _05608_ _05615_ VGND VGND VPWR VPWR _05616_ sky130_fd_sc_hd__or2_1
X_16487_ _06692_ _06693_ VGND VGND VPWR VPWR _06694_ sky130_fd_sc_hd__and2_1
X_19275_ clknet_4_6_0_clock _00071_ VGND VGND VPWR VPWR kp\[5\] sky130_fd_sc_hd__dfxtp_1
X_13699_ _03631_ _03664_ _03662_ VGND VGND VPWR VPWR _03665_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_128_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15438_ _05538_ _05529_ _05537_ VGND VGND VPWR VPWR _05540_ sky130_fd_sc_hd__or3_1
X_18226_ i_error\[12\] _08606_ VGND VGND VPWR VPWR _08607_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_155_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15369_ _05458_ _05461_ _05463_ VGND VGND VPWR VPWR _05464_ sky130_fd_sc_hd__o21ai_2
X_18157_ _06934_ _08530_ VGND VGND VPWR VPWR _08531_ sky130_fd_sc_hd__and2_1
X_17108_ _07089_ _07376_ VGND VGND VPWR VPWR _07377_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18088_ _07351_ _08453_ _08452_ _08451_ VGND VGND VPWR VPWR _08455_ sky130_fd_sc_hd__a211o_1
X_09930_ _04423_ _04500_ _04643_ VGND VGND VPWR VPWR _06579_ sky130_fd_sc_hd__a21oi_4
X_17039_ _07298_ _07299_ _07300_ VGND VGND VPWR VPWR _07301_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09861_ _05743_ _05809_ VGND VGND VPWR VPWR _05820_ sky130_fd_sc_hd__or2_1
X_09792_ _05039_ _05050_ VGND VGND VPWR VPWR _05061_ sky130_fd_sc_hd__nand2_4
XFILLER_0_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11050_ _00938_ _00924_ _00937_ VGND VGND VPWR VPWR _00989_ sky130_fd_sc_hd__and3_1
X_10001_ _07272_ _07349_ VGND VGND VPWR VPWR _07360_ sky130_fd_sc_hd__or2_2
X_14740_ _04752_ _04771_ _04769_ VGND VGND VPWR VPWR _04772_ sky130_fd_sc_hd__a21oi_1
X_11952_ _01889_ _01867_ _01879_ VGND VGND VPWR VPWR _01891_ sky130_fd_sc_hd__nor3_1
XFILLER_0_59_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10903_ _00676_ _00764_ _00766_ VGND VGND VPWR VPWR _00842_ sky130_fd_sc_hd__nand3_1
X_14671_ _04693_ _04695_ VGND VGND VPWR VPWR _04696_ sky130_fd_sc_hd__nand2_1
X_11883_ _01804_ _01820_ VGND VGND VPWR VPWR _01822_ sky130_fd_sc_hd__and2_1
X_16410_ _06372_ _06592_ _06593_ VGND VGND VPWR VPWR _06609_ sky130_fd_sc_hd__or3_1
X_13622_ net248 _02545_ VGND VGND VPWR VPWR _03581_ sky130_fd_sc_hd__nand2_1
X_17390_ _07597_ _07674_ _07686_ VGND VGND VPWR VPWR _07687_ sky130_fd_sc_hd__o21a_1
X_10834_ _00767_ _00763_ VGND VGND VPWR VPWR _00773_ sky130_fd_sc_hd__xnor2_1
X_16341_ _06530_ _06531_ VGND VGND VPWR VPWR _06533_ sky130_fd_sc_hd__nand2_1
X_13553_ net243 _02544_ _02640_ net240 VGND VGND VPWR VPWR _03512_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10765_ net359 _00244_ _00503_ _00703_ VGND VGND VPWR VPWR _00704_ sky130_fd_sc_hd__a31o_1
XFILLER_0_82_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12504_ _02270_ _02439_ _02437_ VGND VGND VPWR VPWR _02443_ sky130_fd_sc_hd__nor3_1
X_19060_ net522 _09484_ VGND VGND VPWR VPWR _09512_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16272_ _06454_ _06456_ VGND VGND VPWR VPWR _06457_ sky130_fd_sc_hd__and2_1
X_13484_ _03402_ _03405_ VGND VGND VPWR VPWR _03443_ sky130_fd_sc_hd__xnor2_1
X_10696_ net384 _05413_ VGND VGND VPWR VPWR _00635_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15223_ prev_d_error\[3\] net477 net157 net153 VGND VGND VPWR VPWR _05304_ sky130_fd_sc_hd__and4_1
X_18011_ _08360_ _08369_ VGND VGND VPWR VPWR _08370_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12435_ net234 _01808_ _02371_ _02373_ VGND VGND VPWR VPWR _02374_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_35_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15154_ net453 net459 net167 net162 VGND VGND VPWR VPWR _05228_ sky130_fd_sc_hd__and4_1
X_12366_ _02203_ _02205_ VGND VGND VPWR VPWR _02305_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_136_Right_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14105_ _03923_ _03939_ _03940_ VGND VGND VPWR VPWR _04077_ sky130_fd_sc_hd__o21ba_1
X_11317_ _01177_ _01255_ VGND VGND VPWR VPWR _01256_ sky130_fd_sc_hd__xor2_1
X_15085_ _05150_ _05151_ VGND VGND VPWR VPWR _05152_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12297_ _02101_ _02235_ VGND VGND VPWR VPWR _02236_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14036_ _04006_ _04007_ VGND VGND VPWR VPWR _04008_ sky130_fd_sc_hd__nor2_1
X_18913_ _01982_ _09319_ _01979_ VGND VGND VPWR VPWR _09363_ sky130_fd_sc_hd__o21ba_1
X_11248_ _01149_ _01148_ VGND VGND VPWR VPWR _01187_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18844_ _02128_ _02129_ _02131_ VGND VGND VPWR VPWR _09287_ sky130_fd_sc_hd__o21ai_1
X_11179_ _01115_ _01117_ VGND VGND VPWR VPWR _01118_ sky130_fd_sc_hd__xnor2_1
X_18775_ _09008_ _09022_ _09203_ VGND VGND VPWR VPWR _09211_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15987_ _01350_ _01677_ _06143_ VGND VGND VPWR VPWR _06144_ sky130_fd_sc_hd__a21o_1
XFILLER_0_145_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17726_ net327 _06720_ _08055_ _08056_ VGND VGND VPWR VPWR _08057_ sky130_fd_sc_hd__nand4_1
XFILLER_0_145_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14938_ _04987_ _04954_ _04988_ _04989_ VGND VGND VPWR VPWR _04990_ sky130_fd_sc_hd__nand4_1
X_17657_ net321 _06801_ _07885_ VGND VGND VPWR VPWR _07981_ sky130_fd_sc_hd__and3_1
X_14869_ net440 net168 net163 net445 VGND VGND VPWR VPWR _04914_ sky130_fd_sc_hd__a22oi_1
X_16608_ _06736_ _06737_ VGND VGND VPWR VPWR _06827_ sky130_fd_sc_hd__xnor2_1
X_17588_ _07852_ _07903_ _07904_ VGND VGND VPWR VPWR _07905_ sky130_fd_sc_hd__and3_1
X_19327_ clknet_4_3_0_clock _00019_ VGND VGND VPWR VPWR kd_2\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16539_ _06671_ _06747_ VGND VGND VPWR VPWR _06751_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_128_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19258_ clknet_4_10_0_clock _00140_ VGND VGND VPWR VPWR prev_d_error\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18209_ _07460_ _08501_ _08511_ VGND VGND VPWR VPWR _08588_ sky130_fd_sc_hd__a21boi_2
X_19189_ _09550_ _06130_ _09592_ net492 VGND VGND VPWR VPWR _00149_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_103_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09913_ _06282_ _06381_ VGND VGND VPWR VPWR _06392_ sky130_fd_sc_hd__xor2_1
XFILLER_0_111_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09844_ _05545_ _05622_ VGND VGND VPWR VPWR _05633_ sky130_fd_sc_hd__and2_1
X_09775_ _04863_ VGND VGND VPWR VPWR _04874_ sky130_fd_sc_hd__buf_6
XFILLER_0_96_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10550_ _00486_ _00487_ _00382_ _00488_ VGND VGND VPWR VPWR _00489_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_134_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10481_ _00418_ _00419_ VGND VGND VPWR VPWR _00420_ sky130_fd_sc_hd__nor2_2
X_12220_ _02157_ _02158_ VGND VGND VPWR VPWR _02159_ sky130_fd_sc_hd__nor2_1
X_12151_ _02089_ VGND VGND VPWR VPWR _02090_ sky130_fd_sc_hd__buf_2
XFILLER_0_114_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11102_ _00951_ _01038_ _01017_ _01037_ VGND VGND VPWR VPWR _01041_ sky130_fd_sc_hd__a211o_1
XFILLER_0_102_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12082_ _01987_ _02010_ _02020_ VGND VGND VPWR VPWR _02021_ sky130_fd_sc_hd__or3b_1
X_15910_ _03863_ _06058_ VGND VGND VPWR VPWR _06059_ sky130_fd_sc_hd__and2_1
X_11033_ _00970_ _00971_ VGND VGND VPWR VPWR _00972_ sky130_fd_sc_hd__xnor2_4
X_16890_ _07130_ _07132_ VGND VGND VPWR VPWR _07137_ sky130_fd_sc_hd__nand2_1
X_15841_ _05975_ _05968_ VGND VGND VPWR VPWR _05983_ sky130_fd_sc_hd__and2b_1
XFILLER_0_99_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18560_ _08739_ VGND VGND VPWR VPWR _08974_ sky130_fd_sc_hd__inv_2
X_15772_ _05884_ _05906_ VGND VGND VPWR VPWR _05907_ sky130_fd_sc_hd__nor2_1
X_12984_ _02919_ _02922_ VGND VGND VPWR VPWR _02923_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17511_ _07807_ _07817_ _07819_ VGND VGND VPWR VPWR _07820_ sky130_fd_sc_hd__a21o_1
X_11935_ _01873_ VGND VGND VPWR VPWR _01874_ sky130_fd_sc_hd__clkbuf_4
X_14723_ net426 net174 _04558_ VGND VGND VPWR VPWR _04754_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18491_ _06266_ _08756_ VGND VGND VPWR VPWR _08898_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14654_ _04675_ _04657_ _04661_ VGND VGND VPWR VPWR _04678_ sky130_fd_sc_hd__or3_1
X_17442_ _07677_ _07738_ _07743_ VGND VGND VPWR VPWR _07744_ sky130_fd_sc_hd__a21oi_1
X_11866_ prev_error\[14\] _05402_ VGND VGND VPWR VPWR _01805_ sky130_fd_sc_hd__xnor2_4
X_13605_ _03560_ _03563_ VGND VGND VPWR VPWR _03564_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10817_ _00564_ _00658_ VGND VGND VPWR VPWR _00756_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_151_Left_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14585_ _04597_ _04601_ VGND VGND VPWR VPWR _04602_ sky130_fd_sc_hd__xnor2_1
X_17373_ _07665_ _07666_ _07667_ VGND VGND VPWR VPWR _07669_ sky130_fd_sc_hd__a21o_1
XFILLER_0_156_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11797_ _01704_ _05908_ _05919_ VGND VGND VPWR VPWR _01736_ sky130_fd_sc_hd__nand3_2
XFILLER_0_144_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19112_ net500 prev_error\[17\] VGND VGND VPWR VPWR _09545_ sky130_fd_sc_hd__or2_1
X_13536_ _03461_ _03493_ VGND VGND VPWR VPWR _03495_ sky130_fd_sc_hd__and2b_1
X_16324_ _06419_ _06514_ VGND VGND VPWR VPWR _06515_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10748_ _00685_ _00686_ VGND VGND VPWR VPWR _00687_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19043_ _09448_ _09485_ _09459_ VGND VGND VPWR VPWR _09500_ sky130_fd_sc_hd__a21oi_1
X_16255_ net279 net275 _06410_ _06404_ VGND VGND VPWR VPWR _06439_ sky130_fd_sc_hd__and4_1
XFILLER_0_152_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13467_ _03421_ _03417_ _03419_ VGND VGND VPWR VPWR _03426_ sky130_fd_sc_hd__and3_1
X_10679_ net340 _00409_ _00617_ VGND VGND VPWR VPWR _00618_ sky130_fd_sc_hd__and3_1
XFILLER_0_153_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15206_ _05185_ _05186_ _05187_ _05168_ VGND VGND VPWR VPWR _05285_ sky130_fd_sc_hd__o22a_1
XFILLER_0_112_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12418_ _02350_ _02349_ VGND VGND VPWR VPWR _02357_ sky130_fd_sc_hd__and2b_1
X_16186_ net566 net317 _01755_ _06314_ VGND VGND VPWR VPWR _06363_ sky130_fd_sc_hd__and4_1
X_13398_ net265 _01873_ _03351_ _03352_ VGND VGND VPWR VPWR _03353_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15137_ net471 net153 net149 net477 VGND VGND VPWR VPWR _05209_ sky130_fd_sc_hd__a22oi_1
X_12349_ net221 _01860_ _02287_ VGND VGND VPWR VPWR _02288_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15068_ _05128_ _05132_ VGND VGND VPWR VPWR _05133_ sky130_fd_sc_hd__xnor2_1
X_14019_ _03989_ _03990_ net420 net146 VGND VGND VPWR VPWR _03991_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_156_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18827_ _09266_ _09267_ VGND VGND VPWR VPWR _09268_ sky130_fd_sc_hd__nor2_1
X_18758_ _09136_ _09184_ _09189_ _09190_ _09191_ VGND VGND VPWR VPWR _09192_ sky130_fd_sc_hd__o221ai_4
X_17709_ _08028_ _08037_ _07938_ VGND VGND VPWR VPWR _08038_ sky130_fd_sc_hd__o21ai_2
X_18689_ _09111_ _09114_ _09115_ VGND VGND VPWR VPWR _09116_ sky130_fd_sc_hd__and3_1
XFILLER_0_148_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout400 net403 VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__clkbuf_2
Xfanout411 net412 VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__buf_2
Xfanout422 net424 VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__clkbuf_4
Xfanout433 prev_d_error\[12\] VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__clkbuf_4
Xfanout444 net445 VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout455 prev_d_error\[7\] VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__buf_2
Xfanout466 net468 VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__buf_2
X_09827_ _05391_ _05435_ VGND VGND VPWR VPWR _05446_ sky130_fd_sc_hd__or2_1
Xfanout477 prev_d_error\[2\] VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__buf_2
Xfanout488 net489 VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__clkbuf_4
Xfanout499 net500 VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__buf_2
X_09758_ _04665_ _04610_ _04676_ VGND VGND VPWR VPWR _04687_ sky130_fd_sc_hd__o21ai_4
X_09689_ net51 _03881_ _03914_ net398 VGND VGND VPWR VPWR _00068_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11720_ _01612_ _01648_ _01657_ _01658_ _01578_ VGND VGND VPWR VPWR _01659_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_139_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11651_ net381 _00810_ _01588_ _01589_ VGND VGND VPWR VPWR _01590_ sky130_fd_sc_hd__nand4_1
XFILLER_0_83_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10602_ _00536_ _00540_ VGND VGND VPWR VPWR _00541_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_37_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14370_ _04337_ VGND VGND VPWR VPWR _04365_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11582_ _01516_ _01519_ _01520_ VGND VGND VPWR VPWR _01521_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13321_ _02880_ _03273_ VGND VGND VPWR VPWR _03274_ sky130_fd_sc_hd__xnor2_1
X_10533_ _00371_ _00370_ VGND VGND VPWR VPWR _00472_ sky130_fd_sc_hd__and2b_1
XFILLER_0_51_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16040_ net349 _05600_ VGND VGND VPWR VPWR _06202_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13252_ net225 _02545_ VGND VGND VPWR VPWR _03205_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10464_ net337 _00325_ _00326_ VGND VGND VPWR VPWR _00403_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12203_ _02121_ _02141_ VGND VGND VPWR VPWR _02142_ sky130_fd_sc_hd__xor2_1
X_13183_ _03066_ _03134_ VGND VGND VPWR VPWR _03136_ sky130_fd_sc_hd__nand2_1
X_10395_ net354 _06645_ _00231_ VGND VGND VPWR VPWR _00334_ sky130_fd_sc_hd__and3_1
X_12134_ _02045_ _02071_ _02019_ _02072_ VGND VGND VPWR VPWR _02073_ sky130_fd_sc_hd__o211a_1
X_17991_ _08323_ _08347_ VGND VGND VPWR VPWR _08348_ sky130_fd_sc_hd__xnor2_2
X_16942_ net297 _06620_ _07193_ VGND VGND VPWR VPWR _07194_ sky130_fd_sc_hd__and3_1
X_12065_ _01984_ _02002_ VGND VGND VPWR VPWR _02004_ sky130_fd_sc_hd__and2_1
X_11016_ _00921_ _00953_ _00954_ VGND VGND VPWR VPWR _00955_ sky130_fd_sc_hd__a21oi_1
X_16873_ net324 _06307_ _06308_ VGND VGND VPWR VPWR _07119_ sky130_fd_sc_hd__and3_2
X_18612_ _06116_ _09025_ _09028_ _09030_ _06134_ VGND VGND VPWR VPWR _09031_ sky130_fd_sc_hd__a32oi_4
X_15824_ _04789_ _04893_ VGND VGND VPWR VPWR _05965_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18543_ _08930_ _08796_ _08932_ VGND VGND VPWR VPWR _08956_ sky130_fd_sc_hd__o21ai_1
X_15755_ _05866_ _05888_ VGND VGND VPWR VPWR _05889_ sky130_fd_sc_hd__or2_1
X_12967_ _02884_ _02891_ _02892_ VGND VGND VPWR VPWR _02906_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11918_ net205 _01836_ VGND VGND VPWR VPWR _01857_ sky130_fd_sc_hd__nand2_1
X_14706_ _04532_ _04734_ VGND VGND VPWR VPWR _04735_ sky130_fd_sc_hd__or2_1
X_18474_ _08730_ _08733_ _08876_ _08879_ VGND VGND VPWR VPWR _08880_ sky130_fd_sc_hd__a22o_4
X_15686_ _05796_ _05812_ VGND VGND VPWR VPWR _05813_ sky130_fd_sc_hd__nor2_1
X_12898_ _02814_ _02836_ VGND VGND VPWR VPWR _02837_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17425_ _07257_ _07725_ VGND VGND VPWR VPWR _07726_ sky130_fd_sc_hd__nor2_1
X_11849_ net223 _01787_ VGND VGND VPWR VPWR _01788_ sky130_fd_sc_hd__nand2_1
X_14637_ _04656_ _04634_ _04639_ VGND VGND VPWR VPWR _04659_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14568_ net465 net121 _04482_ VGND VGND VPWR VPWR _04583_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17356_ _07645_ _07649_ VGND VGND VPWR VPWR _07650_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16307_ net288 _06316_ _06318_ _06389_ VGND VGND VPWR VPWR _06496_ sky130_fd_sc_hd__a31o_1
X_13519_ _03362_ _03364_ VGND VGND VPWR VPWR _03478_ sky130_fd_sc_hd__and2_1
X_14499_ _04505_ _04506_ net435 net151 VGND VGND VPWR VPWR _04507_ sky130_fd_sc_hd__and4bb_1
X_17287_ _07572_ _07573_ VGND VGND VPWR VPWR _07574_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19026_ _04148_ _09486_ net492 VGND VGND VPWR VPWR _00076_ sky130_fd_sc_hd__o21a_1
X_16238_ _06419_ _06406_ VGND VGND VPWR VPWR _06420_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16169_ _01805_ _06343_ VGND VGND VPWR VPWR _06344_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_76_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09612_ net50 _03102_ _03135_ net194 VGND VGND VPWR VPWR _00029_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10180_ net360 _05336_ _09318_ _09296_ VGND VGND VPWR VPWR _09329_ sky130_fd_sc_hd__a31o_1
XFILLER_0_100_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout230 net231 VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__buf_2
Xfanout241 kd_1\[7\] VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__buf_2
Xfanout252 net253 VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__buf_2
Xfanout263 net264 VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__buf_2
Xfanout274 net276 VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__buf_2
Xfanout285 ki\[13\] VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__clkbuf_4
Xfanout296 net297 VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__buf_2
X_13870_ _03821_ _03829_ _03831_ VGND VGND VPWR VPWR _03836_ sky130_fd_sc_hd__or3_1
XFILLER_0_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12821_ _02735_ _02759_ VGND VGND VPWR VPWR _02760_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15540_ _05629_ _05627_ VGND VGND VPWR VPWR _05652_ sky130_fd_sc_hd__xnor2_1
X_12752_ net246 _01806_ VGND VGND VPWR VPWR _02691_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11703_ _01640_ _01641_ VGND VGND VPWR VPWR _01642_ sky130_fd_sc_hd__nor2_1
X_15471_ _05573_ _05575_ VGND VGND VPWR VPWR _05576_ sky130_fd_sc_hd__xnor2_1
X_12683_ _02537_ _02621_ VGND VGND VPWR VPWR _02622_ sky130_fd_sc_hd__or2_1
XFILLER_0_139_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14422_ _04327_ _04329_ VGND VGND VPWR VPWR _04422_ sky130_fd_sc_hd__nor2_1
X_17210_ net311 _06620_ VGND VGND VPWR VPWR _07489_ sky130_fd_sc_hd__nand2_1
X_11634_ _01563_ _01571_ _01544_ _01572_ VGND VGND VPWR VPWR _01573_ sky130_fd_sc_hd__o211a_1
X_18190_ i_error\[3\] _08550_ _08551_ VGND VGND VPWR VPWR _08567_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17141_ _07101_ _07103_ VGND VGND VPWR VPWR _07413_ sky130_fd_sc_hd__or2_1
X_14353_ _04344_ _04345_ net420 net155 VGND VGND VPWR VPWR _04347_ sky130_fd_sc_hd__and4bb_1
X_11565_ _01500_ _01503_ VGND VGND VPWR VPWR _01504_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13304_ _03231_ _03256_ VGND VGND VPWR VPWR _03257_ sky130_fd_sc_hd__nor2_1
X_17072_ _07057_ _07212_ _07336_ VGND VGND VPWR VPWR _07337_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10516_ _00431_ _00454_ VGND VGND VPWR VPWR _00455_ sky130_fd_sc_hd__nor2_1
X_14284_ _03998_ _04000_ _04002_ VGND VGND VPWR VPWR _04271_ sky130_fd_sc_hd__or3_1
XFILLER_0_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11496_ net395 _00322_ _01376_ VGND VGND VPWR VPWR _01435_ sky130_fd_sc_hd__and3_1
XFILLER_0_80_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16023_ _08570_ _06181_ _06182_ VGND VGND VPWR VPWR _06184_ sky130_fd_sc_hd__a21o_1
X_13235_ net268 _01806_ VGND VGND VPWR VPWR _03188_ sky130_fd_sc_hd__nand2_1
X_10447_ net361 _06183_ _00385_ _00383_ VGND VGND VPWR VPWR _00386_ sky130_fd_sc_hd__a31o_1
XFILLER_0_123_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13166_ _03061_ _03116_ VGND VGND VPWR VPWR _03117_ sky130_fd_sc_hd__nor2_1
X_10378_ _00227_ _00316_ VGND VGND VPWR VPWR _00317_ sky130_fd_sc_hd__xnor2_1
X_12117_ _02053_ _02055_ VGND VGND VPWR VPWR _02056_ sky130_fd_sc_hd__and2_1
X_13097_ _03037_ _03017_ _03039_ VGND VGND VPWR VPWR _03041_ sky130_fd_sc_hd__and3_1
X_17974_ _08268_ _08329_ VGND VGND VPWR VPWR _08330_ sky130_fd_sc_hd__nor2_1
X_16925_ _07165_ _07174_ _07175_ VGND VGND VPWR VPWR _07176_ sky130_fd_sc_hd__o21a_1
X_12048_ _01984_ _01986_ VGND VGND VPWR VPWR _01987_ sky130_fd_sc_hd__nor2_1
X_16856_ _07098_ _07099_ VGND VGND VPWR VPWR _07100_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15807_ _05673_ _05943_ _05945_ VGND VGND VPWR VPWR _05946_ sky130_fd_sc_hd__o21a_2
X_16787_ _06552_ _06912_ VGND VGND VPWR VPWR _07024_ sky130_fd_sc_hd__xnor2_1
X_13999_ _03969_ _03966_ VGND VGND VPWR VPWR _03971_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18526_ _08799_ _08935_ _08810_ _08936_ VGND VGND VPWR VPWR _08937_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_153_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15738_ _05843_ _05869_ VGND VGND VPWR VPWR _05870_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18457_ _08860_ _08742_ VGND VGND VPWR VPWR _08861_ sky130_fd_sc_hd__nor2_1
X_15669_ net462 net191 _05792_ _05793_ VGND VGND VPWR VPWR _05794_ sky130_fd_sc_hd__and4_1
XFILLER_0_8_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17408_ _07703_ _07706_ VGND VGND VPWR VPWR _07707_ sky130_fd_sc_hd__xor2_2
XFILLER_0_117_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18388_ _08782_ _08784_ VGND VGND VPWR VPWR _08785_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17339_ _07616_ _07617_ _07629_ VGND VGND VPWR VPWR _07631_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19009_ _09135_ _09106_ _09134_ VGND VGND VPWR VPWR _09468_ sky130_fd_sc_hd__and3_1
XFILLER_0_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold38 net85 VGND VGND VPWR VPWR net545 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 i_error\[2\] VGND VGND VPWR VPWR net556 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11350_ _01284_ _01288_ VGND VGND VPWR VPWR _01289_ sky130_fd_sc_hd__and2b_1
XFILLER_0_104_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10301_ _04379_ _04467_ VGND VGND VPWR VPWR _00240_ sky130_fd_sc_hd__nand2_1
X_11281_ _01217_ _01219_ VGND VGND VPWR VPWR _01220_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13020_ _02956_ _02958_ VGND VGND VPWR VPWR _02959_ sky130_fd_sc_hd__nand2_1
X_10232_ _00165_ _00169_ _08053_ _00170_ VGND VGND VPWR VPWR _00171_ sky130_fd_sc_hd__a211oi_1
X_10163_ net371 _05006_ _05578_ VGND VGND VPWR VPWR _09142_ sky130_fd_sc_hd__a21oi_1
X_10094_ _08097_ _06645_ _08372_ VGND VGND VPWR VPWR _08383_ sky130_fd_sc_hd__or3_1
X_14971_ _04965_ _05021_ _05025_ VGND VGND VPWR VPWR _05026_ sky130_fd_sc_hd__or3_1
X_16710_ net566 _01755_ _06316_ VGND VGND VPWR VPWR _06939_ sky130_fd_sc_hd__and3_1
X_13922_ _02173_ _03890_ VGND VGND VPWR VPWR _03891_ sky130_fd_sc_hd__xnor2_1
X_17690_ net298 _07182_ _07568_ net295 VGND VGND VPWR VPWR _08017_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16641_ _06774_ _06861_ VGND VGND VPWR VPWR _06863_ sky130_fd_sc_hd__nand2_1
X_13853_ _03798_ _03804_ VGND VGND VPWR VPWR _03819_ sky130_fd_sc_hd__xnor2_1
X_12804_ _02644_ _02742_ VGND VGND VPWR VPWR _02743_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16572_ _06784_ _06786_ VGND VGND VPWR VPWR _06787_ sky130_fd_sc_hd__xor2_1
X_13784_ _03746_ _03749_ VGND VGND VPWR VPWR _03750_ sky130_fd_sc_hd__nor2_1
X_10996_ _00932_ _00933_ _00934_ VGND VGND VPWR VPWR _00935_ sky130_fd_sc_hd__or3_2
XFILLER_0_85_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18311_ _06514_ _08634_ VGND VGND VPWR VPWR _08700_ sky130_fd_sc_hd__nor2_1
X_15523_ _05623_ _05630_ _05632_ VGND VGND VPWR VPWR _05634_ sky130_fd_sc_hd__a21oi_2
X_12735_ _02571_ _02671_ VGND VGND VPWR VPWR _02674_ sky130_fd_sc_hd__and2_1
X_19291_ clknet_4_8_0_clock _00049_ VGND VGND VPWR VPWR ki\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18242_ _06577_ _06587_ VGND VGND VPWR VPWR _08624_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12666_ _02590_ _02583_ _02589_ VGND VGND VPWR VPWR _02605_ sky130_fd_sc_hd__nand3_1
X_15454_ net467 net484 net171 net153 VGND VGND VPWR VPWR _05558_ sky130_fd_sc_hd__and4_1
XFILLER_0_26_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14405_ _03911_ _04399_ VGND VGND VPWR VPWR _04404_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11617_ _00439_ _00440_ _00600_ _00612_ VGND VGND VPWR VPWR _01556_ sky130_fd_sc_hd__or4b_2
XFILLER_0_115_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18173_ i_error\[4\] _08547_ VGND VGND VPWR VPWR _08549_ sky130_fd_sc_hd__xor2_2
X_12597_ _02534_ _02535_ VGND VGND VPWR VPWR _02536_ sky130_fd_sc_hd__nor2_1
X_15385_ _05480_ _05481_ VGND VGND VPWR VPWR _05482_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17124_ _07358_ _07362_ VGND VGND VPWR VPWR _07395_ sky130_fd_sc_hd__or2b_1
XFILLER_0_25_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14336_ net420 net151 _04257_ _04259_ VGND VGND VPWR VPWR _04328_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_53_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11548_ net390 _00408_ _00323_ net394 VGND VGND VPWR VPWR _01487_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14267_ _04217_ _04229_ VGND VGND VPWR VPWR _04252_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17055_ _07122_ _07317_ _07318_ VGND VGND VPWR VPWR _07319_ sky130_fd_sc_hd__and3_1
X_11479_ _01367_ _01366_ VGND VGND VPWR VPWR _01418_ sky130_fd_sc_hd__and2b_1
XFILLER_0_150_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13218_ _03167_ _03169_ _03170_ VGND VGND VPWR VPWR _03171_ sky130_fd_sc_hd__nand3_1
X_16006_ _00661_ _06164_ VGND VGND VPWR VPWR _06165_ sky130_fd_sc_hd__xnor2_4
X_14198_ _04107_ _04109_ _04174_ VGND VGND VPWR VPWR _04176_ sky130_fd_sc_hd__or3_1
XFILLER_0_57_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13149_ _03012_ _03015_ VGND VGND VPWR VPWR _03098_ sky130_fd_sc_hd__xor2_1
X_17957_ _08219_ _08310_ VGND VGND VPWR VPWR _08311_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_29_Left_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16908_ _07156_ VGND VGND VPWR VPWR _07157_ sky130_fd_sc_hd__clkbuf_4
X_17888_ _08233_ _08234_ _06801_ VGND VGND VPWR VPWR _08235_ sky130_fd_sc_hd__or3b_1
X_16839_ _07078_ _07080_ VGND VGND VPWR VPWR _07081_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18509_ _06266_ _08780_ VGND VGND VPWR VPWR _08918_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_38_Left_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10850_ _00786_ _00788_ _00784_ VGND VGND VPWR VPWR _00789_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10781_ _00699_ _00719_ VGND VGND VPWR VPWR _00720_ sky130_fd_sc_hd__xor2_1
X_12520_ _02422_ _02397_ VGND VGND VPWR VPWR _02459_ sky130_fd_sc_hd__or2b_1
XFILLER_0_109_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_117_Right_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12451_ _02386_ _02388_ _02389_ VGND VGND VPWR VPWR _02390_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11402_ _01337_ _01339_ _01340_ VGND VGND VPWR VPWR _01341_ sky130_fd_sc_hd__nand3_2
X_15170_ _05143_ _05141_ VGND VGND VPWR VPWR _05245_ sky130_fd_sc_hd__nor2_1
X_12382_ _02315_ _02320_ VGND VGND VPWR VPWR _02321_ sky130_fd_sc_hd__and2b_1
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14121_ _04091_ _04090_ VGND VGND VPWR VPWR _04093_ sky130_fd_sc_hd__and2b_1
XFILLER_0_22_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11333_ _01246_ _01271_ VGND VGND VPWR VPWR _01272_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14052_ net412 net418 net144 net138 VGND VGND VPWR VPWR _04024_ sky130_fd_sc_hd__and4_1
X_11264_ net109 _01170_ _01198_ _01202_ VGND VGND VPWR VPWR _01203_ sky130_fd_sc_hd__o211ai_2
X_13003_ _02918_ _02940_ VGND VGND VPWR VPWR _02942_ sky130_fd_sc_hd__nand2_1
X_10215_ _00152_ _00153_ VGND VGND VPWR VPWR _00154_ sky130_fd_sc_hd__and2b_1
X_18860_ _09281_ _09303_ VGND VGND VPWR VPWR _09304_ sky130_fd_sc_hd__and2b_1
X_11195_ _01130_ _01133_ VGND VGND VPWR VPWR _01134_ sky130_fd_sc_hd__xor2_4
XFILLER_0_101_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17811_ _08135_ _08136_ VGND VGND VPWR VPWR _08150_ sky130_fd_sc_hd__nand2_1
X_10146_ _08933_ _08856_ VGND VGND VPWR VPWR _08955_ sky130_fd_sc_hd__and2b_1
X_18791_ _04188_ _04198_ _04196_ VGND VGND VPWR VPWR _09228_ sky130_fd_sc_hd__a21o_1
X_17742_ _08073_ _07980_ VGND VGND VPWR VPWR _08074_ sky130_fd_sc_hd__xnor2_2
X_14954_ net468 net485 net143 net124 VGND VGND VPWR VPWR _05008_ sky130_fd_sc_hd__and4_1
X_10077_ _08185_ VGND VGND VPWR VPWR _08196_ sky130_fd_sc_hd__clkbuf_4
X_13905_ _02983_ _03869_ _03872_ VGND VGND VPWR VPWR _03873_ sky130_fd_sc_hd__a21o_1
X_17673_ net310 _07094_ VGND VGND VPWR VPWR _07999_ sky130_fd_sc_hd__nand2_1
X_14885_ net427 net181 net177 net432 VGND VGND VPWR VPWR _04932_ sky130_fd_sc_hd__a22o_1
X_16624_ net303 _06353_ VGND VGND VPWR VPWR _06845_ sky130_fd_sc_hd__nand2_1
X_13836_ _03791_ _03796_ _03801_ VGND VGND VPWR VPWR _03802_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_58_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19343_ clknet_4_0_0_clock _00026_ VGND VGND VPWR VPWR kd_2\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16555_ _06694_ _06768_ VGND VGND VPWR VPWR _06769_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13767_ _01763_ _03731_ _03732_ VGND VGND VPWR VPWR _03733_ sky130_fd_sc_hd__o21a_1
X_10979_ _00826_ _00898_ VGND VGND VPWR VPWR _00918_ sky130_fd_sc_hd__nor2_1
X_15506_ _05591_ _05598_ _05607_ VGND VGND VPWR VPWR _05615_ sky130_fd_sc_hd__nor3_1
XFILLER_0_17_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12718_ _02645_ _02656_ _02654_ VGND VGND VPWR VPWR _02657_ sky130_fd_sc_hd__a21oi_2
X_19274_ clknet_4_6_0_clock _00070_ VGND VGND VPWR VPWR kp\[4\] sky130_fd_sc_hd__dfxtp_1
X_16486_ _06629_ _06631_ VGND VGND VPWR VPWR _06693_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13698_ _03662_ _03663_ VGND VGND VPWR VPWR _03664_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18225_ _08604_ _08605_ VGND VGND VPWR VPWR _08606_ sky130_fd_sc_hd__xnor2_4
X_15437_ _05529_ _05537_ _05538_ VGND VGND VPWR VPWR _05539_ sky130_fd_sc_hd__o21ai_2
X_12649_ _02582_ _02580_ VGND VGND VPWR VPWR _02588_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18156_ _06837_ _06933_ VGND VGND VPWR VPWR _08530_ sky130_fd_sc_hd__or2_1
X_15368_ _05376_ _05462_ VGND VGND VPWR VPWR _05463_ sky130_fd_sc_hd__nor2_1
X_17107_ net282 _06803_ _07088_ VGND VGND VPWR VPWR _07376_ sky130_fd_sc_hd__a21oi_1
X_14319_ _04307_ _04308_ net448 net128 VGND VGND VPWR VPWR _04309_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_41_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18087_ _08451_ _08452_ _08453_ _07351_ VGND VGND VPWR VPWR _08454_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_7_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15299_ _05360_ _05386_ VGND VGND VPWR VPWR _05387_ sky130_fd_sc_hd__or2b_1
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17038_ net324 net320 _06351_ _06344_ VGND VGND VPWR VPWR _07300_ sky130_fd_sc_hd__nand4_1
XFILLER_0_1_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09860_ _05765_ _05798_ VGND VGND VPWR VPWR _05809_ sky130_fd_sc_hd__xor2_1
XFILLER_0_21_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09791_ _04929_ _05017_ _05028_ VGND VGND VPWR VPWR _05050_ sky130_fd_sc_hd__nand3_2
X_18989_ _09357_ _09445_ VGND VGND VPWR VPWR _09446_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_84_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_46_Left_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_55_Left_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10000_ _07316_ _07338_ VGND VGND VPWR VPWR _07349_ sky130_fd_sc_hd__nand2_2
X_09989_ _07206_ _07217_ VGND VGND VPWR VPWR _07228_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11951_ _01867_ _01879_ _01889_ VGND VGND VPWR VPWR _01890_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10902_ _00764_ _00766_ _00676_ VGND VGND VPWR VPWR _00841_ sky130_fd_sc_hd__a21o_1
X_14670_ _04688_ _04694_ VGND VGND VPWR VPWR _04695_ sky130_fd_sc_hd__and2_1
X_11882_ _01804_ _01820_ VGND VGND VPWR VPWR _01821_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_64_Left_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13621_ _03574_ _03577_ _03579_ VGND VGND VPWR VPWR _03580_ sky130_fd_sc_hd__o21a_1
X_10833_ _00769_ _00770_ _00771_ VGND VGND VPWR VPWR _00772_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_39_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16340_ _06530_ _06531_ VGND VGND VPWR VPWR _06532_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13552_ _03509_ _03510_ VGND VGND VPWR VPWR _03511_ sky130_fd_sc_hd__and2_1
X_10764_ net565 _00243_ _00226_ _06931_ VGND VGND VPWR VPWR _00703_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_94_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12503_ _02375_ _02441_ VGND VGND VPWR VPWR _02442_ sky130_fd_sc_hd__or2_1
X_13483_ _03435_ _03441_ VGND VGND VPWR VPWR _03442_ sky130_fd_sc_hd__nor2_1
X_16271_ net289 _06353_ _06346_ net286 VGND VGND VPWR VPWR _06456_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10695_ _00568_ _00566_ VGND VGND VPWR VPWR _00634_ sky130_fd_sc_hd__and2b_1
XFILLER_0_152_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18010_ _08367_ _08365_ VGND VGND VPWR VPWR _08369_ sky130_fd_sc_hd__xnor2_1
X_12434_ _02265_ _02372_ VGND VGND VPWR VPWR _02373_ sky130_fd_sc_hd__nor2_1
X_15222_ _05225_ _05227_ _05238_ VGND VGND VPWR VPWR _05302_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12365_ _02301_ _02303_ VGND VGND VPWR VPWR _02304_ sky130_fd_sc_hd__or2_2
X_15153_ _05224_ _05213_ _05222_ VGND VGND VPWR VPWR _05227_ sky130_fd_sc_hd__nand3_1
XFILLER_0_121_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_73_Left_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14104_ net434 net117 VGND VGND VPWR VPWR _04076_ sky130_fd_sc_hd__nand2_1
X_11316_ _01049_ _01180_ VGND VGND VPWR VPWR _01255_ sky130_fd_sc_hd__xnor2_1
X_15084_ _05068_ _05067_ VGND VGND VPWR VPWR _05151_ sky130_fd_sc_hd__and2b_1
X_12296_ _02099_ _02100_ VGND VGND VPWR VPWR _02235_ sky130_fd_sc_hd__nand2_1
X_14035_ net407 net151 _04004_ _04005_ VGND VGND VPWR VPWR _04007_ sky130_fd_sc_hd__o2bb2a_1
X_18912_ _09280_ _09328_ _09326_ VGND VGND VPWR VPWR _09361_ sky130_fd_sc_hd__a21oi_1
X_11247_ _01174_ _01184_ _01185_ VGND VGND VPWR VPWR _01186_ sky130_fd_sc_hd__a21bo_1
X_18843_ _02126_ _02136_ VGND VGND VPWR VPWR _09286_ sky130_fd_sc_hd__nand2_1
X_11178_ _01033_ _01116_ VGND VGND VPWR VPWR _01117_ sky130_fd_sc_hd__xor2_1
X_10129_ _08537_ _08757_ VGND VGND VPWR VPWR _08768_ sky130_fd_sc_hd__xnor2_1
X_18774_ _08996_ _09204_ VGND VGND VPWR VPWR _09210_ sky130_fd_sc_hd__and2_1
X_15986_ _01212_ _01278_ VGND VGND VPWR VPWR _06143_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_145_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17725_ net325 _06800_ _06889_ net318 VGND VGND VPWR VPWR _08056_ sky130_fd_sc_hd__a22o_1
X_14937_ _04851_ _04956_ _04986_ VGND VGND VPWR VPWR _04989_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_82_Left_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17656_ _07885_ _07979_ VGND VGND VPWR VPWR _07980_ sky130_fd_sc_hd__xnor2_2
X_14868_ net439 net445 net168 net163 VGND VGND VPWR VPWR _04913_ sky130_fd_sc_hd__and4_1
XFILLER_0_89_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16607_ _06753_ _06790_ _06825_ VGND VGND VPWR VPWR _06826_ sky130_fd_sc_hd__o21a_1
X_13819_ _03752_ _03784_ VGND VGND VPWR VPWR _03785_ sky130_fd_sc_hd__or2_1
X_17587_ _07849_ _07851_ _07848_ VGND VGND VPWR VPWR _07904_ sky130_fd_sc_hd__o21ai_1
X_14799_ _04835_ _04833_ VGND VGND VPWR VPWR _04837_ sky130_fd_sc_hd__xnor2_1
X_19326_ clknet_4_0_0_clock _00009_ VGND VGND VPWR VPWR kd_1\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16538_ _06748_ _06749_ VGND VGND VPWR VPWR _06750_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19257_ clknet_4_10_0_clock _00139_ VGND VGND VPWR VPWR prev_d_error\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16469_ _06368_ _06379_ _06673_ VGND VGND VPWR VPWR _06674_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18208_ i_error\[11\] _08586_ VGND VGND VPWR VPWR _08587_ sky130_fd_sc_hd__xnor2_2
X_19188_ net507 net414 VGND VGND VPWR VPWR _09592_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18139_ _07444_ _07458_ VGND VGND VPWR VPWR _08511_ sky130_fd_sc_hd__or2b_1
XFILLER_0_14_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09912_ _06359_ _06370_ VGND VGND VPWR VPWR _06381_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09843_ _05589_ _05611_ VGND VGND VPWR VPWR _05622_ sky130_fd_sc_hd__nor2_1
X_09774_ _04841_ _04852_ VGND VGND VPWR VPWR _04863_ sky130_fd_sc_hd__and2_1
XFILLER_0_139_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10480_ _00417_ _00405_ _00416_ VGND VGND VPWR VPWR _00419_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12150_ _02088_ VGND VGND VPWR VPWR _02089_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11101_ _01023_ _01034_ _01021_ VGND VGND VPWR VPWR _01040_ sky130_fd_sc_hd__a21o_1
X_12081_ _02015_ _02019_ VGND VGND VPWR VPWR _02020_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11032_ net383 _06183_ VGND VGND VPWR VPWR _00971_ sky130_fd_sc_hd__nand2_2
X_15840_ _05980_ _05967_ _04787_ VGND VGND VPWR VPWR _05982_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15771_ _05876_ _05883_ VGND VGND VPWR VPWR _05906_ sky130_fd_sc_hd__nor2_1
X_12983_ net211 _02641_ _02921_ VGND VGND VPWR VPWR _02922_ sky130_fd_sc_hd__and3_1
X_17510_ _07576_ _07818_ VGND VGND VPWR VPWR _07819_ sky130_fd_sc_hd__or2_1
X_14722_ _04016_ net186 VGND VGND VPWR VPWR _04752_ sky130_fd_sc_hd__nor2_1
X_11934_ _01872_ VGND VGND VPWR VPWR _01873_ sky130_fd_sc_hd__clkbuf_4
X_18490_ _08894_ _08737_ _08738_ net100 _08750_ VGND VGND VPWR VPWR _08897_ sky130_fd_sc_hd__o32a_1
XFILLER_0_24_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17441_ _07740_ _07742_ VGND VGND VPWR VPWR _07743_ sky130_fd_sc_hd__xnor2_1
X_14653_ _04657_ _04661_ _04675_ VGND VGND VPWR VPWR _04677_ sky130_fd_sc_hd__o21a_1
X_11865_ _01802_ _01803_ VGND VGND VPWR VPWR _01804_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13604_ _03561_ _03562_ VGND VGND VPWR VPWR _03563_ sky130_fd_sc_hd__xnor2_1
X_17372_ net280 net277 _02932_ net540 VGND VGND VPWR VPWR _07667_ sky130_fd_sc_hd__and4_1
X_10816_ _00662_ _00754_ VGND VGND VPWR VPWR _00755_ sky130_fd_sc_hd__nor2_1
X_14584_ _04598_ _04600_ _03917_ VGND VGND VPWR VPWR _04601_ sky130_fd_sc_hd__mux2_1
X_11796_ prev_error\[10\] _06194_ VGND VGND VPWR VPWR _01735_ sky130_fd_sc_hd__or2b_1
XFILLER_0_95_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19111_ _09536_ _04896_ _09544_ net488 VGND VGND VPWR VPWR _00111_ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16323_ net280 _06336_ VGND VGND VPWR VPWR _06514_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13535_ _03461_ _03493_ VGND VGND VPWR VPWR _03494_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_131_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10747_ net368 _06634_ _06183_ net371 VGND VGND VPWR VPWR _00686_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_54_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19042_ _04126_ net95 VGND VGND VPWR VPWR _09498_ sky130_fd_sc_hd__and2_1
X_16254_ _06437_ VGND VGND VPWR VPWR _06438_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13466_ _03423_ _03424_ VGND VGND VPWR VPWR _03425_ sky130_fd_sc_hd__nand2_1
X_10678_ net343 _00515_ VGND VGND VPWR VPWR _00617_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15205_ _05265_ _05282_ _05283_ VGND VGND VPWR VPWR _05284_ sky130_fd_sc_hd__nand3_1
XFILLER_0_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12417_ _02353_ _02355_ VGND VGND VPWR VPWR _02356_ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16185_ net566 net317 VGND VGND VPWR VPWR _06362_ sky130_fd_sc_hd__or2_1
X_13397_ _03349_ _03350_ VGND VGND VPWR VPWR _03352_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15136_ net471 net476 net153 net148 VGND VGND VPWR VPWR _05208_ sky130_fd_sc_hd__and4_1
X_12348_ _02284_ _02286_ VGND VGND VPWR VPWR _02287_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15067_ _05129_ _05130_ _05131_ VGND VGND VPWR VPWR _05132_ sky130_fd_sc_hd__o21ba_1
X_12279_ _01710_ _01728_ VGND VGND VPWR VPWR _02218_ sky130_fd_sc_hd__nand2_2
XFILLER_0_120_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14018_ net425 net141 net137 net430 VGND VGND VPWR VPWR _03990_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_65_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18826_ _09264_ _09265_ VGND VGND VPWR VPWR _09267_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18757_ _09149_ _09162_ _09148_ VGND VGND VPWR VPWR _09191_ sky130_fd_sc_hd__a21oi_1
X_15969_ _06019_ _06122_ _06123_ VGND VGND VPWR VPWR _06124_ sky130_fd_sc_hd__o21bai_4
X_17708_ _08025_ _08030_ VGND VGND VPWR VPWR _08037_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18688_ _08929_ _09075_ _09077_ VGND VGND VPWR VPWR _09115_ sky130_fd_sc_hd__nand3_1
XFILLER_0_78_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17639_ _07952_ _07959_ _07960_ _07872_ VGND VGND VPWR VPWR _07961_ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19309_ clknet_4_1_0_clock _00010_ VGND VGND VPWR VPWR kd_1\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout401 net402 VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__clkbuf_4
Xfanout412 net415 VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__clkbuf_4
Xfanout423 net424 VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__clkbuf_2
Xfanout434 net435 VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__buf_2
Xfanout445 prev_d_error\[9\] VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__clkbuf_4
Xfanout456 net458 VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__buf_2
X_09826_ net353 _05424_ _05182_ net356 VGND VGND VPWR VPWR _05435_ sky130_fd_sc_hd__a22oi_1
Xfanout467 net468 VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__buf_2
Xfanout478 net480 VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__clkbuf_2
Xfanout489 net497 VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__buf_2
X_09757_ _04555_ _04577_ _04544_ VGND VGND VPWR VPWR _04676_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_96_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09688_ net50 _03881_ _03914_ net403 VGND VGND VPWR VPWR _00067_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11650_ net385 _00814_ _01001_ net564 VGND VGND VPWR VPWR _01589_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10601_ _00537_ _00539_ VGND VGND VPWR VPWR _00540_ sky130_fd_sc_hd__and2_2
X_11581_ net366 _00812_ VGND VGND VPWR VPWR _01520_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10532_ net372 _05325_ VGND VGND VPWR VPWR _00471_ sky130_fd_sc_hd__nand2_2
X_13320_ net253 _01907_ VGND VGND VPWR VPWR _03273_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13251_ _03112_ _03111_ VGND VGND VPWR VPWR _03204_ sky130_fd_sc_hd__or2b_1
X_10463_ net350 _09583_ _00401_ VGND VGND VPWR VPWR _00402_ sky130_fd_sc_hd__and3_1
X_12202_ _02122_ _02140_ VGND VGND VPWR VPWR _02141_ sky130_fd_sc_hd__xor2_2
XFILLER_0_20_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13182_ _02225_ _03065_ _02926_ VGND VGND VPWR VPWR _03134_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10394_ net354 _06645_ _00231_ VGND VGND VPWR VPWR _00333_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12133_ _01846_ _02016_ _02018_ VGND VGND VPWR VPWR _02072_ sky130_fd_sc_hd__o21ai_1
X_17990_ _08345_ _08346_ VGND VGND VPWR VPWR _08347_ sky130_fd_sc_hd__nor2_1
X_12064_ _01984_ _02002_ VGND VGND VPWR VPWR _02003_ sky130_fd_sc_hd__nor2_1
X_16941_ net299 _06463_ _06465_ VGND VGND VPWR VPWR _07193_ sky130_fd_sc_hd__and3_2
X_11015_ _00922_ _00952_ VGND VGND VPWR VPWR _00954_ sky130_fd_sc_hd__nor2_1
X_16872_ _07081_ _07116_ VGND VGND VPWR VPWR _07117_ sky130_fd_sc_hd__nor2_1
X_18611_ _09029_ _09028_ VGND VGND VPWR VPWR _09030_ sky130_fd_sc_hd__xnor2_2
X_15823_ _04998_ _05962_ VGND VGND VPWR VPWR _05964_ sky130_fd_sc_hd__or2_1
X_18542_ net524 _08947_ _08949_ _08950_ _08953_ VGND VGND VPWR VPWR _08954_ sky130_fd_sc_hd__a221o_1
X_15754_ _05868_ _05885_ _05887_ VGND VGND VPWR VPWR _05888_ sky130_fd_sc_hd__or3b_1
X_12966_ _02895_ _02900_ _02904_ VGND VGND VPWR VPWR _02905_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14705_ _04526_ _04531_ VGND VGND VPWR VPWR _04734_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11917_ _01837_ _01840_ VGND VGND VPWR VPWR _01856_ sky130_fd_sc_hd__nor2_1
X_18473_ _08728_ _08729_ _08733_ _08877_ _08874_ VGND VGND VPWR VPWR _08879_ sky130_fd_sc_hd__o32a_1
X_15685_ _05795_ _05790_ VGND VGND VPWR VPWR _05812_ sky130_fd_sc_hd__and2b_1
X_12897_ _02830_ _02816_ VGND VGND VPWR VPWR _02836_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17424_ _07254_ _07256_ VGND VGND VPWR VPWR _07725_ sky130_fd_sc_hd__and2_1
XFILLER_0_157_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14636_ _04556_ _04580_ VGND VGND VPWR VPWR _04658_ sky130_fd_sc_hd__xnor2_1
X_11848_ _01786_ VGND VGND VPWR VPWR _01787_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17355_ _07262_ _07648_ VGND VGND VPWR VPWR _07649_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_144_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14567_ net465 net121 _04482_ VGND VGND VPWR VPWR _04582_ sky130_fd_sc_hd__and3_1
X_11779_ prev_error\[1\] _00814_ VGND VGND VPWR VPWR _01718_ sky130_fd_sc_hd__and2b_1
X_16306_ net283 _06336_ VGND VGND VPWR VPWR _06495_ sky130_fd_sc_hd__nand2_1
X_13518_ _03476_ VGND VGND VPWR VPWR _03477_ sky130_fd_sc_hd__inv_2
X_17286_ _07565_ _07566_ _07570_ net281 VGND VGND VPWR VPWR _07573_ sky130_fd_sc_hd__a22o_1
X_14498_ net439 net147 net142 net443 VGND VGND VPWR VPWR _04506_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_24_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19025_ net522 _09485_ _09466_ VGND VGND VPWR VPWR _09486_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16237_ net275 _06386_ VGND VGND VPWR VPWR _06419_ sky130_fd_sc_hd__nand2_1
X_13449_ _03323_ _03385_ _03368_ _03384_ VGND VGND VPWR VPWR _03408_ sky130_fd_sc_hd__a211o_1
XFILLER_0_3_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16168_ _06298_ _01742_ _06297_ _06302_ VGND VGND VPWR VPWR _06343_ sky130_fd_sc_hd__a31o_2
XFILLER_0_23_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15119_ _05087_ _05088_ _05089_ _05064_ VGND VGND VPWR VPWR _05189_ sky130_fd_sc_hd__a22o_1
X_16099_ _06174_ _01698_ VGND VGND VPWR VPWR _06267_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_10_Left_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09611_ net40 _03102_ _03135_ kd_2\[0\] VGND VGND VPWR VPWR _00019_ sky130_fd_sc_hd__a22o_1
X_18809_ _04178_ _04182_ _09246_ VGND VGND VPWR VPWR _09248_ sky130_fd_sc_hd__nand3_1
XFILLER_0_78_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout220 kd_1\[12\] VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__buf_2
Xfanout231 net233 VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__clkbuf_4
Xfanout242 net245 VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__clkbuf_4
Xfanout253 kd_1\[4\] VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__clkbuf_2
Xfanout264 net266 VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__clkbuf_4
Xfanout275 net276 VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__clkbuf_4
Xfanout286 net287 VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__clkbuf_4
X_09809_ _05116_ _05237_ VGND VGND VPWR VPWR _05248_ sky130_fd_sc_hd__or2b_1
Xfanout297 ki\[10\] VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__clkbuf_4
X_12820_ _02756_ _02758_ VGND VGND VPWR VPWR _02759_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12751_ _01813_ _02364_ _02689_ VGND VGND VPWR VPWR _02690_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_38_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11702_ _01636_ _01639_ VGND VGND VPWR VPWR _01641_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15470_ _05495_ _05574_ VGND VGND VPWR VPWR _05575_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12682_ net209 _02224_ _02536_ VGND VGND VPWR VPWR _02621_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14421_ _04418_ _04420_ VGND VGND VPWR VPWR _04421_ sky130_fd_sc_hd__and2_1
X_11633_ _01540_ _01543_ _01542_ VGND VGND VPWR VPWR _01572_ sky130_fd_sc_hd__a21o_1
XFILLER_0_108_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17140_ _07164_ _07171_ VGND VGND VPWR VPWR _07412_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14352_ net425 net152 net147 net430 VGND VGND VPWR VPWR _04345_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_25_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11564_ _01501_ _01502_ VGND VGND VPWR VPWR _01503_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13303_ _03251_ _03255_ VGND VGND VPWR VPWR _03256_ sky130_fd_sc_hd__and2_1
X_17071_ net305 _06409_ _06345_ net308 VGND VGND VPWR VPWR _07336_ sky130_fd_sc_hd__a22o_1
X_10515_ _00432_ _00452_ _00453_ VGND VGND VPWR VPWR _00454_ sky130_fd_sc_hd__a21oi_1
X_14283_ _04264_ _04266_ _04268_ VGND VGND VPWR VPWR _04270_ sky130_fd_sc_hd__o21ai_2
X_11495_ net395 _00243_ _00323_ net390 VGND VGND VPWR VPWR _01434_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16022_ net342 _04896_ _05677_ net344 VGND VGND VPWR VPWR _06182_ sky130_fd_sc_hd__a22oi_1
X_13234_ net252 _01873_ VGND VGND VPWR VPWR _03187_ sky130_fd_sc_hd__nand2_1
X_10446_ _00383_ _00384_ VGND VGND VPWR VPWR _00385_ sky130_fd_sc_hd__nor2_1
X_13165_ net211 _02746_ _03060_ VGND VGND VPWR VPWR _03116_ sky130_fd_sc_hd__a21oi_1
X_10377_ _00253_ _00252_ VGND VGND VPWR VPWR _00316_ sky130_fd_sc_hd__nor2_1
X_12116_ net226 _01814_ _01799_ net230 VGND VGND VPWR VPWR _02055_ sky130_fd_sc_hd__a22o_1
X_13096_ _03037_ _03017_ _03039_ VGND VGND VPWR VPWR _03040_ sky130_fd_sc_hd__a21oi_2
X_17973_ net326 _07094_ _08267_ VGND VGND VPWR VPWR _08329_ sky130_fd_sc_hd__a21oi_1
X_16924_ net288 _06803_ _06891_ net285 VGND VGND VPWR VPWR _07175_ sky130_fd_sc_hd__a22o_1
X_12047_ _01951_ _01985_ VGND VGND VPWR VPWR _01986_ sky130_fd_sc_hd__or2_1
X_16855_ _06989_ _07097_ VGND VGND VPWR VPWR _07099_ sky130_fd_sc_hd__and2_1
X_15806_ _05613_ _05944_ VGND VGND VPWR VPWR _05945_ sky130_fd_sc_hd__xnor2_1
X_16786_ _07016_ _07021_ _07022_ _06542_ VGND VGND VPWR VPWR _07023_ sky130_fd_sc_hd__a211o_1
X_13998_ _03966_ _03969_ VGND VGND VPWR VPWR _03970_ sky130_fd_sc_hd__and2b_1
X_18525_ _06261_ _06264_ _08808_ VGND VGND VPWR VPWR _08936_ sky130_fd_sc_hd__a21oi_1
X_15737_ _05839_ _05841_ VGND VGND VPWR VPWR _05869_ sky130_fd_sc_hd__and2_1
X_12949_ net245 _01852_ _02887_ VGND VGND VPWR VPWR _02888_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_88_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18456_ _06166_ _08859_ VGND VGND VPWR VPWR _08860_ sky130_fd_sc_hd__nand2_1
X_15668_ net466 net187 net171 net483 VGND VGND VPWR VPWR _05793_ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17407_ _07704_ _07705_ VGND VGND VPWR VPWR _07706_ sky130_fd_sc_hd__xnor2_2
X_14619_ _04636_ _04638_ VGND VGND VPWR VPWR _04639_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18387_ _08783_ _08544_ VGND VGND VPWR VPWR _08784_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15599_ _05713_ _05714_ _05716_ VGND VGND VPWR VPWR _05717_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17338_ _07616_ _07617_ _07629_ VGND VGND VPWR VPWR _07630_ sky130_fd_sc_hd__or3_4
XFILLER_0_43_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17269_ net292 _07094_ _07552_ VGND VGND VPWR VPWR _07554_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_153_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19008_ _09135_ _09106_ _09134_ VGND VGND VPWR VPWR _09467_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold39 net88 VGND VGND VPWR VPWR net546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_127_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10300_ _04346_ VGND VGND VPWR VPWR _00239_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11280_ _01147_ _01218_ VGND VGND VPWR VPWR _01219_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10231_ _08020_ _08031_ _08042_ VGND VGND VPWR VPWR _00170_ sky130_fd_sc_hd__o21a_1
XFILLER_0_131_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10162_ _08504_ _09120_ VGND VGND VPWR VPWR _09131_ sky130_fd_sc_hd__xnor2_4
X_10093_ _08152_ _08361_ VGND VGND VPWR VPWR _08372_ sky130_fd_sc_hd__xnor2_1
X_14970_ _05022_ _05023_ _05024_ VGND VGND VPWR VPWR _05025_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_100_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13921_ _02252_ _02254_ _03889_ VGND VGND VPWR VPWR _03890_ sky130_fd_sc_hd__a21boi_2
X_16640_ _06774_ _06861_ VGND VGND VPWR VPWR _06862_ sky130_fd_sc_hd__nor2_1
X_13852_ _03813_ _03815_ _03817_ VGND VGND VPWR VPWR _03818_ sky130_fd_sc_hd__o21a_1
X_12803_ net202 _02641_ _02643_ VGND VGND VPWR VPWR _02742_ sky130_fd_sc_hd__a21oi_1
X_16571_ _06649_ _06785_ _06548_ VGND VGND VPWR VPWR _06786_ sky130_fd_sc_hd__a21bo_1
X_13783_ _03747_ _03746_ _03748_ VGND VGND VPWR VPWR _03749_ sky130_fd_sc_hd__nor3_1
XFILLER_0_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10995_ _00926_ _00930_ VGND VGND VPWR VPWR _00934_ sky130_fd_sc_hd__xor2_1
X_18310_ _08631_ _08641_ _08639_ VGND VGND VPWR VPWR _08699_ sky130_fd_sc_hd__a21oi_1
X_15522_ _05597_ _05631_ VGND VGND VPWR VPWR _05632_ sky130_fd_sc_hd__or2_1
X_12734_ _02570_ _02672_ VGND VGND VPWR VPWR _02673_ sky130_fd_sc_hd__nand2_1
X_19290_ clknet_4_8_0_clock _00048_ VGND VGND VPWR VPWR ki\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18241_ _08622_ VGND VGND VPWR VPWR _08623_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15453_ net467 net171 VGND VGND VPWR VPWR _05557_ sky130_fd_sc_hd__nand2_1
X_12665_ _02597_ _02603_ VGND VGND VPWR VPWR _02604_ sky130_fd_sc_hd__xor2_1
XFILLER_0_26_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14404_ _04399_ _04402_ VGND VGND VPWR VPWR _04403_ sky130_fd_sc_hd__nor2_1
X_11616_ _01554_ _01532_ VGND VGND VPWR VPWR _01555_ sky130_fd_sc_hd__xnor2_1
X_18172_ _08546_ _08439_ VGND VGND VPWR VPWR _08547_ sky130_fd_sc_hd__xnor2_2
X_15384_ net463 net172 _05477_ _05478_ VGND VGND VPWR VPWR _05481_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_154_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12596_ net214 _02091_ _01909_ net217 VGND VGND VPWR VPWR _02535_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_52_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17123_ _07375_ _07377_ VGND VGND VPWR VPWR _07394_ sky130_fd_sc_hd__and2b_1
X_14335_ _04325_ _04322_ VGND VGND VPWR VPWR _04327_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11547_ net400 _09577_ _01485_ _01434_ VGND VGND VPWR VPWR _01486_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17054_ net329 _06324_ _07120_ _07121_ VGND VGND VPWR VPWR _07318_ sky130_fd_sc_hd__a22o_1
X_14266_ _04248_ _04250_ VGND VGND VPWR VPWR _04251_ sky130_fd_sc_hd__nand2_1
X_11478_ net370 _00614_ VGND VGND VPWR VPWR _01417_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16005_ _00759_ _01690_ _00757_ VGND VGND VPWR VPWR _06164_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_0_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13217_ _03048_ _03166_ _03161_ _03165_ VGND VGND VPWR VPWR _03170_ sky130_fd_sc_hd__a211o_1
XFILLER_0_111_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10429_ _00365_ _00366_ _00367_ VGND VGND VPWR VPWR _00368_ sky130_fd_sc_hd__a21o_1
X_14197_ _04107_ _04109_ _04174_ VGND VGND VPWR VPWR _04175_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13148_ net248 _01874_ _03096_ _03095_ VGND VGND VPWR VPWR _03097_ sky130_fd_sc_hd__a31o_1
XFILLER_0_148_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13079_ _03019_ _03020_ VGND VGND VPWR VPWR _03021_ sky130_fd_sc_hd__nor2_1
X_17956_ _08216_ _08217_ _08210_ VGND VGND VPWR VPWR _08310_ sky130_fd_sc_hd__o21ai_1
X_16907_ _07155_ VGND VGND VPWR VPWR _07156_ sky130_fd_sc_hd__clkbuf_4
X_17887_ net331 _07155_ VGND VGND VPWR VPWR _08234_ sky130_fd_sc_hd__nand2_1
X_16838_ _07066_ _07079_ VGND VGND VPWR VPWR _07080_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16769_ _06891_ _07003_ net270 VGND VGND VPWR VPWR _07004_ sky130_fd_sc_hd__and3b_1
X_18508_ _08893_ _08739_ _08897_ net99 _08916_ VGND VGND VPWR VPWR _08917_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_119_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18439_ _08840_ _08743_ VGND VGND VPWR VPWR _08841_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_102_Left_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10780_ _00700_ _00717_ _00718_ VGND VGND VPWR VPWR _00719_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12450_ _02381_ _02384_ _02379_ VGND VGND VPWR VPWR _02389_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11401_ _01268_ _01336_ _01331_ _01335_ VGND VGND VPWR VPWR _01340_ sky130_fd_sc_hd__a211o_1
XFILLER_0_124_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12381_ _02316_ _02319_ VGND VGND VPWR VPWR _02320_ sky130_fd_sc_hd__or2_1
X_14120_ _04090_ _04091_ VGND VGND VPWR VPWR _04092_ sky130_fd_sc_hd__and2b_1
XFILLER_0_105_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11332_ _01248_ _01269_ _01270_ VGND VGND VPWR VPWR _01271_ sky130_fd_sc_hd__a21bo_2
X_14051_ _04017_ net151 VGND VGND VPWR VPWR _04023_ sky130_fd_sc_hd__nor2_1
X_11263_ _01198_ _01200_ _01201_ VGND VGND VPWR VPWR _01202_ sky130_fd_sc_hd__nand3_2
X_13002_ _02918_ _02940_ VGND VGND VPWR VPWR _02941_ sky130_fd_sc_hd__or2_1
X_10214_ _09527_ _09491_ VGND VGND VPWR VPWR _00153_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11194_ _01131_ _01132_ VGND VGND VPWR VPWR _01133_ sky130_fd_sc_hd__xor2_4
X_10145_ _08856_ _08933_ VGND VGND VPWR VPWR _08944_ sky130_fd_sc_hd__and2b_1
X_17810_ _08126_ _08142_ VGND VGND VPWR VPWR _08149_ sky130_fd_sc_hd__nand2_1
X_18790_ _04163_ _04184_ _04186_ VGND VGND VPWR VPWR _09227_ sky130_fd_sc_hd__a21oi_2
X_17741_ net327 _06619_ VGND VGND VPWR VPWR _08073_ sky130_fd_sc_hd__nand2_1
X_14953_ net462 net148 VGND VGND VPWR VPWR _05007_ sky130_fd_sc_hd__nand2_1
X_10076_ _08174_ VGND VGND VPWR VPWR _08185_ sky130_fd_sc_hd__buf_2
X_13904_ _02873_ _03871_ VGND VGND VPWR VPWR _03872_ sky130_fd_sc_hd__nand2_1
X_17672_ net310 _06992_ _07094_ net307 VGND VGND VPWR VPWR _07997_ sky130_fd_sc_hd__a22o_1
X_14884_ net427 net432 net181 net177 VGND VGND VPWR VPWR _04931_ sky130_fd_sc_hd__and4_1
X_16623_ _06841_ _06842_ VGND VGND VPWR VPWR _06844_ sky130_fd_sc_hd__or2b_1
X_13835_ _03799_ _03800_ VGND VGND VPWR VPWR _03801_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16554_ _06692_ _06693_ VGND VGND VPWR VPWR _06768_ sky130_fd_sc_hd__nor2_1
X_19342_ clknet_4_0_0_clock _00025_ VGND VGND VPWR VPWR kd_2\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13766_ net247 _02913_ _03730_ VGND VGND VPWR VPWR _03732_ sky130_fd_sc_hd__a21o_1
X_10978_ _00899_ _00915_ _00916_ VGND VGND VPWR VPWR _00917_ sky130_fd_sc_hd__o21ba_1
X_15505_ _05461_ _05543_ _05539_ _05542_ VGND VGND VPWR VPWR _05614_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_128_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12717_ _02654_ _02655_ VGND VGND VPWR VPWR _02656_ sky130_fd_sc_hd__nor2_1
X_19273_ clknet_4_6_0_clock _00069_ VGND VGND VPWR VPWR kp\[3\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_155_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16485_ _06686_ _06691_ VGND VGND VPWR VPWR _06692_ sky130_fd_sc_hd__xor2_1
XFILLER_0_57_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13697_ net105 _03661_ _03656_ _03660_ VGND VGND VPWR VPWR _03663_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_84_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18224_ _08513_ _08518_ _08516_ VGND VGND VPWR VPWR _08605_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_150_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15436_ _05449_ _05454_ VGND VGND VPWR VPWR _05538_ sky130_fd_sc_hd__xnor2_1
X_12648_ _02585_ _02586_ VGND VGND VPWR VPWR _02587_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18155_ i_error\[15\] _08528_ VGND VGND VPWR VPWR _08529_ sky130_fd_sc_hd__nand2_1
X_15367_ _05373_ _05375_ _05365_ VGND VGND VPWR VPWR _05462_ sky130_fd_sc_hd__a21oi_1
X_12579_ _02479_ _02482_ VGND VGND VPWR VPWR _02518_ sky130_fd_sc_hd__nand2_1
X_17106_ _07373_ _07374_ VGND VGND VPWR VPWR _07375_ sky130_fd_sc_hd__or2_1
X_14318_ net451 net123 net120 net456 VGND VGND VPWR VPWR _04308_ sky130_fd_sc_hd__a22oi_1
X_18086_ _07346_ _07347_ _07350_ VGND VGND VPWR VPWR _08453_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15298_ _05357_ _05359_ _05337_ VGND VGND VPWR VPWR _05386_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17037_ net325 _06351_ _06344_ net320 VGND VGND VPWR VPWR _07299_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14249_ net438 net136 net132 net443 VGND VGND VPWR VPWR _04232_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_68_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09790_ _04929_ _05017_ _05028_ VGND VGND VPWR VPWR _05039_ sky130_fd_sc_hd__a21o_1
X_18988_ _09359_ _09444_ VGND VGND VPWR VPWR _09445_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17939_ _08282_ _08272_ _08281_ VGND VGND VPWR VPWR _08291_ sky130_fd_sc_hd__nor3_1
XFILLER_0_96_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09988_ _05941_ _06414_ _06403_ VGND VGND VPWR VPWR _07217_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_150_Right_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11950_ _01880_ _01888_ VGND VGND VPWR VPWR _01889_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10901_ _00833_ _00839_ VGND VGND VPWR VPWR _00840_ sky130_fd_sc_hd__or2b_1
XFILLER_0_86_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11881_ _01809_ _01819_ VGND VGND VPWR VPWR _01820_ sky130_fd_sc_hd__xor2_1
X_13620_ _03532_ _03578_ VGND VGND VPWR VPWR _03579_ sky130_fd_sc_hd__and2b_1
X_10832_ net379 net375 _05985_ _06183_ VGND VGND VPWR VPWR _00771_ sky130_fd_sc_hd__and4_1
XFILLER_0_149_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13551_ _03506_ _03508_ VGND VGND VPWR VPWR _03510_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10763_ net351 _00325_ VGND VGND VPWR VPWR _00702_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12502_ _02370_ _02374_ VGND VGND VPWR VPWR _02441_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16270_ net283 _06410_ VGND VGND VPWR VPWR _06455_ sky130_fd_sc_hd__nand2_1
X_13482_ _03436_ _03440_ VGND VGND VPWR VPWR _03441_ sky130_fd_sc_hd__nor2_1
X_10694_ _00535_ _00541_ VGND VGND VPWR VPWR _00633_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_81_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15221_ _05263_ _05300_ VGND VGND VPWR VPWR _05301_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12433_ net242 _01813_ VGND VGND VPWR VPWR _02372_ sky130_fd_sc_hd__nand2_2
XFILLER_0_152_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15152_ _05213_ _05222_ _05224_ VGND VGND VPWR VPWR _05225_ sky130_fd_sc_hd__a21o_1
X_12364_ _02279_ _02302_ VGND VGND VPWR VPWR _02303_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14103_ _04071_ _04074_ VGND VGND VPWR VPWR _04075_ sky130_fd_sc_hd__xnor2_1
X_11315_ _01252_ _01253_ VGND VGND VPWR VPWR _01254_ sky130_fd_sc_hd__xnor2_1
X_15083_ net423 net189 VGND VGND VPWR VPWR _05150_ sky130_fd_sc_hd__nand2_1
X_12295_ net199 _02210_ _02232_ _02233_ VGND VGND VPWR VPWR _02234_ sky130_fd_sc_hd__a31oi_1
X_14034_ _04004_ _04005_ net407 net151 VGND VGND VPWR VPWR _04006_ sky130_fd_sc_hd__and4bb_1
X_18911_ _09343_ _09344_ _09341_ VGND VGND VPWR VPWR _09360_ sky130_fd_sc_hd__o21ai_4
X_11246_ _01175_ _01176_ _01183_ VGND VGND VPWR VPWR _01185_ sky130_fd_sc_hd__nand3_1
X_18842_ _01848_ _01808_ VGND VGND VPWR VPWR _09284_ sky130_fd_sc_hd__or2_1
X_11177_ _00912_ _01031_ VGND VGND VPWR VPWR _01116_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10128_ _08724_ _08746_ VGND VGND VPWR VPWR _08757_ sky130_fd_sc_hd__and2_1
X_18773_ _08983_ _09207_ VGND VGND VPWR VPWR _09209_ sky130_fd_sc_hd__xnor2_1
X_15985_ _01679_ _01280_ VGND VGND VPWR VPWR _06142_ sky130_fd_sc_hd__xnor2_2
X_10059_ _05468_ _07987_ VGND VGND VPWR VPWR _07998_ sky130_fd_sc_hd__and2_1
X_14936_ _04930_ _04953_ _04947_ _04952_ VGND VGND VPWR VPWR _04988_ sky130_fd_sc_hd__a211o_1
X_17724_ _06539_ _08054_ _06800_ VGND VGND VPWR VPWR _08055_ sky130_fd_sc_hd__or3b_1
XFILLER_0_89_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14867_ _04902_ _04909_ _04911_ VGND VGND VPWR VPWR _04912_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17655_ net318 _06801_ VGND VGND VPWR VPWR _07979_ sky130_fd_sc_hd__nand2_1
X_16606_ _06823_ _06824_ VGND VGND VPWR VPWR _06825_ sky130_fd_sc_hd__or2_1
X_13818_ _03758_ _03783_ _03780_ VGND VGND VPWR VPWR _03784_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_147_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17586_ _07893_ _07901_ _07902_ VGND VGND VPWR VPWR _07903_ sky130_fd_sc_hd__a21o_1
X_14798_ _04833_ _04835_ VGND VGND VPWR VPWR _04836_ sky130_fd_sc_hd__and2b_1
XFILLER_0_57_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19325_ clknet_4_0_0_clock _00008_ VGND VGND VPWR VPWR kd_1\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16537_ _06671_ _06747_ _06670_ VGND VGND VPWR VPWR _06749_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13749_ _03672_ _03712_ _03714_ VGND VGND VPWR VPWR _03715_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19256_ clknet_4_10_0_clock _00138_ VGND VGND VPWR VPWR prev_d_error\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16468_ _06328_ _06367_ _06320_ net303 VGND VGND VPWR VPWR _06673_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_156_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15419_ _05492_ _05516_ _05518_ VGND VGND VPWR VPWR _05519_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_72_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18207_ _08513_ _08518_ VGND VGND VPWR VPWR _08586_ sky130_fd_sc_hd__xor2_2
XFILLER_0_143_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19187_ net498 net417 net487 _09591_ VGND VGND VPWR VPWR _00148_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16399_ _06595_ _06596_ VGND VGND VPWR VPWR _06597_ sky130_fd_sc_hd__xor2_1
XFILLER_0_115_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18138_ _08502_ _08509_ VGND VGND VPWR VPWR _08510_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_41_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18069_ net102 _08430_ net512 _08433_ VGND VGND VPWR VPWR _08434_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_111_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09911_ _06348_ _06337_ VGND VGND VPWR VPWR _06370_ sky130_fd_sc_hd__and2b_1
XFILLER_0_22_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09842_ net371 _05600_ _05578_ VGND VGND VPWR VPWR _05611_ sky130_fd_sc_hd__a21oi_1
X_09773_ _04159_ _04786_ _04830_ VGND VGND VPWR VPWR _04852_ sky130_fd_sc_hd__nand3_4
XFILLER_0_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_14_0_clock clknet_0_clock VGND VGND VPWR VPWR clknet_4_14_0_clock sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11100_ _01017_ _01037_ _00951_ _01038_ VGND VGND VPWR VPWR _01039_ sky130_fd_sc_hd__o211ai_2
X_12080_ _01846_ _02016_ _02018_ VGND VGND VPWR VPWR _02019_ sky130_fd_sc_hd__or3_1
XFILLER_0_130_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11031_ _00969_ _00567_ VGND VGND VPWR VPWR _00970_ sky130_fd_sc_hd__xnor2_4
X_15770_ _05879_ _05894_ _05904_ VGND VGND VPWR VPWR _05905_ sky130_fd_sc_hd__or3b_1
X_12982_ _02919_ _02920_ VGND VGND VPWR VPWR _02921_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14721_ _04749_ _04750_ VGND VGND VPWR VPWR _04751_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11933_ _01734_ _01871_ VGND VGND VPWR VPWR _01872_ sky130_fd_sc_hd__xor2_2
XFILLER_0_59_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17440_ _07266_ _07741_ VGND VGND VPWR VPWR _07742_ sky130_fd_sc_hd__and2_1
XFILLER_0_157_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14652_ _04673_ _04674_ VGND VGND VPWR VPWR _04675_ sky130_fd_sc_hd__nor2_1
X_11864_ _01792_ _01801_ VGND VGND VPWR VPWR _01803_ sky130_fd_sc_hd__and2_1
X_13603_ _03513_ _03512_ VGND VGND VPWR VPWR _03562_ sky130_fd_sc_hd__and2b_1
XFILLER_0_67_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17371_ net277 _02933_ VGND VGND VPWR VPWR _07666_ sky130_fd_sc_hd__nand2_1
X_10815_ _00663_ _00749_ _00753_ VGND VGND VPWR VPWR _00754_ sky130_fd_sc_hd__o21a_2
X_14583_ net121 _03912_ VGND VGND VPWR VPWR _04600_ sky130_fd_sc_hd__and2_1
X_11795_ _01708_ _01709_ _01732_ _01733_ VGND VGND VPWR VPWR _01734_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_27_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16322_ net273 _06346_ VGND VGND VPWR VPWR _06512_ sky130_fd_sc_hd__nand2_1
X_19110_ net500 prev_error\[16\] VGND VGND VPWR VPWR _09544_ sky130_fd_sc_hd__or2_1
X_13534_ _03458_ _03462_ _03492_ _03491_ _03464_ VGND VGND VPWR VPWR _03493_ sky130_fd_sc_hd__o32ai_4
XFILLER_0_138_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10746_ net371 _06623_ _00488_ VGND VGND VPWR VPWR _00685_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19041_ _09496_ _09497_ net493 VGND VGND VPWR VPWR _00081_ sky130_fd_sc_hd__o21a_1
X_16253_ _06435_ VGND VGND VPWR VPWR _06437_ sky130_fd_sc_hd__buf_4
X_13465_ _03341_ _03422_ VGND VGND VPWR VPWR _03424_ sky130_fd_sc_hd__or2_1
X_10677_ net343 _00409_ _00516_ kp\[16\] VGND VGND VPWR VPWR _00616_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15204_ _05165_ _05206_ _05264_ VGND VGND VPWR VPWR _05283_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12416_ _02249_ _02352_ _02347_ _02351_ VGND VGND VPWR VPWR _02355_ sky130_fd_sc_hd__a211oi_1
X_16184_ _06331_ _06332_ _06340_ _06360_ VGND VGND VPWR VPWR _06361_ sky130_fd_sc_hd__a31o_1
X_13396_ _03349_ _03350_ VGND VGND VPWR VPWR _03351_ sky130_fd_sc_hd__xor2_1
XFILLER_0_112_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15135_ _05123_ _05134_ _05133_ VGND VGND VPWR VPWR _05207_ sky130_fd_sc_hd__a21o_1
X_12347_ net230 _01807_ _02285_ VGND VGND VPWR VPWR _02286_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_2_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15066_ net453 net460 net163 net157 VGND VGND VPWR VPWR _05131_ sky130_fd_sc_hd__and4_1
X_12278_ net205 net203 _02091_ _01910_ VGND VGND VPWR VPWR _02217_ sky130_fd_sc_hd__and4_1
X_14017_ net425 net430 net141 net137 VGND VGND VPWR VPWR _03989_ sky130_fd_sc_hd__and4_1
X_11229_ _01114_ _01167_ VGND VGND VPWR VPWR _01168_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18825_ _09264_ _09265_ VGND VGND VPWR VPWR _09266_ sky130_fd_sc_hd__and2_1
XFILLER_0_156_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18756_ _09150_ _09165_ VGND VGND VPWR VPWR _09190_ sky130_fd_sc_hd__or2_1
X_15968_ _06015_ _06017_ VGND VGND VPWR VPWR _06123_ sky130_fd_sc_hd__and2_1
X_17707_ _08034_ _08035_ VGND VGND VPWR VPWR _08036_ sky130_fd_sc_hd__or2_1
X_14919_ _04820_ _04968_ VGND VGND VPWR VPWR _04969_ sky130_fd_sc_hd__xnor2_1
X_15899_ _03868_ _03087_ _03866_ VGND VGND VPWR VPWR _06047_ sky130_fd_sc_hd__nand3_1
X_18687_ _09075_ _09077_ _09113_ VGND VGND VPWR VPWR _09114_ sky130_fd_sc_hd__a21o_1
X_17638_ _07868_ _07869_ _07871_ VGND VGND VPWR VPWR _07960_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17569_ _07798_ _07883_ VGND VGND VPWR VPWR _07884_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19308_ clknet_4_1_0_clock _00000_ VGND VGND VPWR VPWR kd_1\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19239_ clknet_4_9_0_clock _00121_ VGND VGND VPWR VPWR i_error\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout402 net403 VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__buf_2
Xfanout413 net415 VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__buf_2
XFILLER_0_10_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout424 prev_d_error\[14\] VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__clkbuf_2
Xfanout435 prev_d_error\[11\] VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__buf_2
Xfanout446 net447 VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__clkbuf_4
Xfanout457 net458 VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__clkbuf_4
X_09825_ _05413_ VGND VGND VPWR VPWR _05424_ sky130_fd_sc_hd__buf_2
Xfanout468 prev_d_error\[4\] VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__clkbuf_4
Xfanout479 net480 VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__clkbuf_2
X_09756_ _04621_ _04522_ _04511_ VGND VGND VPWR VPWR _04665_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_68_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09687_ net40 _03881_ _03914_ net406 VGND VGND VPWR VPWR _00057_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10600_ net401 _05061_ _00537_ _00538_ VGND VGND VPWR VPWR _00539_ sky130_fd_sc_hd__nand4_1
X_11580_ _01472_ _01517_ _01518_ VGND VGND VPWR VPWR _01519_ sky130_fd_sc_hd__or3_1
XFILLER_0_119_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10531_ net383 _05182_ _00469_ _00468_ VGND VGND VPWR VPWR _00470_ sky130_fd_sc_hd__a31o_2
XFILLER_0_134_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13250_ _03133_ _03202_ VGND VGND VPWR VPWR _03203_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10462_ _00399_ _00400_ VGND VGND VPWR VPWR _00401_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12201_ _02138_ _02139_ VGND VGND VPWR VPWR _02140_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13181_ net211 _02915_ _03132_ VGND VGND VPWR VPWR _03133_ sky130_fd_sc_hd__nand3_1
XFILLER_0_33_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10393_ net350 _08207_ VGND VGND VPWR VPWR _00332_ sky130_fd_sc_hd__nand2_1
X_12132_ _02067_ _02068_ _02070_ VGND VGND VPWR VPWR _02071_ sky130_fd_sc_hd__and3_2
XFILLER_0_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16940_ _07157_ _07191_ net270 VGND VGND VPWR VPWR _07192_ sky130_fd_sc_hd__and3b_1
X_12063_ _02000_ _02001_ VGND VGND VPWR VPWR _02002_ sky130_fd_sc_hd__nand2_1
X_11014_ _00922_ _00952_ VGND VGND VPWR VPWR _00953_ sky130_fd_sc_hd__xor2_4
X_16871_ _07078_ _07080_ VGND VGND VPWR VPWR _07116_ sky130_fd_sc_hd__nor2_1
X_18610_ _06116_ _09025_ VGND VGND VPWR VPWR _09029_ sky130_fd_sc_hd__nand2_1
X_15822_ _05960_ _05961_ VGND VGND VPWR VPWR _05962_ sky130_fd_sc_hd__nand2_1
X_15753_ _05837_ _05857_ VGND VGND VPWR VPWR _05887_ sky130_fd_sc_hd__xor2_1
X_18541_ _08897_ _08952_ _08893_ _08739_ VGND VGND VPWR VPWR _08953_ sky130_fd_sc_hd__o2bb2a_1
X_12965_ _02901_ _02903_ VGND VGND VPWR VPWR _02904_ sky130_fd_sc_hd__and2_1
X_11916_ _01848_ _01854_ VGND VGND VPWR VPWR _01855_ sky130_fd_sc_hd__or2_1
X_14704_ _04729_ _04732_ VGND VGND VPWR VPWR _04733_ sky130_fd_sc_hd__and2_1
X_15684_ _05740_ _05800_ _05804_ _05810_ VGND VGND VPWR VPWR _05811_ sky130_fd_sc_hd__o31ai_4
X_18472_ net532 _08870_ _08872_ _08622_ _08615_ VGND VGND VPWR VPWR _08877_ sky130_fd_sc_hd__a32oi_1
X_12896_ _02809_ _02833_ _02730_ _02834_ VGND VGND VPWR VPWR _02835_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_68_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14635_ _04634_ _04639_ _04656_ VGND VGND VPWR VPWR _04657_ sky130_fd_sc_hd__a21oi_1
X_17423_ _07721_ _07722_ VGND VGND VPWR VPWR _07724_ sky130_fd_sc_hd__nand2_2
X_11847_ _01785_ VGND VGND VPWR VPWR _01786_ sky130_fd_sc_hd__buf_2
XFILLER_0_157_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14566_ _04556_ _04580_ _04553_ VGND VGND VPWR VPWR _04581_ sky130_fd_sc_hd__o21ai_1
X_17354_ _07254_ _07590_ _07647_ VGND VGND VPWR VPWR _07648_ sky130_fd_sc_hd__o21a_1
X_11778_ prev_error\[1\] _00813_ VGND VGND VPWR VPWR _01717_ sky130_fd_sc_hd__xnor2_4
X_13517_ _03474_ _03475_ VGND VGND VPWR VPWR _03476_ sky130_fd_sc_hd__nand2_1
X_16305_ _06492_ _06493_ VGND VGND VPWR VPWR _06494_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17285_ net281 _07565_ _07566_ net540 VGND VGND VPWR VPWR _07572_ sky130_fd_sc_hd__nand4_2
X_10729_ _00664_ _00666_ _00667_ VGND VGND VPWR VPWR _00668_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_126_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14497_ net439 net443 net147 net142 VGND VGND VPWR VPWR _04505_ sky130_fd_sc_hd__and4_1
XFILLER_0_82_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19024_ _09484_ VGND VGND VPWR VPWR _09485_ sky130_fd_sc_hd__buf_6
XFILLER_0_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16236_ net273 _06410_ VGND VGND VPWR VPWR _06418_ sky130_fd_sc_hd__nand2_1
X_13448_ _03390_ _03406_ VGND VGND VPWR VPWR _03407_ sky130_fd_sc_hd__xor2_1
X_16167_ _06341_ _06340_ VGND VGND VPWR VPWR _06342_ sky130_fd_sc_hd__xor2_1
X_13379_ _03272_ _03331_ VGND VGND VPWR VPWR _03332_ sky130_fd_sc_hd__xor2_1
XFILLER_0_51_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15118_ _05168_ _05185_ _05186_ _05187_ VGND VGND VPWR VPWR _05188_ sky130_fd_sc_hd__nor4_1
XFILLER_0_11_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16098_ _06265_ VGND VGND VPWR VPWR _06266_ sky130_fd_sc_hd__buf_2
XFILLER_0_11_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15049_ _05110_ _05106_ _05108_ VGND VGND VPWR VPWR _05112_ sky130_fd_sc_hd__or3_1
X_09610_ _03124_ VGND VGND VPWR VPWR _03135_ sky130_fd_sc_hd__buf_2
X_18808_ _04178_ _04182_ _09246_ VGND VGND VPWR VPWR _09247_ sky130_fd_sc_hd__a21o_1
X_18739_ _08961_ _09077_ _09170_ VGND VGND VPWR VPWR _09171_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout210 net212 VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_4
Xfanout221 net223 VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__buf_2
Xfanout232 net233 VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout243 net244 VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__clkbuf_4
Xfanout254 net255 VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__buf_2
Xfanout265 net266 VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__clkbuf_4
Xfanout276 net277 VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__clkbuf_4
X_09808_ net360 _05193_ _05226_ _05204_ VGND VGND VPWR VPWR _05237_ sky130_fd_sc_hd__a31o_1
Xfanout287 ki\[13\] VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__clkbuf_4
Xfanout298 ki\[9\] VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__clkbuf_4
X_09739_ _04379_ _04467_ VGND VGND VPWR VPWR _04478_ sky130_fd_sc_hd__or2_2
X_12750_ net250 _01813_ _01759_ net268 VGND VGND VPWR VPWR _02689_ sky130_fd_sc_hd__a22o_1
X_11701_ net564 _00516_ VGND VGND VPWR VPWR _01640_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12681_ _02612_ _02619_ VGND VGND VPWR VPWR _02620_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14420_ _04347_ _04419_ VGND VGND VPWR VPWR _04420_ sky130_fd_sc_hd__nor2_1
X_11632_ _01568_ _01570_ VGND VGND VPWR VPWR _01571_ sky130_fd_sc_hd__and2b_1
X_14351_ net425 net430 net152 net147 VGND VGND VPWR VPWR _04344_ sky130_fd_sc_hd__and4_1
XFILLER_0_37_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11563_ _01499_ _01498_ VGND VGND VPWR VPWR _01502_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13302_ _03251_ _03253_ _03254_ VGND VGND VPWR VPWR _03255_ sky130_fd_sc_hd__nand3_1
X_10514_ _00451_ _00433_ VGND VGND VPWR VPWR _00453_ sky130_fd_sc_hd__and2b_1
X_17070_ _07293_ _07290_ _06353_ _06364_ VGND VGND VPWR VPWR _07335_ sky130_fd_sc_hd__a2bb2o_1
X_14282_ _04263_ _04267_ VGND VGND VPWR VPWR _04268_ sky130_fd_sc_hd__and2_1
X_11494_ net400 _08196_ _01377_ _01378_ VGND VGND VPWR VPWR _01433_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16021_ kp\[16\] _05677_ VGND VGND VPWR VPWR _06181_ sky130_fd_sc_hd__and2_1
X_13233_ _03181_ _03185_ _03183_ VGND VGND VPWR VPWR _03186_ sky130_fd_sc_hd__o21ai_2
X_10445_ _00293_ _00382_ VGND VGND VPWR VPWR _00384_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13164_ _03110_ _03114_ VGND VGND VPWR VPWR _03115_ sky130_fd_sc_hd__xor2_1
X_10376_ _00288_ _00298_ _00286_ VGND VGND VPWR VPWR _00315_ sky130_fd_sc_hd__o21ai_1
X_12115_ net221 _01808_ VGND VGND VPWR VPWR _02054_ sky130_fd_sc_hd__nand2_1
X_13095_ _02904_ _03038_ VGND VGND VPWR VPWR _03039_ sky130_fd_sc_hd__or2_1
X_17972_ net326 _07156_ _08326_ VGND VGND VPWR VPWR _08327_ sky130_fd_sc_hd__and3_1
X_16923_ net288 _06890_ VGND VGND VPWR VPWR _07174_ sky130_fd_sc_hd__nand2_1
X_12046_ _01802_ _01821_ _01950_ VGND VGND VPWR VPWR _01985_ sky130_fd_sc_hd__nor3_1
X_16854_ _06989_ _07097_ VGND VGND VPWR VPWR _07098_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15805_ _05544_ _05614_ VGND VGND VPWR VPWR _05944_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_148_Left_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13997_ _03967_ _03968_ VGND VGND VPWR VPWR _03969_ sky130_fd_sc_hd__xnor2_1
X_16785_ _06938_ _06941_ VGND VGND VPWR VPWR _07022_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18524_ _06261_ _06264_ _08803_ VGND VGND VPWR VPWR _08935_ sky130_fd_sc_hd__a21oi_1
X_15736_ _05862_ _05867_ VGND VGND VPWR VPWR _05868_ sky130_fd_sc_hd__or2_1
X_12948_ net239 _01873_ VGND VGND VPWR VPWR _02887_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18455_ _06163_ _06165_ _06134_ VGND VGND VPWR VPWR _08859_ sky130_fd_sc_hd__o21ai_1
X_15667_ _05557_ _05791_ VGND VGND VPWR VPWR _05792_ sky130_fd_sc_hd__or2_1
X_12879_ net228 _02089_ VGND VGND VPWR VPWR _02818_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17406_ _07212_ _07226_ _07225_ VGND VGND VPWR VPWR _07705_ sky130_fd_sc_hd__o21a_1
XFILLER_0_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14618_ _04634_ _04637_ VGND VGND VPWR VPWR _04638_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15598_ _05596_ _05715_ VGND VGND VPWR VPWR _05716_ sky130_fd_sc_hd__or2_1
X_18386_ i_error\[5\] _08543_ VGND VGND VPWR VPWR _08783_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14549_ net409 net182 _04540_ _04541_ VGND VGND VPWR VPWR _04562_ sky130_fd_sc_hd__o2bb2a_1
X_17337_ _07618_ _07628_ VGND VGND VPWR VPWR _07629_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_157_Left_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17268_ net292 _07094_ _07552_ VGND VGND VPWR VPWR _07553_ sky130_fd_sc_hd__and3_1
X_19007_ _06146_ _09129_ VGND VGND VPWR VPWR _09466_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_114_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16219_ _06398_ VGND VGND VPWR VPWR _06399_ sky130_fd_sc_hd__clkbuf_4
X_17199_ _07469_ _07471_ _07475_ VGND VGND VPWR VPWR _07477_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10230_ _00166_ _00168_ VGND VGND VPWR VPWR _00169_ sky130_fd_sc_hd__nand2_1
X_10161_ _09098_ _09109_ VGND VGND VPWR VPWR _09120_ sky130_fd_sc_hd__nor2_2
XFILLER_0_100_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10092_ _08262_ _08339_ _08350_ VGND VGND VPWR VPWR _08361_ sky130_fd_sc_hd__o21ba_1
X_13920_ _02354_ _03887_ _03888_ VGND VGND VPWR VPWR _03889_ sky130_fd_sc_hd__a21o_1
X_13851_ _03801_ _03816_ VGND VGND VPWR VPWR _03817_ sky130_fd_sc_hd__nor2_1
X_12802_ net211 _02410_ _02740_ _02738_ VGND VGND VPWR VPWR _02741_ sky130_fd_sc_hd__a31o_1
X_13782_ net108 _03745_ _03738_ _03744_ VGND VGND VPWR VPWR _03748_ sky130_fd_sc_hd__o211a_1
X_16570_ _06763_ _06764_ VGND VGND VPWR VPWR _06785_ sky130_fd_sc_hd__xnor2_1
X_10994_ _00869_ _00873_ _00870_ VGND VGND VPWR VPWR _00933_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12733_ _02571_ _02671_ VGND VGND VPWR VPWR _02672_ sky130_fd_sc_hd__nor2_1
X_15521_ _05595_ _05596_ VGND VGND VPWR VPWR _05631_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15452_ _05550_ _05552_ _05554_ VGND VGND VPWR VPWR _05555_ sky130_fd_sc_hd__o21ai_1
X_18240_ _08620_ _08621_ VGND VGND VPWR VPWR _08622_ sky130_fd_sc_hd__nand2_2
X_12664_ _02484_ _02598_ _02602_ VGND VGND VPWR VPWR _02603_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14403_ _04400_ _04389_ VGND VGND VPWR VPWR _04402_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11615_ net399 _00323_ VGND VGND VPWR VPWR _01554_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15383_ _05477_ _05478_ net463 net172 VGND VGND VPWR VPWR _05480_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_93_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18171_ _08545_ net515 _07972_ VGND VGND VPWR VPWR _08546_ sky130_fd_sc_hd__a21oi_2
X_12595_ net217 net214 _02091_ _01909_ VGND VGND VPWR VPWR _02534_ sky130_fd_sc_hd__and4_1
XFILLER_0_108_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17122_ _07390_ _07391_ VGND VGND VPWR VPWR _07392_ sky130_fd_sc_hd__xor2_2
X_14334_ _04322_ _04325_ VGND VGND VPWR VPWR _04326_ sky130_fd_sc_hd__and2b_1
XFILLER_0_80_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11546_ net394 _01001_ _01376_ VGND VGND VPWR VPWR _01485_ sky130_fd_sc_hd__nand3_1
XFILLER_0_13_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17053_ _06537_ _06492_ _07287_ _07315_ VGND VGND VPWR VPWR _07317_ sky130_fd_sc_hd__o31ai_1
X_14265_ _04249_ VGND VGND VPWR VPWR _04250_ sky130_fd_sc_hd__inv_2
X_11477_ _01413_ _01415_ VGND VGND VPWR VPWR _01416_ sky130_fd_sc_hd__nand2_1
X_16004_ _06135_ _06159_ _06162_ VGND VGND VPWR VPWR _06163_ sky130_fd_sc_hd__or3_4
X_13216_ _03127_ _03168_ VGND VGND VPWR VPWR _03169_ sky130_fd_sc_hd__xnor2_1
X_10428_ net387 _00363_ net539 VGND VGND VPWR VPWR _00367_ sky130_fd_sc_hd__and3_1
X_14196_ _04172_ _04173_ VGND VGND VPWR VPWR _04174_ sky130_fd_sc_hd__and2_1
X_13147_ _03093_ _03095_ VGND VGND VPWR VPWR _03096_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10359_ _00235_ _00296_ _00297_ _00290_ _00295_ VGND VGND VPWR VPWR _00298_ sky130_fd_sc_hd__o32a_2
X_13078_ _02988_ _03004_ VGND VGND VPWR VPWR _03020_ sky130_fd_sc_hd__xor2_2
X_17955_ _08302_ _08308_ VGND VGND VPWR VPWR _08309_ sky130_fd_sc_hd__or2_1
X_12029_ _01855_ _01891_ _01890_ VGND VGND VPWR VPWR _01968_ sky130_fd_sc_hd__o21ba_1
X_16906_ _02637_ _06278_ VGND VGND VPWR VPWR _07155_ sky130_fd_sc_hd__xor2_4
X_17886_ net314 VGND VGND VPWR VPWR _08233_ sky130_fd_sc_hd__inv_2
X_16837_ _07055_ _07064_ _07065_ VGND VGND VPWR VPWR _07079_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16768_ _07002_ _07001_ VGND VGND VPWR VPWR _07003_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18507_ _08906_ _08910_ _08914_ _08915_ VGND VGND VPWR VPWR _08916_ sky130_fd_sc_hd__and4bb_1
X_15719_ _05845_ _05838_ _05843_ VGND VGND VPWR VPWR _05849_ sky130_fd_sc_hd__or3_1
X_16699_ _06839_ _06926_ VGND VGND VPWR VPWR _06927_ sky130_fd_sc_hd__xnor2_2
X_18438_ _08838_ _08839_ VGND VGND VPWR VPWR _08840_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18369_ _08763_ _08607_ VGND VGND VPWR VPWR _08764_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_90_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_131_Right_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11400_ _01310_ _01338_ VGND VGND VPWR VPWR _01339_ sky130_fd_sc_hd__nor2_1
X_12380_ net209 _01910_ _02318_ VGND VGND VPWR VPWR _02319_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11331_ _01265_ _01268_ _01190_ _01249_ VGND VGND VPWR VPWR _01270_ sky130_fd_sc_hd__a211o_1
XFILLER_0_6_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14050_ _03983_ VGND VGND VPWR VPWR _04022_ sky130_fd_sc_hd__inv_2
X_11262_ _01196_ _01197_ _01192_ _01195_ VGND VGND VPWR VPWR _01201_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_132_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13001_ _02923_ _02925_ _02939_ VGND VGND VPWR VPWR _02940_ sky130_fd_sc_hd__a21oi_1
X_10213_ _09546_ _09596_ VGND VGND VPWR VPWR _00152_ sky130_fd_sc_hd__nor2_1
X_11193_ _01040_ _01041_ _01039_ VGND VGND VPWR VPWR _01132_ sky130_fd_sc_hd__a21boi_4
X_10144_ _05666_ _08922_ VGND VGND VPWR VPWR _08933_ sky130_fd_sc_hd__xor2_1
XFILLER_0_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17740_ _08055_ _08057_ VGND VGND VPWR VPWR _08072_ sky130_fd_sc_hd__nand2_1
X_14952_ net467 net144 net124 net485 VGND VGND VPWR VPWR _05005_ sky130_fd_sc_hd__a22oi_2
X_10075_ _06579_ _08163_ VGND VGND VPWR VPWR _08174_ sky130_fd_sc_hd__nor2_1
X_13903_ _02772_ _02872_ VGND VGND VPWR VPWR _03871_ sky130_fd_sc_hd__or2_1
X_17671_ _07992_ _07994_ VGND VGND VPWR VPWR _07996_ sky130_fd_sc_hd__xnor2_2
X_14883_ _04912_ _04927_ _04928_ VGND VGND VPWR VPWR _04930_ sky130_fd_sc_hd__a21o_1
X_16622_ net312 _06545_ _06320_ _06364_ VGND VGND VPWR VPWR _06842_ sky130_fd_sc_hd__a31o_1
X_13834_ _03791_ _03796_ VGND VGND VPWR VPWR _03800_ sky130_fd_sc_hd__xnor2_1
X_19341_ clknet_4_0_0_clock _00024_ VGND VGND VPWR VPWR kd_2\[14\] sky130_fd_sc_hd__dfxtp_1
X_13765_ _02913_ _03730_ VGND VGND VPWR VPWR _03731_ sky130_fd_sc_hd__nand2_1
X_16553_ _06758_ _06765_ VGND VGND VPWR VPWR _06767_ sky130_fd_sc_hd__nor2_1
X_10977_ _00901_ _00914_ VGND VGND VPWR VPWR _00916_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15504_ _05548_ _05612_ VGND VGND VPWR VPWR _05613_ sky130_fd_sc_hd__nor2_1
X_12716_ _02646_ _02650_ _02653_ VGND VGND VPWR VPWR _02655_ sky130_fd_sc_hd__and3_1
X_19272_ clknet_4_6_0_clock _00068_ VGND VGND VPWR VPWR kp\[2\] sky130_fd_sc_hd__dfxtp_1
X_13696_ _03656_ _03660_ net105 _03661_ VGND VGND VPWR VPWR _03662_ sky130_fd_sc_hd__a211o_1
X_16484_ net293 _06346_ _06688_ _06690_ VGND VGND VPWR VPWR _06691_ sky130_fd_sc_hd__a31o_1
XFILLER_0_116_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18223_ _07154_ _08602_ VGND VGND VPWR VPWR _08604_ sky130_fd_sc_hd__and2_2
X_12647_ net246 _01814_ VGND VGND VPWR VPWR _02586_ sky130_fd_sc_hd__nand2_1
X_15435_ _05533_ _05536_ VGND VGND VPWR VPWR _05537_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15366_ _05452_ _05459_ _05460_ VGND VGND VPWR VPWR _05461_ sky130_fd_sc_hd__and3_1
X_18154_ _06836_ _08522_ VGND VGND VPWR VPWR _08528_ sky130_fd_sc_hd__xor2_2
X_12578_ _02512_ _02515_ _02516_ VGND VGND VPWR VPWR _02517_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17105_ _07372_ _07370_ VGND VGND VPWR VPWR _07374_ sky130_fd_sc_hd__and2b_1
XFILLER_0_25_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14317_ net451 net456 net123 net120 VGND VGND VPWR VPWR _04307_ sky130_fd_sc_hd__and4_1
XFILLER_0_41_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11529_ _01423_ _01426_ VGND VGND VPWR VPWR _01468_ sky130_fd_sc_hd__xor2_2
X_15297_ _05384_ _05368_ VGND VGND VPWR VPWR _05385_ sky130_fd_sc_hd__xnor2_1
X_18085_ _07772_ _07779_ VGND VGND VPWR VPWR _08452_ sky130_fd_sc_hd__and2b_1
XFILLER_0_151_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14248_ net438 net443 net136 net132 VGND VGND VPWR VPWR _04231_ sky130_fd_sc_hd__and4_1
X_17036_ net329 _06334_ VGND VGND VPWR VPWR _07298_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14179_ _03950_ _04047_ _04064_ VGND VGND VPWR VPWR _04155_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18987_ _09438_ _09443_ VGND VGND VPWR VPWR _09444_ sky130_fd_sc_hd__xnor2_1
X_17938_ _08286_ _08289_ VGND VGND VPWR VPWR _08290_ sky130_fd_sc_hd__xnor2_1
X_17869_ _08212_ _08213_ VGND VGND VPWR VPWR _08214_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_10_0_clock clknet_0_clock VGND VGND VPWR VPWR clknet_4_10_0_clock sky130_fd_sc_hd__clkbuf_8
XFILLER_0_31_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09987_ _06997_ _07195_ VGND VGND VPWR VPWR _07206_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10900_ _00834_ _00732_ _00835_ _00838_ VGND VGND VPWR VPWR _00839_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11880_ _01816_ _01818_ VGND VGND VPWR VPWR _01819_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10831_ net379 _05985_ _06183_ net375 VGND VGND VPWR VPWR _00770_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_67_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13550_ _03506_ _03508_ VGND VGND VPWR VPWR _03509_ sky130_fd_sc_hd__nand2_1
X_10762_ _00619_ _00621_ VGND VGND VPWR VPWR _00701_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12501_ _02270_ _02437_ _02439_ VGND VGND VPWR VPWR _02440_ sky130_fd_sc_hd__o21a_1
XFILLER_0_137_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13481_ _03371_ _03437_ _03439_ VGND VGND VPWR VPWR _03440_ sky130_fd_sc_hd__o21ba_1
X_10693_ _00576_ _00631_ VGND VGND VPWR VPWR _00632_ sky130_fd_sc_hd__nor2_2
X_15220_ _05258_ _05260_ _05262_ VGND VGND VPWR VPWR _05300_ sky130_fd_sc_hd__a21oi_1
X_12432_ net238 _01814_ _01798_ net242 VGND VGND VPWR VPWR _02371_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15151_ _05120_ _05223_ VGND VGND VPWR VPWR _05224_ sky130_fd_sc_hd__nand2_1
X_12363_ _02257_ _02278_ VGND VGND VPWR VPWR _02302_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14102_ _04072_ _04073_ VGND VGND VPWR VPWR _04074_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11314_ net381 _09577_ VGND VGND VPWR VPWR _01253_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15082_ _05146_ _05144_ VGND VGND VPWR VPWR _05148_ sky130_fd_sc_hd__xnor2_1
X_12294_ _02212_ _02231_ VGND VGND VPWR VPWR _02233_ sky130_fd_sc_hd__and2b_1
X_14033_ net411 net146 net141 net416 VGND VGND VPWR VPWR _04005_ sky130_fd_sc_hd__a22oi_1
X_18910_ _09345_ _09348_ _09358_ VGND VGND VPWR VPWR _09359_ sky130_fd_sc_hd__o21a_1
X_11245_ _01175_ _01176_ _01183_ VGND VGND VPWR VPWR _01184_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18841_ _02147_ _02155_ _09282_ VGND VGND VPWR VPWR _09283_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_38_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11176_ _01009_ _01082_ _01083_ _01098_ VGND VGND VPWR VPWR _01115_ sky130_fd_sc_hd__a31oi_2
X_10127_ net336 _08735_ _08713_ VGND VGND VPWR VPWR _08746_ sky130_fd_sc_hd__a21o_1
X_18772_ _08996_ _09206_ VGND VGND VPWR VPWR _09207_ sky130_fd_sc_hd__nand2_1
X_15984_ _01134_ _06140_ VGND VGND VPWR VPWR _06141_ sky130_fd_sc_hd__xnor2_4
X_17723_ net322 _06889_ VGND VGND VPWR VPWR _08054_ sky130_fd_sc_hd__nand2_1
X_10058_ _05270_ _05457_ VGND VGND VPWR VPWR _07987_ sky130_fd_sc_hd__nand2_1
X_14935_ _04851_ _04956_ _04986_ VGND VGND VPWR VPWR _04987_ sky130_fd_sc_hd__or3_2
XFILLER_0_145_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17654_ _07952_ _07958_ _07957_ VGND VGND VPWR VPWR _07978_ sky130_fd_sc_hd__o21a_1
X_14866_ _04840_ _04910_ VGND VGND VPWR VPWR _04911_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_121_Left_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16605_ _06753_ _06790_ VGND VGND VPWR VPWR _06824_ sky130_fd_sc_hd__xnor2_2
X_13817_ _03782_ VGND VGND VPWR VPWR _03783_ sky130_fd_sc_hd__inv_2
X_17585_ _07892_ _07890_ VGND VGND VPWR VPWR _07902_ sky130_fd_sc_hd__and2b_1
X_14797_ _04724_ _04834_ VGND VGND VPWR VPWR _04835_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19324_ clknet_4_0_0_clock _00007_ VGND VGND VPWR VPWR kd_1\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16536_ _06670_ _06671_ _06747_ VGND VGND VPWR VPWR _06748_ sky130_fd_sc_hd__nor3_1
X_13748_ _03707_ _03713_ VGND VGND VPWR VPWR _03714_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19255_ clknet_4_11_0_clock _00137_ VGND VGND VPWR VPWR prev_d_error\[4\] sky130_fd_sc_hd__dfxtp_1
X_16467_ _06654_ _06657_ VGND VGND VPWR VPWR _06672_ sky130_fd_sc_hd__xnor2_1
X_13679_ _03615_ _03613_ VGND VGND VPWR VPWR _03643_ sky130_fd_sc_hd__and2b_1
X_18206_ _08542_ _08579_ _08583_ _08584_ VGND VGND VPWR VPWR _08585_ sky130_fd_sc_hd__or4_4
X_15418_ _05433_ _05517_ VGND VGND VPWR VPWR _05518_ sky130_fd_sc_hd__nand2_1
X_19186_ net498 _08973_ VGND VGND VPWR VPWR _09591_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16398_ _06339_ _06338_ VGND VGND VPWR VPWR _06596_ sky130_fd_sc_hd__and2b_1
X_18137_ _08507_ _08508_ VGND VGND VPWR VPWR _08509_ sky130_fd_sc_hd__nor2_2
X_15349_ _05426_ _05433_ _05440_ _05441_ VGND VGND VPWR VPWR _05442_ sky130_fd_sc_hd__a211o_1
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_130_Left_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18068_ _08048_ _08431_ _08165_ _08052_ VGND VGND VPWR VPWR _08433_ sky130_fd_sc_hd__o22ai_4
X_09910_ _06337_ _06348_ VGND VGND VPWR VPWR _06359_ sky130_fd_sc_hd__and2b_1
X_17019_ net320 net270 _06352_ VGND VGND VPWR VPWR _07279_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09841_ _05072_ VGND VGND VPWR VPWR _05600_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09772_ _04159_ _04786_ _04830_ VGND VGND VPWR VPWR _04841_ sky130_fd_sc_hd__a21o_2
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11030_ net388 _05985_ VGND VGND VPWR VPWR _00969_ sky130_fd_sc_hd__nand2_2
XFILLER_0_99_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12981_ net216 _02544_ _02409_ net220 VGND VGND VPWR VPWR _02920_ sky130_fd_sc_hd__a22oi_1
X_14720_ _04736_ _04738_ _04748_ VGND VGND VPWR VPWR _04750_ sky130_fd_sc_hd__nand3_1
X_11932_ prev_error\[10\] _06172_ VGND VGND VPWR VPWR _01871_ sky130_fd_sc_hd__xor2_4
XFILLER_0_115_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11863_ _01792_ _01801_ VGND VGND VPWR VPWR _01802_ sky130_fd_sc_hd__nor2_1
X_14651_ _04669_ _04672_ VGND VGND VPWR VPWR _04674_ sky130_fd_sc_hd__and2_1
XFILLER_0_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13602_ net237 _02747_ VGND VGND VPWR VPWR _03561_ sky130_fd_sc_hd__nand2_1
X_10814_ _00750_ _00752_ VGND VGND VPWR VPWR _00753_ sky130_fd_sc_hd__or2b_1
X_17370_ net280 _07570_ VGND VGND VPWR VPWR _07665_ sky130_fd_sc_hd__nand2_1
X_14582_ net470 net121 net118 net475 VGND VGND VPWR VPWR _04598_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_83_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11794_ _06590_ _06601_ prev_error\[9\] VGND VGND VPWR VPWR _01733_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_156_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16321_ _06495_ _06498_ _06497_ VGND VGND VPWR VPWR _06511_ sky130_fd_sc_hd__o21ai_1
X_13533_ _03464_ _03491_ VGND VGND VPWR VPWR _03492_ sky130_fd_sc_hd__xnor2_2
X_10745_ _00683_ VGND VGND VPWR VPWR _00684_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19040_ net522 _09485_ _09462_ VGND VGND VPWR VPWR _09497_ sky130_fd_sc_hd__a21oi_1
X_13464_ _03341_ _03422_ VGND VGND VPWR VPWR _03423_ sky130_fd_sc_hd__nand2_1
X_16252_ _06431_ _06434_ VGND VGND VPWR VPWR _06435_ sky130_fd_sc_hd__and2_1
X_10676_ _00614_ VGND VGND VPWR VPWR _00615_ sky130_fd_sc_hd__buf_4
XFILLER_0_152_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12415_ _02256_ _02353_ VGND VGND VPWR VPWR _02354_ sky130_fd_sc_hd__nand2_1
X_15203_ _05279_ _05280_ VGND VGND VPWR VPWR _05282_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13395_ net258 _02088_ VGND VGND VPWR VPWR _03350_ sky130_fd_sc_hd__nand2_1
X_16183_ _06342_ _06358_ VGND VGND VPWR VPWR _06360_ sky130_fd_sc_hd__and2b_1
XFILLER_0_23_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12346_ net227 _01835_ VGND VGND VPWR VPWR _02285_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15134_ _05162_ _05163_ _05164_ _05140_ VGND VGND VPWR VPWR _05206_ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15065_ net449 net166 VGND VGND VPWR VPWR _05130_ sky130_fd_sc_hd__nand2_1
X_12277_ _02092_ _02094_ VGND VGND VPWR VPWR _02216_ sky130_fd_sc_hd__xnor2_1
X_14016_ _03954_ _03987_ VGND VGND VPWR VPWR _03988_ sky130_fd_sc_hd__and2_1
X_11228_ _01111_ _01113_ VGND VGND VPWR VPWR _01167_ sky130_fd_sc_hd__or2_1
X_18824_ _04202_ _04204_ _04206_ VGND VGND VPWR VPWR _09265_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_156_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11159_ _01085_ _01097_ VGND VGND VPWR VPWR _01098_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18755_ _09185_ _09187_ _09188_ VGND VGND VPWR VPWR _09189_ sky130_fd_sc_hd__a21oi_2
X_15967_ _06021_ _06022_ _06121_ VGND VGND VPWR VPWR _06122_ sky130_fd_sc_hd__a21oi_4
X_17706_ _07924_ _07948_ VGND VGND VPWR VPWR _08035_ sky130_fd_sc_hd__xnor2_2
X_14918_ _04897_ _04898_ VGND VGND VPWR VPWR _04968_ sky130_fd_sc_hd__nor2_1
X_18686_ _08792_ _09112_ _08881_ VGND VGND VPWR VPWR _09113_ sky130_fd_sc_hd__mux2_1
X_15898_ _06043_ _06045_ VGND VGND VPWR VPWR _06046_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17637_ _07952_ _07957_ _07958_ VGND VGND VPWR VPWR _07959_ sky130_fd_sc_hd__nor3_2
X_14849_ _04783_ _04782_ VGND VGND VPWR VPWR _04892_ sky130_fd_sc_hd__xor2_1
XFILLER_0_148_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17568_ _07799_ _07881_ _07882_ VGND VGND VPWR VPWR _07883_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_74_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19307_ clknet_4_7_0_clock _00047_ VGND VGND VPWR VPWR ki\[18\] sky130_fd_sc_hd__dfxtp_2
X_16519_ _06727_ _06728_ VGND VGND VPWR VPWR _06729_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17499_ _07804_ _07806_ VGND VGND VPWR VPWR _07807_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19238_ clknet_4_13_0_clock _00120_ VGND VGND VPWR VPWR i_error\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19169_ _09550_ _09144_ _09580_ net491 VGND VGND VPWR VPWR _00139_ sky130_fd_sc_hd__o211a_1
XFILLER_0_143_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout403 kp\[1\] VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__clkbuf_4
Xfanout414 net415 VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__clkbuf_2
Xfanout425 net426 VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__buf_2
Xfanout436 prev_d_error\[11\] VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__clkbuf_4
Xfanout447 prev_d_error\[9\] VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__buf_2
X_09824_ _05402_ VGND VGND VPWR VPWR _05413_ sky130_fd_sc_hd__buf_2
Xfanout458 net460 VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__buf_2
Xfanout469 net470 VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__buf_2
X_09755_ _04423_ _04500_ _04533_ _04610_ _04643_ VGND VGND VPWR VPWR _04654_ sky130_fd_sc_hd__a2111oi_4
X_09686_ _03903_ VGND VGND VPWR VPWR _03914_ sky130_fd_sc_hd__buf_2
XFILLER_0_139_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout10 net355 VGND VGND VPWR VPWR net565 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10530_ _00467_ _00468_ VGND VGND VPWR VPWR _00469_ sky130_fd_sc_hd__nor2_2
XFILLER_0_17_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10461_ net354 _08196_ _06634_ net356 VGND VGND VPWR VPWR _00400_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_122_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12200_ _02123_ _02124_ _02137_ VGND VGND VPWR VPWR _02139_ sky130_fd_sc_hd__nand3_1
XFILLER_0_134_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13180_ _03130_ _03131_ VGND VGND VPWR VPWR _03132_ sky130_fd_sc_hd__and2_1
X_10392_ _00329_ _00330_ VGND VGND VPWR VPWR _00331_ sky130_fd_sc_hd__xor2_1
X_12131_ _02045_ _02069_ VGND VGND VPWR VPWR _02070_ sky130_fd_sc_hd__nor2_1
X_12062_ _01936_ _01945_ _01999_ VGND VGND VPWR VPWR _02001_ sky130_fd_sc_hd__or3_1
X_11013_ _00948_ _00951_ VGND VGND VPWR VPWR _00952_ sky130_fd_sc_hd__and2_2
X_16870_ _07112_ _07110_ VGND VGND VPWR VPWR _07115_ sky130_fd_sc_hd__xnor2_1
X_15821_ _05959_ _05100_ _05957_ VGND VGND VPWR VPWR _05961_ sky130_fd_sc_hd__nand3_1
XFILLER_0_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18540_ _08750_ net100 _08951_ _08902_ VGND VGND VPWR VPWR _08952_ sky130_fd_sc_hd__a211o_1
X_15752_ _05882_ _05884_ VGND VGND VPWR VPWR _05885_ sky130_fd_sc_hd__nor2_1
X_12964_ _02844_ _02902_ VGND VGND VPWR VPWR _02903_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14703_ _04561_ _04730_ VGND VGND VPWR VPWR _04732_ sky130_fd_sc_hd__nor2_1
X_11915_ _01853_ VGND VGND VPWR VPWR _01854_ sky130_fd_sc_hd__buf_2
X_18471_ _08767_ _08869_ _08873_ _08874_ _08875_ VGND VGND VPWR VPWR _08876_ sky130_fd_sc_hd__a2111o_1
X_15683_ _05806_ _05808_ VGND VGND VPWR VPWR _05810_ sky130_fd_sc_hd__nand2_1
X_12895_ _02711_ _02729_ _02728_ VGND VGND VPWR VPWR _02834_ sky130_fd_sc_hd__a21o_1
X_17422_ _07720_ _07719_ VGND VGND VPWR VPWR _07722_ sky130_fd_sc_hd__or2b_1
X_14634_ _04653_ _04655_ VGND VGND VPWR VPWR _04656_ sky130_fd_sc_hd__or2b_1
X_11846_ _01784_ _01752_ VGND VGND VPWR VPWR _01785_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_55_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17353_ net288 _06993_ _07095_ net285 VGND VGND VPWR VPWR _07647_ sky130_fd_sc_hd__a22o_1
X_14565_ _04557_ _04579_ _04576_ VGND VGND VPWR VPWR _04580_ sky130_fd_sc_hd__a21oi_1
X_11777_ prev_error\[0\] _04236_ _00808_ VGND VGND VPWR VPWR _01716_ sky130_fd_sc_hd__nand3_4
XFILLER_0_67_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16304_ net292 _06378_ VGND VGND VPWR VPWR _06493_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13516_ _03471_ _03469_ VGND VGND VPWR VPWR _03475_ sky130_fd_sc_hd__xnor2_1
X_10728_ net401 _00363_ _04984_ VGND VGND VPWR VPWR _00667_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17284_ _07570_ VGND VGND VPWR VPWR _07571_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14496_ _04413_ _04503_ VGND VGND VPWR VPWR _04504_ sky130_fd_sc_hd__nor2_1
X_19023_ _09482_ VGND VGND VPWR VPWR _09484_ sky130_fd_sc_hd__clkbuf_2
X_16235_ net283 _06386_ _06391_ _06390_ VGND VGND VPWR VPWR _06417_ sky130_fd_sc_hd__a31o_1
X_13447_ _03402_ _03405_ _03400_ VGND VGND VPWR VPWR _03406_ sky130_fd_sc_hd__a21oi_1
X_10659_ _00579_ _00594_ _00596_ VGND VGND VPWR VPWR _00598_ sky130_fd_sc_hd__nand3_1
XFILLER_0_153_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13378_ _03305_ _03329_ _03330_ VGND VGND VPWR VPWR _03331_ sky130_fd_sc_hd__a21boi_1
X_16166_ _06331_ _06332_ VGND VGND VPWR VPWR _06341_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15117_ _05167_ _05140_ net114 VGND VGND VPWR VPWR _05187_ sky130_fd_sc_hd__nor3_1
X_12329_ net234 _01817_ _02266_ _02267_ VGND VGND VPWR VPWR _02268_ sky130_fd_sc_hd__a31o_1
X_16097_ _06261_ _06264_ VGND VGND VPWR VPWR _06265_ sky130_fd_sc_hd__and2_4
X_15048_ _05106_ _05108_ _05110_ VGND VGND VPWR VPWR _05111_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18807_ _09228_ _09245_ VGND VGND VPWR VPWR _09246_ sky130_fd_sc_hd__xnor2_1
X_16999_ _07254_ _07256_ VGND VGND VPWR VPWR _07257_ sky130_fd_sc_hd__nor2_2
X_18738_ _08819_ _09169_ _08880_ VGND VGND VPWR VPWR _09170_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18669_ _06094_ _06083_ _06092_ VGND VGND VPWR VPWR _09094_ sky130_fd_sc_hd__nand3_1
XFILLER_0_148_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout200 net201 VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__buf_2
XFILLER_0_100_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout211 net212 VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__buf_2
Xfanout222 net223 VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout233 kd_1\[9\] VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__buf_2
Xfanout244 net245 VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__clkbuf_4
Xfanout255 net257 VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout266 kd_1\[1\] VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__clkbuf_4
X_09807_ _05204_ _05215_ VGND VGND VPWR VPWR _05226_ sky130_fd_sc_hd__nor2_1
Xfanout277 ki\[16\] VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__buf_2
Xfanout288 ki\[12\] VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__clkbuf_4
Xfanout299 ki\[9\] VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__buf_4
X_09738_ _04434_ _04445_ _04456_ VGND VGND VPWR VPWR _04467_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09669_ net56 _03625_ _03658_ net307 VGND VGND VPWR VPWR _00054_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11700_ net394 _00811_ _01638_ VGND VGND VPWR VPWR _01639_ sky130_fd_sc_hd__and3_1
X_12680_ net227 _01853_ _02615_ _02618_ VGND VGND VPWR VPWR _02619_ sky130_fd_sc_hd__a31o_1
XFILLER_0_49_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11631_ _01563_ _01569_ VGND VGND VPWR VPWR _01570_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_145_Right_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14350_ _04318_ _04341_ _04342_ VGND VGND VPWR VPWR _04343_ sky130_fd_sc_hd__a21o_1
X_11562_ _01476_ _01478_ VGND VGND VPWR VPWR _01501_ sky130_fd_sc_hd__xor2_1
XFILLER_0_108_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13301_ _03159_ _03250_ _03246_ _03249_ VGND VGND VPWR VPWR _03254_ sky130_fd_sc_hd__a211o_1
XFILLER_0_80_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10513_ _00433_ _00451_ VGND VGND VPWR VPWR _00452_ sky130_fd_sc_hd__xnor2_1
X_14281_ _04257_ _04260_ _04262_ VGND VGND VPWR VPWR _04267_ sky130_fd_sc_hd__or3_1
X_11493_ _01373_ _01381_ VGND VGND VPWR VPWR _01432_ sky130_fd_sc_hd__xnor2_1
X_16020_ net339 _05193_ VGND VGND VPWR VPWR _06180_ sky130_fd_sc_hd__nand2_1
X_13232_ _03183_ _03184_ VGND VGND VPWR VPWR _03185_ sky130_fd_sc_hd__nand2_1
X_10444_ _00293_ _00382_ VGND VGND VPWR VPWR _00383_ sky130_fd_sc_hd__and2_1
XFILLER_0_150_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13163_ net225 _02545_ _03111_ _03112_ VGND VGND VPWR VPWR _03114_ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10375_ _00299_ _00312_ _00313_ VGND VGND VPWR VPWR _00314_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_131_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12114_ net230 net226 _01814_ _01799_ VGND VGND VPWR VPWR _02053_ sky130_fd_sc_hd__nand4_2
XFILLER_0_130_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13094_ _02901_ _02903_ VGND VGND VPWR VPWR _03038_ sky130_fd_sc_hd__nor2_1
X_17971_ _08324_ _08325_ VGND VGND VPWR VPWR _08326_ sky130_fd_sc_hd__nor2_1
X_16922_ _07164_ _07171_ VGND VGND VPWR VPWR _07172_ sky130_fd_sc_hd__xnor2_1
X_12045_ _01983_ VGND VGND VPWR VPWR _01984_ sky130_fd_sc_hd__clkbuf_2
X_16853_ net276 _06993_ VGND VGND VPWR VPWR _07097_ sky130_fd_sc_hd__nand2_1
X_15804_ _05675_ _05942_ VGND VGND VPWR VPWR _05943_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16784_ _06492_ _06540_ _07014_ _07020_ VGND VGND VPWR VPWR _07021_ sky130_fd_sc_hd__o22a_1
X_13996_ _03928_ _03927_ VGND VGND VPWR VPWR _03968_ sky130_fd_sc_hd__and2b_1
X_18523_ _08819_ _08924_ VGND VGND VPWR VPWR _08934_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15735_ _05860_ _05861_ VGND VGND VPWR VPWR _05867_ sky130_fd_sc_hd__and2_1
X_12947_ net244 net239 _01852_ _01873_ VGND VGND VPWR VPWR _02886_ sky130_fd_sc_hd__and4_1
X_18454_ _08587_ _08857_ VGND VGND VPWR VPWR _08858_ sky130_fd_sc_hd__xor2_2
X_15666_ net484 net187 VGND VGND VPWR VPWR _05791_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12878_ net236 _01907_ _02615_ VGND VGND VPWR VPWR _02817_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17405_ net305 _06437_ VGND VGND VPWR VPWR _07704_ sky130_fd_sc_hd__nand2_1
X_14617_ _04612_ _04633_ VGND VGND VPWR VPWR _04637_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11829_ _01767_ VGND VGND VPWR VPWR _01768_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_8_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18385_ net518 _08568_ _08569_ VGND VGND VPWR VPWR _08782_ sky130_fd_sc_hd__a21o_1
X_15597_ net442 net195 net192 net447 VGND VGND VPWR VPWR _05715_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_145_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17336_ _07619_ _07627_ VGND VGND VPWR VPWR _07628_ sky130_fd_sc_hd__xor2_1
X_14548_ _04559_ _04560_ net421 net170 VGND VGND VPWR VPWR _04561_ sky130_fd_sc_hd__and4bb_1
XPHY_EDGE_ROW_112_Right_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17267_ _07550_ _07551_ VGND VGND VPWR VPWR _07552_ sky130_fd_sc_hd__xor2_1
X_14479_ _04484_ _04483_ VGND VGND VPWR VPWR _04485_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19006_ net508 _09179_ VGND VGND VPWR VPWR _09465_ sky130_fd_sc_hd__xor2_2
X_16218_ net270 VGND VGND VPWR VPWR _06398_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_11_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17198_ _07469_ _07471_ _07475_ VGND VGND VPWR VPWR _07476_ sky130_fd_sc_hd__nand3_1
XFILLER_0_140_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16149_ _06313_ _06307_ _01757_ VGND VGND VPWR VPWR _06322_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10160_ _09076_ _09087_ VGND VGND VPWR VPWR _09109_ sky130_fd_sc_hd__and2_1
X_10091_ _08284_ _08317_ _08328_ VGND VGND VPWR VPWR _08350_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13850_ _03799_ _03800_ VGND VGND VPWR VPWR _03816_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12801_ _02738_ _02739_ VGND VGND VPWR VPWR _02740_ sky130_fd_sc_hd__nor2_1
X_13781_ _03739_ _03741_ VGND VGND VPWR VPWR _03747_ sky130_fd_sc_hd__nand2_1
X_10993_ _00869_ _00873_ _00870_ VGND VGND VPWR VPWR _00932_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15520_ _05627_ _05629_ VGND VGND VPWR VPWR _05630_ sky130_fd_sc_hd__or2b_1
XFILLER_0_85_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12732_ _02573_ _02667_ _02670_ VGND VGND VPWR VPWR _02671_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15451_ _05473_ _05553_ VGND VGND VPWR VPWR _05554_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12663_ _02599_ _02601_ VGND VGND VPWR VPWR _02602_ sky130_fd_sc_hd__or2b_1
XFILLER_0_84_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14402_ net461 net120 _03910_ VGND VGND VPWR VPWR _04400_ sky130_fd_sc_hd__a21oi_1
X_11614_ _01551_ _01552_ VGND VGND VPWR VPWR _01553_ sky130_fd_sc_hd__xor2_1
X_18170_ _07971_ _07970_ _07969_ VGND VGND VPWR VPWR _08545_ sky130_fd_sc_hd__a21bo_1
X_15382_ prev_d_error\[4\] net166 net148 net486 VGND VGND VPWR VPWR _05478_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_154_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12594_ _02405_ _02414_ _02415_ VGND VGND VPWR VPWR _02533_ sky130_fd_sc_hd__or3_1
X_17121_ _07133_ _07136_ VGND VGND VPWR VPWR _07391_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14333_ _04233_ _04323_ VGND VGND VPWR VPWR _04325_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11545_ _00964_ _00226_ _01435_ _01434_ VGND VGND VPWR VPWR _01484_ sky130_fd_sc_hd__or4b_1
XFILLER_0_123_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17052_ net321 _06335_ _07119_ VGND VGND VPWR VPWR _07315_ sky130_fd_sc_hd__nand3_1
X_14264_ _04245_ _04246_ _04238_ _04242_ VGND VGND VPWR VPWR _04249_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_12_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11476_ net381 _00409_ _01413_ _01414_ VGND VGND VPWR VPWR _01415_ sky130_fd_sc_hd__nand4_1
XFILLER_0_40_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16003_ _00866_ _06160_ VGND VGND VPWR VPWR _06162_ sky130_fd_sc_hd__xnor2_4
X_10427_ net383 _04841_ _04852_ VGND VGND VPWR VPWR _00366_ sky130_fd_sc_hd__and3_2
X_13215_ _03128_ _03137_ VGND VGND VPWR VPWR _03168_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14195_ _04132_ _04134_ _04171_ VGND VGND VPWR VPWR _04173_ sky130_fd_sc_hd__or3_1
XFILLER_0_110_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13146_ net252 _03094_ _01812_ VGND VGND VPWR VPWR _03095_ sky130_fd_sc_hd__and3_1
X_10358_ net350 _06645_ _00234_ VGND VGND VPWR VPWR _00297_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13077_ _03017_ _03018_ VGND VGND VPWR VPWR _03019_ sky130_fd_sc_hd__nand2_1
X_17954_ _08303_ _08307_ VGND VGND VPWR VPWR _08308_ sky130_fd_sc_hd__xnor2_2
X_10289_ _00152_ _00153_ VGND VGND VPWR VPWR _00228_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12028_ _01952_ _01966_ VGND VGND VPWR VPWR _01967_ sky130_fd_sc_hd__xnor2_1
X_16905_ _07047_ _07153_ VGND VGND VPWR VPWR _07154_ sky130_fd_sc_hd__nand2_1
X_17885_ _08228_ _08231_ VGND VGND VPWR VPWR _08232_ sky130_fd_sc_hd__and2b_1
X_16836_ _07068_ _07072_ _07077_ VGND VGND VPWR VPWR _07078_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16767_ _06896_ _06979_ VGND VGND VPWR VPWR _07002_ sky130_fd_sc_hd__nand2_1
X_13979_ _03902_ _03907_ _03949_ VGND VGND VPWR VPWR _03951_ sky130_fd_sc_hd__or3_1
X_18506_ _08905_ _08858_ _08851_ _08907_ VGND VGND VPWR VPWR _08915_ sky130_fd_sc_hd__o2bb2a_1
X_15718_ _05847_ _05834_ VGND VGND VPWR VPWR _05848_ sky130_fd_sc_hd__xor2_1
XFILLER_0_75_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16698_ _06904_ _06925_ _06923_ VGND VGND VPWR VPWR _06926_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_76_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18437_ _06159_ _06162_ VGND VGND VPWR VPWR _08839_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15649_ _05756_ _05769_ _05771_ VGND VGND VPWR VPWR _05772_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18368_ _08596_ _08600_ VGND VGND VPWR VPWR _08763_ sky130_fd_sc_hd__nand2_2
XFILLER_0_113_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17319_ _07605_ _07607_ _07606_ VGND VGND VPWR VPWR _07609_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18299_ _08677_ _06589_ _06666_ VGND VGND VPWR VPWR _08687_ sky130_fd_sc_hd__or3_1
XFILLER_0_154_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_16_Left_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_25_Left_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11330_ _01190_ _01249_ _01265_ _01268_ VGND VGND VPWR VPWR _01269_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_104_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11261_ _01169_ _01199_ VGND VGND VPWR VPWR _01200_ sky130_fd_sc_hd__nor2_1
X_13000_ _02927_ _02937_ _02938_ VGND VGND VPWR VPWR _02939_ sky130_fd_sc_hd__a21oi_1
X_10212_ net338 _09583_ _09595_ VGND VGND VPWR VPWR _09596_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11192_ _00921_ _00953_ VGND VGND VPWR VPWR _01131_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_101_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10143_ _06920_ _08911_ VGND VGND VPWR VPWR _08922_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_118_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14951_ _04976_ _04978_ _04977_ VGND VGND VPWR VPWR _05004_ sky130_fd_sc_hd__a21o_1
X_10074_ _04643_ _04423_ _04500_ VGND VGND VPWR VPWR _08163_ sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_34_Left_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13902_ _03087_ _03866_ _03868_ VGND VGND VPWR VPWR _03869_ sky130_fd_sc_hd__a21o_1
X_17670_ _07992_ _07994_ VGND VGND VPWR VPWR _07995_ sky130_fd_sc_hd__and2_1
X_14882_ _04859_ _04879_ VGND VGND VPWR VPWR _04928_ sky130_fd_sc_hd__xnor2_1
X_16621_ _06840_ _06761_ VGND VGND VPWR VPWR _06841_ sky130_fd_sc_hd__xor2_1
X_13833_ _03797_ _03798_ VGND VGND VPWR VPWR _03799_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19340_ clknet_4_2_0_clock _00023_ VGND VGND VPWR VPWR kd_2\[13\] sky130_fd_sc_hd__dfxtp_1
X_16552_ _06763_ _06764_ VGND VGND VPWR VPWR _06765_ sky130_fd_sc_hd__and2b_1
X_13764_ _03728_ _03729_ VGND VGND VPWR VPWR _03730_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10976_ _00901_ _00914_ VGND VGND VPWR VPWR _00915_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15503_ _05605_ _05608_ _05610_ VGND VGND VPWR VPWR _05612_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_97_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12715_ _02646_ _02650_ _02653_ VGND VGND VPWR VPWR _02654_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19271_ clknet_4_6_0_clock _00067_ VGND VGND VPWR VPWR kp\[1\] sky130_fd_sc_hd__dfxtp_1
X_16483_ net296 _06353_ _06598_ VGND VGND VPWR VPWR _06690_ sky130_fd_sc_hd__and3_1
X_13695_ _03596_ _03599_ _03598_ VGND VGND VPWR VPWR _03661_ sky130_fd_sc_hd__o21a_1
XFILLER_0_127_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18222_ _07047_ _07153_ VGND VGND VPWR VPWR _08602_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15434_ _05529_ _05535_ VGND VGND VPWR VPWR _05536_ sky130_fd_sc_hd__or2_1
X_12646_ _01761_ _02584_ VGND VGND VPWR VPWR _02585_ sky130_fd_sc_hd__xor2_1
XFILLER_0_38_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18153_ i_error\[16\] _08525_ VGND VGND VPWR VPWR _08527_ sky130_fd_sc_hd__xnor2_2
X_15365_ _05385_ _05456_ VGND VGND VPWR VPWR _05460_ sky130_fd_sc_hd__or2_1
X_12577_ _02506_ _02510_ VGND VGND VPWR VPWR _02516_ sky130_fd_sc_hd__and2b_1
X_17104_ _07370_ _07372_ VGND VGND VPWR VPWR _07373_ sky130_fd_sc_hd__and2b_1
X_14316_ _03955_ _04305_ VGND VGND VPWR VPWR _04306_ sky130_fd_sc_hd__xnor2_1
X_11528_ _01464_ _01465_ _01466_ VGND VGND VPWR VPWR _01467_ sky130_fd_sc_hd__o21bai_1
X_18084_ _07770_ _07771_ VGND VGND VPWR VPWR _08451_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15296_ _05365_ _05366_ VGND VGND VPWR VPWR _05384_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17035_ _07289_ _07296_ VGND VGND VPWR VPWR _07297_ sky130_fd_sc_hd__xnor2_2
X_14247_ _04217_ _04229_ VGND VGND VPWR VPWR _04230_ sky130_fd_sc_hd__nand2_1
X_11459_ _01355_ _01386_ VGND VGND VPWR VPWR _01398_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14178_ _04151_ _04152_ _04092_ _04102_ VGND VGND VPWR VPWR _04154_ sky130_fd_sc_hd__a211o_1
X_13129_ _02987_ _03049_ _03075_ VGND VGND VPWR VPWR _03076_ sky130_fd_sc_hd__o21ba_1
X_18986_ _09442_ _09441_ _06261_ VGND VGND VPWR VPWR _09443_ sky130_fd_sc_hd__mux2_1
X_17937_ _08287_ _08288_ _08250_ VGND VGND VPWR VPWR _08289_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17868_ _08202_ _08203_ VGND VGND VPWR VPWR _08213_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_84_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16819_ _07056_ _07057_ VGND VGND VPWR VPWR _07059_ sky130_fd_sc_hd__xor2_2
XFILLER_0_17_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17799_ _08135_ _08136_ VGND VGND VPWR VPWR _08137_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09986_ _07173_ _07184_ VGND VGND VPWR VPWR _07195_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10830_ net371 _06634_ VGND VGND VPWR VPWR _00769_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10761_ _08086_ _00615_ VGND VGND VPWR VPWR _00700_ sky130_fd_sc_hd__nor2_2
XFILLER_0_94_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12500_ _02273_ _02438_ VGND VGND VPWR VPWR _02439_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13480_ net236 _02641_ _03438_ VGND VGND VPWR VPWR _03439_ sky130_fd_sc_hd__and3_1
X_10692_ _00575_ _00574_ VGND VGND VPWR VPWR _00631_ sky130_fd_sc_hd__and2b_1
XFILLER_0_109_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12431_ _02366_ _02369_ VGND VGND VPWR VPWR _02370_ sky130_fd_sc_hd__xnor2_1
X_15150_ _05113_ _05119_ VGND VGND VPWR VPWR _05223_ sky130_fd_sc_hd__or2_1
X_12362_ _02299_ _02300_ VGND VGND VPWR VPWR _02301_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14101_ net428 net433 net124 net119 VGND VGND VPWR VPWR _04073_ sky130_fd_sc_hd__and4_1
XFILLER_0_121_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11313_ _01216_ _01215_ VGND VGND VPWR VPWR _01252_ sky130_fd_sc_hd__and2b_1
X_12293_ _02212_ _02231_ VGND VGND VPWR VPWR _02232_ sky130_fd_sc_hd__xnor2_1
X_15081_ _05144_ _05146_ VGND VGND VPWR VPWR _05147_ sky130_fd_sc_hd__and2b_1
XFILLER_0_31_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14032_ net411 net416 net146 net141 VGND VGND VPWR VPWR _04004_ sky130_fd_sc_hd__and4_1
X_11244_ _01177_ _01181_ _01182_ VGND VGND VPWR VPWR _01183_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18840_ _01929_ _02154_ VGND VGND VPWR VPWR _09282_ sky130_fd_sc_hd__or2b_1
X_11175_ _01111_ _01113_ VGND VGND VPWR VPWR _01114_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_42_Left_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10126_ _05292_ _05303_ VGND VGND VPWR VPWR _08735_ sky130_fd_sc_hd__nand2_2
X_18771_ _09008_ _09022_ _09203_ _09205_ VGND VGND VPWR VPWR _09206_ sky130_fd_sc_hd__a31o_1
X_15983_ _01209_ _01681_ VGND VGND VPWR VPWR _06140_ sky130_fd_sc_hd__nor2_2
X_17722_ _08050_ _08051_ VGND VGND VPWR VPWR _08052_ sky130_fd_sc_hd__nand2_2
X_10057_ _05633_ _07965_ VGND VGND VPWR VPWR _07976_ sky130_fd_sc_hd__or2_1
X_14934_ _04826_ _04957_ _04980_ _04985_ VGND VGND VPWR VPWR _04986_ sky130_fd_sc_hd__a31oi_2
X_17653_ _07879_ _07968_ _07967_ VGND VGND VPWR VPWR _07977_ sky130_fd_sc_hd__o21ai_2
X_14865_ _04837_ _04839_ VGND VGND VPWR VPWR _04910_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16604_ _06795_ _06822_ VGND VGND VPWR VPWR _06823_ sky130_fd_sc_hd__xor2_2
X_13816_ _03780_ _03781_ VGND VGND VPWR VPWR _03782_ sky130_fd_sc_hd__or2_2
X_17584_ _07894_ _07900_ VGND VGND VPWR VPWR _07901_ sky130_fd_sc_hd__xnor2_2
X_14796_ net436 net161 _04722_ _04723_ VGND VGND VPWR VPWR _04834_ sky130_fd_sc_hd__o2bb2a_1
X_19323_ clknet_4_0_0_clock _00006_ VGND VGND VPWR VPWR kd_1\[15\] sky130_fd_sc_hd__dfxtp_1
X_16535_ _06741_ _06746_ VGND VGND VPWR VPWR _06747_ sky130_fd_sc_hd__nor2_2
X_13747_ _03672_ _03712_ VGND VGND VPWR VPWR _03713_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10959_ _08086_ _00818_ _00825_ VGND VGND VPWR VPWR _00898_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_128_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19254_ clknet_4_11_0_clock _00136_ VGND VGND VPWR VPWR prev_d_error\[3\] sky130_fd_sc_hd__dfxtp_2
X_16466_ _06646_ _06664_ VGND VGND VPWR VPWR _06671_ sky130_fd_sc_hd__xnor2_2
X_13678_ _03638_ _03641_ VGND VGND VPWR VPWR _03642_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18205_ _08580_ _08582_ i_error\[8\] VGND VGND VPWR VPWR _08584_ sky130_fd_sc_hd__a21oi_1
X_15417_ _05428_ _05432_ VGND VGND VPWR VPWR _05517_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12629_ _02470_ _02567_ VGND VGND VPWR VPWR _02568_ sky130_fd_sc_hd__nor2_1
X_19185_ net498 net424 net487 _09590_ VGND VGND VPWR VPWR _00147_ sky130_fd_sc_hd__o211a_1
X_16397_ net293 _06336_ VGND VGND VPWR VPWR _06595_ sky130_fd_sc_hd__nand2_1
X_18136_ _08505_ _08506_ VGND VGND VPWR VPWR _08508_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15348_ _05434_ _05436_ _05438_ VGND VGND VPWR VPWR _05441_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18067_ _08048_ _08431_ _08165_ _08052_ VGND VGND VPWR VPWR _08432_ sky130_fd_sc_hd__or4_4
XFILLER_0_110_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15279_ _05355_ _05357_ _05364_ VGND VGND VPWR VPWR _05365_ sky130_fd_sc_hd__a21oi_1
X_17018_ _07192_ _07246_ _07247_ _07277_ VGND VGND VPWR VPWR _07278_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_1_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09840_ net371 _05578_ VGND VGND VPWR VPWR _05589_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09771_ _04797_ _04819_ VGND VGND VPWR VPWR _04830_ sky130_fd_sc_hd__nand2_1
X_18969_ _09409_ _09423_ VGND VGND VPWR VPWR _09424_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_8_0_clock clknet_0_clock VGND VGND VPWR VPWR clknet_4_8_0_clock sky130_fd_sc_hd__clkbuf_8
X_09969_ _06051_ VGND VGND VPWR VPWR _07008_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12980_ net220 net216 _02544_ _02408_ VGND VGND VPWR VPWR _02919_ sky130_fd_sc_hd__and4_1
X_11931_ net203 _01854_ VGND VGND VPWR VPWR _01870_ sky130_fd_sc_hd__nand2_1
X_14650_ _04669_ _04672_ VGND VGND VPWR VPWR _04673_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11862_ _01793_ _01800_ VGND VGND VPWR VPWR _01801_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13601_ net248 _02546_ _03559_ _03557_ VGND VGND VPWR VPWR _03560_ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10813_ _00696_ _00698_ _00751_ VGND VGND VPWR VPWR _00752_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_156_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14581_ _03912_ _03918_ VGND VGND VPWR VPWR _04597_ sky130_fd_sc_hd__nor2_1
X_11793_ _01710_ _01728_ _01729_ _01730_ _01731_ VGND VGND VPWR VPWR _01732_ sky130_fd_sc_hd__a311o_2
XFILLER_0_39_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16320_ _06418_ _06422_ VGND VGND VPWR VPWR _06510_ sky130_fd_sc_hd__or2b_1
X_13532_ _03486_ _03490_ VGND VGND VPWR VPWR _03491_ sky130_fd_sc_hd__nor2_2
X_10744_ _00583_ _00586_ VGND VGND VPWR VPWR _00683_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_131_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16251_ _06432_ _06433_ _06290_ _01849_ VGND VGND VPWR VPWR _06434_ sky130_fd_sc_hd__a211o_2
X_13463_ _03417_ _03419_ _03421_ VGND VGND VPWR VPWR _03422_ sky130_fd_sc_hd__a21oi_1
X_10675_ _00613_ VGND VGND VPWR VPWR _00614_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15202_ _05271_ _05278_ VGND VGND VPWR VPWR _05280_ sky130_fd_sc_hd__nor2_1
X_12414_ _02347_ _02351_ _02249_ _02352_ VGND VGND VPWR VPWR _02353_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16182_ _06356_ _06357_ VGND VGND VPWR VPWR _06358_ sky130_fd_sc_hd__nor2_1
X_13394_ net262 _01907_ VGND VGND VPWR VPWR _03349_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15133_ _05194_ _05203_ VGND VGND VPWR VPWR _05205_ sky130_fd_sc_hd__or2b_1
X_12345_ net230 net226 _01835_ _01807_ VGND VGND VPWR VPWR _02284_ sky130_fd_sc_hd__and4_1
XFILLER_0_105_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15064_ net453 net162 net158 net460 VGND VGND VPWR VPWR _05129_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_120_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12276_ net208 _01875_ _02213_ _02214_ VGND VGND VPWR VPWR _02215_ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14015_ _03961_ _03962_ _03986_ VGND VGND VPWR VPWR _03987_ sky130_fd_sc_hd__a21o_1
X_11227_ _01163_ _01165_ VGND VGND VPWR VPWR _01166_ sky130_fd_sc_hd__or2b_1
X_18823_ _09249_ _09262_ VGND VGND VPWR VPWR _09264_ sky130_fd_sc_hd__xnor2_1
X_11158_ _01087_ _01095_ _01096_ VGND VGND VPWR VPWR _01097_ sky130_fd_sc_hd__o21a_1
X_10109_ net339 _05336_ _07074_ _07063_ VGND VGND VPWR VPWR _08548_ sky130_fd_sc_hd__a31o_1
X_15966_ _06028_ _06119_ _06120_ VGND VGND VPWR VPWR _06121_ sky130_fd_sc_hd__a21oi_4
X_18754_ _09181_ _09182_ VGND VGND VPWR VPWR _09188_ sky130_fd_sc_hd__and2b_1
X_11089_ net346 _00818_ _01027_ VGND VGND VPWR VPWR _01028_ sky130_fd_sc_hd__nand3_1
X_14917_ _04798_ _04959_ _04966_ VGND VGND VPWR VPWR _04967_ sky130_fd_sc_hd__or3_1
X_17705_ _08013_ _08033_ VGND VGND VPWR VPWR _08034_ sky130_fd_sc_hd__or2_1
X_15897_ _03873_ _06044_ VGND VGND VPWR VPWR _06045_ sky130_fd_sc_hd__and2_1
X_18685_ _08794_ _08620_ VGND VGND VPWR VPWR _09112_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14848_ _04889_ _04890_ VGND VGND VPWR VPWR _04891_ sky130_fd_sc_hd__or2b_1
X_17636_ _07950_ _07951_ _07923_ _07949_ VGND VGND VPWR VPWR _07958_ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17567_ _07880_ _07879_ _07801_ _07763_ VGND VGND VPWR VPWR _07882_ sky130_fd_sc_hd__o211ai_2
X_14779_ _04701_ _04814_ VGND VGND VPWR VPWR _04815_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16518_ _06715_ _06717_ VGND VGND VPWR VPWR _06728_ sky130_fd_sc_hd__xor2_1
X_19306_ clknet_4_7_0_clock _00046_ VGND VGND VPWR VPWR ki\[17\] sky130_fd_sc_hd__dfxtp_2
X_17498_ _07805_ _07502_ VGND VGND VPWR VPWR _07806_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19237_ clknet_4_13_0_clock _00119_ VGND VGND VPWR VPWR i_error\[5\] sky130_fd_sc_hd__dfxtp_1
X_16449_ _06536_ _06649_ VGND VGND VPWR VPWR _06652_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19168_ net501 net459 VGND VGND VPWR VPWR _09580_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18119_ _08475_ _08487_ _08485_ _08486_ VGND VGND VPWR VPWR _08489_ sky130_fd_sc_hd__a211o_1
X_19099_ _09536_ _06194_ _09537_ net488 VGND VGND VPWR VPWR _00105_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout404 net406 VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__buf_1
XFILLER_0_111_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout415 prev_d_error\[16\] VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__buf_2
XFILLER_0_39_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout426 net429 VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__clkbuf_4
Xfanout437 prev_d_error\[11\] VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__buf_2
X_09823_ _04764_ _05369_ VGND VGND VPWR VPWR _05402_ sky130_fd_sc_hd__and2_2
Xfanout448 net450 VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__buf_2
Xfanout459 net460 VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__clkbuf_4
X_09754_ _04621_ _04632_ VGND VGND VPWR VPWR _04643_ sky130_fd_sc_hd__or2_2
X_09685_ _03892_ VGND VGND VPWR VPWR _03903_ sky130_fd_sc_hd__buf_2
XFILLER_0_146_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_126_Right_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout11 net333 VGND VGND VPWR VPWR net566 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10460_ net352 _06623_ _00398_ VGND VGND VPWR VPWR _00399_ sky130_fd_sc_hd__and3_1
XFILLER_0_150_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10391_ _00248_ _00246_ VGND VGND VPWR VPWR _00330_ sky130_fd_sc_hd__and2b_1
XFILLER_0_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12130_ _02035_ _02044_ VGND VGND VPWR VPWR _02069_ sky130_fd_sc_hd__and2_1
X_12061_ _01936_ _01945_ _01999_ VGND VGND VPWR VPWR _02000_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_102_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11012_ _00948_ _00949_ _00950_ VGND VGND VPWR VPWR _00951_ sky130_fd_sc_hd__nand3_2
XPHY_EDGE_ROW_8_Left_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15820_ _05100_ _05957_ _05959_ VGND VGND VPWR VPWR _05960_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15751_ _05876_ _05883_ VGND VGND VPWR VPWR _05884_ sky130_fd_sc_hd__and2_1
X_12963_ net216 _02410_ _02843_ VGND VGND VPWR VPWR _02902_ sky130_fd_sc_hd__a21oi_1
X_14702_ net421 net170 _04559_ _04560_ VGND VGND VPWR VPWR _04730_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_99_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11914_ _01852_ VGND VGND VPWR VPWR _01853_ sky130_fd_sc_hd__buf_2
X_18470_ _08615_ _08622_ VGND VGND VPWR VPWR _08875_ sky130_fd_sc_hd__nor2_1
X_15682_ _05807_ _05804_ VGND VGND VPWR VPWR _05808_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12894_ _02808_ _02831_ _02832_ VGND VGND VPWR VPWR _02833_ sky130_fd_sc_hd__and3_1
X_17421_ _07719_ _07720_ VGND VGND VPWR VPWR _07721_ sky130_fd_sc_hd__or2b_1
X_14633_ _04649_ _04652_ VGND VGND VPWR VPWR _04655_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11845_ _01700_ _01753_ VGND VGND VPWR VPWR _01784_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_157_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17352_ _07643_ _07644_ VGND VGND VPWR VPWR _07645_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14564_ _04576_ _04578_ VGND VGND VPWR VPWR _04579_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11776_ _00613_ prev_error\[2\] VGND VGND VPWR VPWR _01715_ sky130_fd_sc_hd__or2b_1
XFILLER_0_138_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16303_ _06316_ _06318_ VGND VGND VPWR VPWR _06492_ sky130_fd_sc_hd__nand2_1
X_13515_ _03433_ _03473_ VGND VGND VPWR VPWR _03474_ sky130_fd_sc_hd__nor2_1
X_17283_ _07568_ VGND VGND VPWR VPWR _07570_ sky130_fd_sc_hd__buf_2
X_10727_ _00363_ _00665_ VGND VGND VPWR VPWR _00666_ sky130_fd_sc_hd__xnor2_4
X_14495_ net435 net146 _04410_ _04411_ VGND VGND VPWR VPWR _04503_ sky130_fd_sc_hd__o2bb2a_1
X_19022_ _04126_ _09446_ _09355_ _09481_ VGND VGND VPWR VPWR _09482_ sky130_fd_sc_hd__or4b_1
X_16234_ net272 _06404_ _06415_ _06412_ VGND VGND VPWR VPWR _06416_ sky130_fd_sc_hd__a31o_1
XFILLER_0_153_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13446_ _03403_ _03221_ _03404_ VGND VGND VPWR VPWR _03405_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10658_ _00579_ _00594_ _00596_ VGND VGND VPWR VPWR _00597_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16165_ net293 _06336_ _06338_ _06339_ VGND VGND VPWR VPWR _06340_ sky130_fd_sc_hd__a31o_1
XFILLER_0_24_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13377_ _03325_ _03328_ _03255_ _03306_ VGND VGND VPWR VPWR _03330_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10589_ _00432_ _00452_ VGND VGND VPWR VPWR _00528_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15116_ _05184_ _05170_ _05178_ VGND VGND VPWR VPWR _05186_ sky130_fd_sc_hd__and3_1
X_12328_ net242 net238 _01786_ _01798_ VGND VGND VPWR VPWR _02267_ sky130_fd_sc_hd__and4_1
X_16096_ _06262_ net101 _01698_ VGND VGND VPWR VPWR _06264_ sky130_fd_sc_hd__nand3b_1
X_15047_ _05109_ _05023_ VGND VGND VPWR VPWR _05110_ sky130_fd_sc_hd__xnor2_1
X_12259_ _02079_ _02197_ VGND VGND VPWR VPWR _02198_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18806_ _09229_ _09244_ VGND VGND VPWR VPWR _09245_ sky130_fd_sc_hd__xnor2_1
X_16998_ _07253_ _07255_ VGND VGND VPWR VPWR _07256_ sky130_fd_sc_hd__or2_1
X_18737_ _08818_ VGND VGND VPWR VPWR _09169_ sky130_fd_sc_hd__inv_2
X_15949_ _06061_ _06064_ VGND VGND VPWR VPWR _06102_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_149_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18668_ _06145_ _09092_ VGND VGND VPWR VPWR _09093_ sky130_fd_sc_hd__xor2_1
XFILLER_0_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17619_ _07659_ _07937_ _07938_ VGND VGND VPWR VPWR _07939_ sky130_fd_sc_hd__a21oi_1
X_18599_ _09014_ _09016_ _08964_ VGND VGND VPWR VPWR _09017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout201 kd_1\[17\] VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout212 kd_1\[14\] VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_2
Xfanout223 kd_1\[11\] VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__clkbuf_4
Xfanout234 net235 VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__buf_2
Xfanout245 kd_1\[6\] VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__buf_2
Xfanout256 net257 VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__clkbuf_4
X_09806_ net365 _04885_ net539 net368 VGND VGND VPWR VPWR _05215_ sky130_fd_sc_hd__a22oi_1
Xfanout267 net268 VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout278 ki\[15\] VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__buf_2
Xfanout289 net290 VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__buf_2
X_09737_ net74 net16 VGND VGND VPWR VPWR _04456_ sky130_fd_sc_hd__or2b_1
XFILLER_0_97_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09668_ net55 _03625_ _03658_ net310 VGND VGND VPWR VPWR _00053_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09599_ net35 net34 net37 net36 VGND VGND VPWR VPWR _03014_ sky130_fd_sc_hd__or4_1
XFILLER_0_38_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11630_ _01538_ _01548_ _01562_ VGND VGND VPWR VPWR _01569_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11561_ _01498_ _01499_ VGND VGND VPWR VPWR _01500_ sky130_fd_sc_hd__or2b_1
X_13300_ _03215_ _03252_ VGND VGND VPWR VPWR _03253_ sky130_fd_sc_hd__and2_1
X_10512_ _00434_ _00449_ _00450_ VGND VGND VPWR VPWR _00451_ sky130_fd_sc_hd__a21oi_1
X_14280_ _04264_ _04265_ net407 net165 VGND VGND VPWR VPWR _04266_ sky130_fd_sc_hd__and4bb_1
X_11492_ _01420_ _01428_ _01430_ VGND VGND VPWR VPWR _01431_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13231_ net239 _02222_ _02089_ net244 VGND VGND VPWR VPWR _03184_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10443_ net364 _05963_ _05974_ VGND VGND VPWR VPWR _00382_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13162_ net232 net228 _02330_ _02408_ VGND VGND VPWR VPWR _03112_ sky130_fd_sc_hd__and4_1
XFILLER_0_60_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10374_ _00307_ _00311_ _00300_ VGND VGND VPWR VPWR _00313_ sky130_fd_sc_hd__o21ai_1
X_12113_ _02050_ _02051_ VGND VGND VPWR VPWR _02052_ sky130_fd_sc_hd__and2_1
X_13093_ _03007_ _03009_ VGND VGND VPWR VPWR _03037_ sky130_fd_sc_hd__nand2_1
X_17970_ net322 _07181_ _07567_ net318 VGND VGND VPWR VPWR _08325_ sky130_fd_sc_hd__a22oi_1
X_16921_ _07168_ _07170_ VGND VGND VPWR VPWR _07171_ sky130_fd_sc_hd__xnor2_1
X_12044_ _01979_ _01982_ VGND VGND VPWR VPWR _01983_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16852_ _07094_ VGND VGND VPWR VPWR _07095_ sky130_fd_sc_hd__clkbuf_4
X_15803_ _05671_ _05733_ _05939_ _05940_ VGND VGND VPWR VPWR _05942_ sky130_fd_sc_hd__o22a_1
X_16783_ _07017_ _07018_ VGND VGND VPWR VPWR _07020_ sky130_fd_sc_hd__xnor2_2
X_13995_ net434 net128 VGND VGND VPWR VPWR _03967_ sky130_fd_sc_hd__nand2_1
X_15734_ _05829_ _05863_ VGND VGND VPWR VPWR _05866_ sky130_fd_sc_hd__xnor2_1
X_18522_ _08792_ _08929_ VGND VGND VPWR VPWR _08932_ sky130_fd_sc_hd__or2_1
X_12946_ _02883_ _02878_ VGND VGND VPWR VPWR _02885_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15665_ _05763_ _05789_ VGND VGND VPWR VPWR _05790_ sky130_fd_sc_hd__or2_1
X_18453_ _08590_ _08848_ _08849_ _08855_ VGND VGND VPWR VPWR _08857_ sky130_fd_sc_hd__o31a_1
X_12877_ _02814_ _02815_ VGND VGND VPWR VPWR _02816_ sky130_fd_sc_hd__nor2_1
X_14616_ _04535_ _04635_ VGND VGND VPWR VPWR _04636_ sky130_fd_sc_hd__and2_1
X_17404_ _07700_ _07702_ _07611_ _07226_ VGND VGND VPWR VPWR _07703_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_157_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11828_ _01762_ _01766_ VGND VGND VPWR VPWR _01767_ sky130_fd_sc_hd__and2_1
X_18384_ _08780_ _08743_ VGND VGND VPWR VPWR _08781_ sky130_fd_sc_hd__nor2_1
X_15596_ _05706_ _05702_ VGND VGND VPWR VPWR _05714_ sky130_fd_sc_hd__or2b_1
XFILLER_0_55_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17335_ _07625_ _07626_ VGND VGND VPWR VPWR _07627_ sky130_fd_sc_hd__nor2_1
X_14547_ net426 net169 net160 prev_d_error\[12\] VGND VGND VPWR VPWR _04560_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_44_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11759_ _09131_ _01697_ VGND VGND VPWR VPWR _01698_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_55_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17266_ net295 _06991_ VGND VGND VPWR VPWR _07551_ sky130_fd_sc_hd__nand2_2
X_14478_ net465 net125 _04482_ VGND VGND VPWR VPWR _04484_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19005_ _09463_ _09192_ VGND VGND VPWR VPWR _09464_ sky130_fd_sc_hd__xor2_1
X_16217_ _06361_ _06395_ _06396_ VGND VGND VPWR VPWR _06397_ sky130_fd_sc_hd__a21o_1
X_13429_ _03293_ _03295_ VGND VGND VPWR VPWR _03387_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17197_ net328 net514 _07472_ _07474_ VGND VGND VPWR VPWR _07475_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16148_ prev_error\[18\] _05072_ VGND VGND VPWR VPWR _06321_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16079_ _06230_ _06244_ VGND VGND VPWR VPWR _06245_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput1 iterate_enable VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_89_Left_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10090_ _08284_ _08317_ _08328_ VGND VGND VPWR VPWR _08339_ sky130_fd_sc_hd__nor3_1
XFILLER_0_11_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_98_Left_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12800_ net218 _02224_ _02332_ net216 VGND VGND VPWR VPWR _02739_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_97_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13780_ _03738_ _03744_ net108 _03745_ VGND VGND VPWR VPWR _03746_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_97_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10992_ _00926_ _00930_ VGND VGND VPWR VPWR _00931_ sky130_fd_sc_hd__or2b_1
X_12731_ _02668_ _02669_ VGND VGND VPWR VPWR _02670_ sky130_fd_sc_hd__or2b_1
X_15450_ net480 net157 _05471_ _05472_ VGND VGND VPWR VPWR _05553_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_155_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12662_ _02484_ _02598_ _02600_ VGND VGND VPWR VPWR _02601_ sky130_fd_sc_hd__o21a_1
X_14401_ _03917_ _03918_ _03913_ VGND VGND VPWR VPWR _04399_ sky130_fd_sc_hd__a21o_1
X_11613_ net381 _00815_ VGND VGND VPWR VPWR _01552_ sky130_fd_sc_hd__nand2_1
X_15381_ net468 net486 net166 net148 VGND VGND VPWR VPWR _05477_ sky130_fd_sc_hd__and4_1
X_12593_ _02529_ _02531_ VGND VGND VPWR VPWR _02532_ sky130_fd_sc_hd__xnor2_1
X_17120_ _07357_ _07363_ _07389_ VGND VGND VPWR VPWR _07390_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_37_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14332_ net434 net137 _04231_ _04232_ VGND VGND VPWR VPWR _04323_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_52_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11544_ _01464_ _01465_ VGND VGND VPWR VPWR _01483_ sky130_fd_sc_hd__xor2_1
XFILLER_0_37_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17051_ _07311_ _07313_ VGND VGND VPWR VPWR _07314_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14263_ _04238_ _04242_ _04245_ _04246_ VGND VGND VPWR VPWR _04248_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_123_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11475_ net405 _01178_ _01179_ net388 _01001_ VGND VGND VPWR VPWR _01414_ sky130_fd_sc_hd__a32o_1
X_16002_ _00959_ net569 _00957_ VGND VGND VPWR VPWR _06160_ sky130_fd_sc_hd__a21boi_2
X_13214_ _03161_ _03165_ _03048_ _03166_ VGND VGND VPWR VPWR _03167_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_61_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10426_ _00363_ _00364_ VGND VGND VPWR VPWR _00365_ sky130_fd_sc_hd__xnor2_4
X_14194_ _04132_ _04134_ _04171_ VGND VGND VPWR VPWR _04172_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_104_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13145_ net269 _01851_ VGND VGND VPWR VPWR _03094_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10357_ _00290_ _00295_ VGND VGND VPWR VPWR _00296_ sky130_fd_sc_hd__xnor2_1
X_13076_ _03010_ _03016_ VGND VGND VPWR VPWR _03018_ sky130_fd_sc_hd__nand2_1
X_17953_ _08304_ _08305_ VGND VGND VPWR VPWR _08307_ sky130_fd_sc_hd__xor2_2
X_10288_ net568 _00226_ VGND VGND VPWR VPWR _00227_ sky130_fd_sc_hd__nand2_1
X_16904_ _07048_ _07152_ VGND VGND VPWR VPWR _07153_ sky130_fd_sc_hd__or2_1
X_12027_ _01953_ _01965_ VGND VGND VPWR VPWR _01966_ sky130_fd_sc_hd__xor2_1
X_17884_ _08180_ _08230_ VGND VGND VPWR VPWR _08231_ sky130_fd_sc_hd__nor2_1
X_16835_ _07073_ _07076_ VGND VGND VPWR VPWR _07077_ sky130_fd_sc_hd__or2_1
X_16766_ _06984_ _06987_ _07000_ VGND VGND VPWR VPWR _07001_ sky130_fd_sc_hd__a21bo_1
X_13978_ _03902_ _03907_ _03949_ VGND VGND VPWR VPWR _03950_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_87_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18505_ _08843_ _08912_ _08913_ VGND VGND VPWR VPWR _08914_ sky130_fd_sc_hd__a21oi_1
X_15717_ _05833_ _05835_ VGND VGND VPWR VPWR _05847_ sky130_fd_sc_hd__nor2_1
X_12929_ _02862_ _02840_ VGND VGND VPWR VPWR _02868_ sky130_fd_sc_hd__or2b_1
X_16697_ _06923_ _06924_ VGND VGND VPWR VPWR _06925_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18436_ _06159_ _06162_ VGND VGND VPWR VPWR _08838_ sky130_fd_sc_hd__nor2_1
X_15648_ _05709_ _05770_ VGND VGND VPWR VPWR _05771_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15579_ _05645_ _05647_ VGND VGND VPWR VPWR _05695_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18367_ _08761_ _08743_ VGND VGND VPWR VPWR _08762_ sky130_fd_sc_hd__or2_2
X_17318_ _07605_ _07606_ _07607_ VGND VGND VPWR VPWR _07608_ sky130_fd_sc_hd__nand3_1
XFILLER_0_113_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18298_ _08683_ _08684_ _08685_ VGND VGND VPWR VPWR _08686_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17249_ _07517_ _07530_ _07531_ VGND VGND VPWR VPWR _07532_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11260_ _01152_ _01166_ _01168_ VGND VGND VPWR VPWR _01199_ sky130_fd_sc_hd__and3_1
X_10211_ _09546_ _09589_ VGND VGND VPWR VPWR _09595_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11191_ _01044_ _01129_ VGND VGND VPWR VPWR _01130_ sky130_fd_sc_hd__nand2_2
XFILLER_0_101_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10142_ _08889_ _08900_ VGND VGND VPWR VPWR _08911_ sky130_fd_sc_hd__xnor2_2
X_10073_ _06711_ _08141_ VGND VGND VPWR VPWR _08152_ sky130_fd_sc_hd__or2_1
X_14950_ _04927_ _04981_ _04983_ VGND VGND VPWR VPWR _05003_ sky130_fd_sc_hd__a21oi_1
X_13901_ _02983_ _03867_ VGND VGND VPWR VPWR _03868_ sky130_fd_sc_hd__nand2_1
X_14881_ _04920_ _04925_ _04912_ _04926_ VGND VGND VPWR VPWR _04927_ sky130_fd_sc_hd__o211ai_2
X_13832_ _03611_ _03065_ _03612_ VGND VGND VPWR VPWR _03798_ sky130_fd_sc_hd__or3_2
X_16620_ net303 _06335_ VGND VGND VPWR VPWR _06840_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16551_ _06365_ _06757_ VGND VGND VPWR VPWR _06764_ sky130_fd_sc_hd__xnor2_1
X_13763_ _03611_ _03503_ _02745_ VGND VGND VPWR VPWR _03729_ sky130_fd_sc_hd__or3b_1
X_10975_ _00910_ _00912_ _00913_ VGND VGND VPWR VPWR _00914_ sky130_fd_sc_hd__a21o_1
X_12714_ _02651_ _02652_ VGND VGND VPWR VPWR _02653_ sky130_fd_sc_hd__xnor2_1
X_15502_ _05537_ _05609_ VGND VGND VPWR VPWR _05610_ sky130_fd_sc_hd__nor2_1
X_16482_ _06598_ _06687_ VGND VGND VPWR VPWR _06688_ sky130_fd_sc_hd__xnor2_1
X_19270_ clknet_4_6_0_clock _00057_ VGND VGND VPWR VPWR kp\[0\] sky130_fd_sc_hd__dfxtp_1
X_13694_ _03656_ _03657_ _03659_ VGND VGND VPWR VPWR _03660_ sky130_fd_sc_hd__nand3_1
XFILLER_0_128_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15433_ _05447_ _05527_ _05505_ _05526_ VGND VGND VPWR VPWR _05535_ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18221_ i_error\[13\] _08535_ VGND VGND VPWR VPWR _08601_ sky130_fd_sc_hd__xnor2_2
X_12645_ net250 _01798_ VGND VGND VPWR VPWR _02584_ sky130_fd_sc_hd__nand2_2
XFILLER_0_150_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15364_ _05385_ _05456_ VGND VGND VPWR VPWR _05459_ sky130_fd_sc_hd__nand2_1
X_18152_ _06750_ _08524_ VGND VGND VPWR VPWR _08525_ sky130_fd_sc_hd__xor2_2
X_12576_ _02513_ _02514_ VGND VGND VPWR VPWR _02515_ sky130_fd_sc_hd__xnor2_1
X_17103_ _07232_ _07233_ _07069_ _07193_ VGND VGND VPWR VPWR _07372_ sky130_fd_sc_hd__a2bb2o_1
X_14315_ _04227_ _04228_ VGND VGND VPWR VPWR _04305_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11527_ _01462_ _01463_ VGND VGND VPWR VPWR _01466_ sky130_fd_sc_hd__nor2_1
X_18083_ _08443_ _08445_ _08448_ VGND VGND VPWR VPWR _08450_ sky130_fd_sc_hd__a21bo_2
X_15295_ _05379_ _05382_ VGND VGND VPWR VPWR _05383_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17034_ _07290_ _07295_ VGND VGND VPWR VPWR _07296_ sky130_fd_sc_hd__xnor2_2
X_14246_ _03955_ _04227_ _04228_ _03915_ VGND VGND VPWR VPWR _04229_ sky130_fd_sc_hd__a31o_1
XFILLER_0_151_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11458_ _01391_ _01396_ VGND VGND VPWR VPWR _01397_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10409_ _00346_ _00347_ VGND VGND VPWR VPWR _00348_ sky130_fd_sc_hd__nand2_1
X_14177_ _04092_ _04102_ _04151_ _04152_ VGND VGND VPWR VPWR _04153_ sky130_fd_sc_hd__o211ai_4
X_11389_ _01260_ _01318_ _01322_ VGND VGND VPWR VPWR _01328_ sky130_fd_sc_hd__a21o_1
X_13128_ _03073_ _03074_ VGND VGND VPWR VPWR _03075_ sky130_fd_sc_hd__and2_1
X_18985_ _09440_ _09075_ _09441_ VGND VGND VPWR VPWR _09442_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13059_ _02998_ _02948_ VGND VGND VPWR VPWR _02999_ sky130_fd_sc_hd__nor2_1
X_17936_ net307 _02932_ VGND VGND VPWR VPWR _08288_ sky130_fd_sc_hd__nand2_1
X_17867_ _08210_ _08211_ VGND VGND VPWR VPWR _08212_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16818_ net303 _06409_ VGND VGND VPWR VPWR _07058_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17798_ _07996_ _08010_ VGND VGND VPWR VPWR _08136_ sky130_fd_sc_hd__xor2_2
X_16749_ net288 _06468_ _06621_ net285 VGND VGND VPWR VPWR _06982_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_48_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18419_ net516 _08568_ VGND VGND VPWR VPWR _08819_ sky130_fd_sc_hd__xor2_2
XFILLER_0_118_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput70 target[1] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_6
XFILLER_0_3_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09985_ net336 _07008_ _07162_ VGND VGND VPWR VPWR _07184_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10760_ _00696_ _00698_ VGND VGND VPWR VPWR _00699_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_149_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_4_0_clock clknet_0_clock VGND VGND VPWR VPWR clknet_4_4_0_clock sky130_fd_sc_hd__clkbuf_8
XFILLER_0_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10691_ _00532_ _00544_ VGND VGND VPWR VPWR _00630_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_109_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12430_ _02367_ _02368_ VGND VGND VPWR VPWR _02369_ sky130_fd_sc_hd__xor2_2
XFILLER_0_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12361_ _02283_ _02298_ VGND VGND VPWR VPWR _02300_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14100_ net428 net124 net121 net433 VGND VGND VPWR VPWR _04072_ sky130_fd_sc_hd__a22oi_2
X_11312_ _01185_ _01184_ _01174_ VGND VGND VPWR VPWR _01251_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15080_ _05040_ _05145_ VGND VGND VPWR VPWR _05146_ sky130_fd_sc_hd__nor2_1
X_12292_ _02215_ _02216_ _02230_ VGND VGND VPWR VPWR _02231_ sky130_fd_sc_hd__a21bo_1
X_14031_ _03998_ _04000_ _04002_ VGND VGND VPWR VPWR _04003_ sky130_fd_sc_hd__o21ai_2
X_11243_ _01049_ _01180_ VGND VGND VPWR VPWR _01182_ sky130_fd_sc_hd__and2_1
XFILLER_0_132_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11174_ _01031_ _01112_ VGND VGND VPWR VPWR _01113_ sky130_fd_sc_hd__and2_1
X_10125_ _08097_ _05336_ _08713_ VGND VGND VPWR VPWR _08724_ sky130_fd_sc_hd__or3b_1
X_18770_ _08998_ _09007_ _09204_ VGND VGND VPWR VPWR _09205_ sky130_fd_sc_hd__o21ai_1
X_15982_ _01685_ _06137_ VGND VGND VPWR VPWR _06138_ sky130_fd_sc_hd__xor2_4
X_17721_ _08044_ _08045_ _08038_ VGND VGND VPWR VPWR _08051_ sky130_fd_sc_hd__o21ai_2
X_10056_ _07789_ _05644_ VGND VGND VPWR VPWR _07965_ sky130_fd_sc_hd__and2b_1
X_14933_ _04927_ _04981_ _04983_ VGND VGND VPWR VPWR _04985_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17652_ _07971_ _07970_ _07969_ VGND VGND VPWR VPWR _07975_ sky130_fd_sc_hd__a21boi_1
X_14864_ _04906_ _04908_ VGND VGND VPWR VPWR _04909_ sky130_fd_sc_hd__or2b_1
XFILLER_0_98_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16603_ _06797_ _06818_ _06820_ VGND VGND VPWR VPWR _06822_ sky130_fd_sc_hd__o21a_1
XFILLER_0_86_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13815_ _03744_ _03779_ _03772_ _03777_ VGND VGND VPWR VPWR _03781_ sky130_fd_sc_hd__a211oi_1
X_14795_ _04829_ _04832_ VGND VGND VPWR VPWR _04833_ sky130_fd_sc_hd__nor2_1
X_17583_ _07896_ _07898_ VGND VGND VPWR VPWR _07900_ sky130_fd_sc_hd__nor2_1
X_19322_ clknet_4_0_0_clock _00005_ VGND VGND VPWR VPWR kd_1\[14\] sky130_fd_sc_hd__dfxtp_1
X_13746_ _03705_ _03711_ VGND VGND VPWR VPWR _03712_ sky130_fd_sc_hd__or2b_1
X_16534_ _06742_ _06745_ VGND VGND VPWR VPWR _06746_ sky130_fd_sc_hd__and2b_1
X_10958_ _00884_ _00896_ VGND VGND VPWR VPWR _00897_ sky130_fd_sc_hd__nor2_2
XFILLER_0_57_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19253_ clknet_4_11_0_clock _00135_ VGND VGND VPWR VPWR prev_d_error\[2\] sky130_fd_sc_hd__dfxtp_1
X_13677_ net263 _02330_ _03640_ VGND VGND VPWR VPWR _03641_ sky130_fd_sc_hd__and3_1
X_16465_ _06668_ _06669_ VGND VGND VPWR VPWR _06670_ sky130_fd_sc_hd__or2_1
X_10889_ _00796_ _00827_ VGND VGND VPWR VPWR _00828_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_156_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18204_ i_error\[8\] _08580_ _08582_ VGND VGND VPWR VPWR _08583_ sky130_fd_sc_hd__and3_1
X_12628_ _02471_ _02562_ _02566_ VGND VGND VPWR VPWR _02567_ sky130_fd_sc_hd__o21a_1
X_15416_ _05498_ _05494_ VGND VGND VPWR VPWR _05516_ sky130_fd_sc_hd__or2b_1
XFILLER_0_66_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19184_ net498 _08987_ VGND VGND VPWR VPWR _09590_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16396_ _06372_ _06592_ _06593_ VGND VGND VPWR VPWR _06594_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_143_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18135_ _08505_ _08506_ VGND VGND VPWR VPWR _08507_ sky130_fd_sc_hd__nor2_1
X_15347_ _05439_ VGND VGND VPWR VPWR _05440_ sky130_fd_sc_hd__inv_2
X_12559_ _02491_ _02494_ VGND VGND VPWR VPWR _02498_ sky130_fd_sc_hd__xor2_1
XFILLER_0_54_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15278_ _05278_ _05363_ VGND VGND VPWR VPWR _05364_ sky130_fd_sc_hd__nand2_1
X_18066_ net523 _08047_ _08046_ _08044_ VGND VGND VPWR VPWR _08431_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_123_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17017_ _07274_ _07276_ VGND VGND VPWR VPWR _07277_ sky130_fd_sc_hd__or2b_1
XFILLER_0_10_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14229_ _04208_ _04147_ _04151_ VGND VGND VPWR VPWR _04210_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_107_Right_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09770_ _04808_ VGND VGND VPWR VPWR _04819_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18968_ _09419_ _09422_ VGND VGND VPWR VPWR _09423_ sky130_fd_sc_hd__xnor2_1
X_17919_ _08226_ _08266_ _08268_ VGND VGND VPWR VPWR _08269_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_119_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18899_ _09346_ _08872_ _08882_ VGND VGND VPWR VPWR _09347_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09968_ _06810_ _06975_ _06986_ VGND VGND VPWR VPWR _06997_ sky130_fd_sc_hd__a21o_1
X_09899_ _06139_ _06227_ VGND VGND VPWR VPWR _06238_ sky130_fd_sc_hd__nor2_1
X_11930_ net205 _01860_ VGND VGND VPWR VPWR _01869_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11861_ _01793_ _01794_ net221 _01799_ VGND VGND VPWR VPWR _01800_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_24_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13600_ _03557_ _03558_ VGND VGND VPWR VPWR _03559_ sky130_fd_sc_hd__nor2_1
X_10812_ _00699_ _00719_ VGND VGND VPWR VPWR _00751_ sky130_fd_sc_hd__or2_1
X_14580_ _04595_ _04586_ VGND VGND VPWR VPWR _04596_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11792_ prev_error\[8\] _08174_ VGND VGND VPWR VPWR _01731_ sky130_fd_sc_hd__and2b_1
X_13531_ _03486_ _03488_ _03489_ VGND VGND VPWR VPWR _03490_ sky130_fd_sc_hd__nor3_1
XFILLER_0_27_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10743_ _00680_ _00681_ VGND VGND VPWR VPWR _00682_ sky130_fd_sc_hd__and2b_1
XFILLER_0_54_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16250_ prev_error\[9\] _06623_ _01871_ VGND VGND VPWR VPWR _06433_ sky130_fd_sc_hd__o21a_1
X_13462_ _03333_ _03420_ VGND VGND VPWR VPWR _03421_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10674_ _00612_ VGND VGND VPWR VPWR _00613_ sky130_fd_sc_hd__buf_2
XFILLER_0_125_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15201_ _05271_ _05278_ VGND VGND VPWR VPWR _05279_ sky130_fd_sc_hd__and2_1
X_12413_ _02246_ _02247_ _02237_ _02240_ VGND VGND VPWR VPWR _02352_ sky130_fd_sc_hd__a211o_1
XFILLER_0_51_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16181_ net283 _06346_ _06355_ VGND VGND VPWR VPWR _06357_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13393_ _03310_ _03346_ VGND VGND VPWR VPWR _03348_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15132_ _05181_ _05186_ _05192_ VGND VGND VPWR VPWR _05203_ sky130_fd_sc_hd__or3b_1
X_12344_ _02280_ _02282_ VGND VGND VPWR VPWR _02283_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15063_ _05124_ _05126_ VGND VGND VPWR VPWR _05128_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12275_ net217 net213 _01854_ _01861_ VGND VGND VPWR VPWR _02214_ sky130_fd_sc_hd__and4_1
X_14014_ _03983_ _03984_ _03985_ VGND VGND VPWR VPWR _03986_ sky130_fd_sc_hd__nor3_1
X_11226_ _01152_ _01164_ VGND VGND VPWR VPWR _01165_ sky130_fd_sc_hd__and2_2
X_18822_ _09260_ _09261_ VGND VGND VPWR VPWR _09262_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11157_ _01089_ _01094_ VGND VGND VPWR VPWR _01096_ sky130_fd_sc_hd__or2b_1
X_10108_ _05666_ _07492_ _08526_ VGND VGND VPWR VPWR _08537_ sky130_fd_sc_hd__o21ai_1
X_18753_ _09182_ _09181_ VGND VGND VPWR VPWR _09187_ sky130_fd_sc_hd__or2b_1
X_15965_ _06021_ _06022_ VGND VGND VPWR VPWR _06120_ sky130_fd_sc_hd__xnor2_2
X_11088_ _01025_ _01026_ VGND VGND VPWR VPWR _01027_ sky130_fd_sc_hd__and2_1
X_17704_ _08013_ _08014_ _08032_ VGND VGND VPWR VPWR _08033_ sky130_fd_sc_hd__nor3_2
X_10039_ _07316_ _07371_ _07349_ VGND VGND VPWR VPWR _07778_ sky130_fd_sc_hd__o21ai_4
X_14916_ _04960_ _04965_ VGND VGND VPWR VPWR _04966_ sky130_fd_sc_hd__nor2_1
X_18684_ _06092_ _09110_ VGND VGND VPWR VPWR _09111_ sky130_fd_sc_hd__nand2_1
X_15896_ _03872_ _02983_ _03869_ VGND VGND VPWR VPWR _06044_ sky130_fd_sc_hd__nand3_1
X_17635_ _07955_ _07956_ VGND VGND VPWR VPWR _07957_ sky130_fd_sc_hd__xnor2_1
X_14847_ _04858_ _04880_ _04856_ VGND VGND VPWR VPWR _04890_ sky130_fd_sc_hd__o21ai_1
X_17566_ _07763_ _07801_ _07879_ _07880_ VGND VGND VPWR VPWR _07881_ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14778_ _04704_ _04703_ VGND VGND VPWR VPWR _04814_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19305_ clknet_4_8_0_clock _00045_ VGND VGND VPWR VPWR ki\[16\] sky130_fd_sc_hd__dfxtp_1
X_16517_ net272 _06724_ _06725_ _06726_ VGND VGND VPWR VPWR _06727_ sky130_fd_sc_hd__a31o_1
X_13729_ _03691_ _03694_ VGND VGND VPWR VPWR _03695_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17497_ net302 _06890_ VGND VGND VPWR VPWR _07805_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19236_ clknet_4_9_0_clock _00118_ VGND VGND VPWR VPWR i_error\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16448_ _06649_ _06650_ _06548_ VGND VGND VPWR VPWR _06651_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_26_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19167_ _09559_ _09158_ _09579_ net490 VGND VGND VPWR VPWR _00138_ sky130_fd_sc_hd__o211a_1
X_16379_ _06549_ _06573_ _06558_ VGND VGND VPWR VPWR _06575_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18118_ _08485_ _08486_ _08475_ _08487_ VGND VGND VPWR VPWR _08488_ sky130_fd_sc_hd__o211a_1
X_19098_ net499 prev_error\[10\] VGND VGND VPWR VPWR _09537_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18049_ _08299_ _08409_ _08407_ _08408_ VGND VGND VPWR VPWR _08412_ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout405 net406 VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__clkbuf_4
Xfanout416 prev_d_error\[15\] VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__buf_2
X_09822_ net353 _05182_ _05380_ VGND VGND VPWR VPWR _05391_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout427 net428 VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__buf_2
Xfanout438 net440 VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__buf_2
Xfanout449 net450 VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__clkbuf_4
X_09753_ net77 net19 VGND VGND VPWR VPWR _04632_ sky130_fd_sc_hd__and2b_1
XFILLER_0_146_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09684_ net79 _03859_ net487 VGND VGND VPWR VPWR _03892_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_61_Left_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout12 net431 VGND VGND VPWR VPWR net567 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_70_Left_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10390_ net339 _00245_ VGND VGND VPWR VPWR _00329_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12060_ _01929_ _01998_ VGND VGND VPWR VPWR _01999_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11011_ _00946_ _00947_ _00941_ _00945_ VGND VGND VPWR VPWR _00950_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_99_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15750_ _05881_ _05880_ VGND VGND VPWR VPWR _05883_ sky130_fd_sc_hd__xnor2_1
X_12962_ _02895_ _02900_ VGND VGND VPWR VPWR _02901_ sky130_fd_sc_hd__xor2_1
X_14701_ _04727_ _04725_ VGND VGND VPWR VPWR _04729_ sky130_fd_sc_hd__xnor2_1
X_11913_ _01851_ VGND VGND VPWR VPWR _01852_ sky130_fd_sc_hd__buf_2
XFILLER_0_99_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15681_ _05740_ _05800_ VGND VGND VPWR VPWR _05807_ sky130_fd_sc_hd__nor2_1
X_12893_ _02709_ _02807_ _02793_ _02806_ VGND VGND VPWR VPWR _02832_ sky130_fd_sc_hd__o211ai_2
X_17420_ _07201_ _07640_ _07642_ _07639_ VGND VGND VPWR VPWR _07720_ sky130_fd_sc_hd__o22ai_1
X_14632_ _04649_ _04652_ VGND VGND VPWR VPWR _04653_ sky130_fd_sc_hd__nor2_1
X_11844_ _01775_ _01782_ VGND VGND VPWR VPWR _01783_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14563_ _04575_ _04564_ _04573_ VGND VGND VPWR VPWR _04578_ sky130_fd_sc_hd__and3_1
X_17351_ _07550_ _07581_ _07584_ VGND VGND VPWR VPWR _07644_ sky130_fd_sc_hd__o21ba_1
X_11775_ prev_error\[3\] VGND VGND VPWR VPWR _01714_ sky130_fd_sc_hd__inv_2
X_16302_ _06328_ _06489_ VGND VGND VPWR VPWR _06490_ sky130_fd_sc_hd__nand2_1
X_13514_ net249 _02332_ _03432_ VGND VGND VPWR VPWR _03473_ sky130_fd_sc_hd__a21oi_1
X_10726_ net401 _04973_ VGND VGND VPWR VPWR _00665_ sky130_fd_sc_hd__nand2_1
X_14494_ _04498_ _04501_ VGND VGND VPWR VPWR _04502_ sky130_fd_sc_hd__or2b_1
X_17282_ _07567_ VGND VGND VPWR VPWR _07568_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_109_Left_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19021_ _09209_ _09213_ _09480_ VGND VGND VPWR VPWR _09481_ sky130_fd_sc_hd__and3_1
X_13445_ kd_1\[13\] _02935_ _02915_ net220 VGND VGND VPWR VPWR _03404_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16233_ _06412_ _06413_ VGND VGND VPWR VPWR _06415_ sky130_fd_sc_hd__and2b_1
XFILLER_0_126_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10657_ _00525_ _00595_ VGND VGND VPWR VPWR _00596_ sky130_fd_sc_hd__or2_1
XFILLER_0_141_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13376_ _03255_ _03306_ _03325_ _03328_ VGND VGND VPWR VPWR _03329_ sky130_fd_sc_hd__a211o_1
XFILLER_0_106_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16164_ net300 net297 _06310_ _06320_ VGND VGND VPWR VPWR _06339_ sky130_fd_sc_hd__and4_1
X_10588_ _00500_ _00526_ VGND VGND VPWR VPWR _00527_ sky130_fd_sc_hd__xor2_4
XFILLER_0_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12327_ net242 _01786_ _02265_ VGND VGND VPWR VPWR _02266_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_51_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15115_ _05170_ _05178_ _05184_ VGND VGND VPWR VPWR _05185_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16095_ _06225_ _06228_ VGND VGND VPWR VPWR _06263_ sky130_fd_sc_hd__xnor2_1
X_15046_ _05024_ _05022_ VGND VGND VPWR VPWR _05109_ sky130_fd_sc_hd__nor2_1
X_12258_ net208 _01854_ _02078_ VGND VGND VPWR VPWR _02197_ sky130_fd_sc_hd__a21oi_1
X_11209_ _01145_ _01065_ _01147_ VGND VGND VPWR VPWR _01148_ sky130_fd_sc_hd__a21oi_1
X_12189_ net204 _01817_ VGND VGND VPWR VPWR _02128_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_118_Left_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18805_ _09242_ _09243_ VGND VGND VPWR VPWR _09244_ sky130_fd_sc_hd__nor2_1
X_16997_ _07174_ _07252_ VGND VGND VPWR VPWR _07255_ sky130_fd_sc_hd__and2_1
X_18736_ _06101_ _09167_ VGND VGND VPWR VPWR _09168_ sky130_fd_sc_hd__and2_1
X_15948_ _06075_ _06099_ _06100_ VGND VGND VPWR VPWR _06101_ sky130_fd_sc_hd__a21o_1
X_18667_ _09089_ _09091_ VGND VGND VPWR VPWR _09092_ sky130_fd_sc_hd__xor2_1
X_15879_ _04480_ _05990_ _05993_ VGND VGND VPWR VPWR _06025_ sky130_fd_sc_hd__nor3_1
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17618_ net290 net287 _02932_ net540 VGND VGND VPWR VPWR _07938_ sky130_fd_sc_hd__and4_1
XFILLER_0_25_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18598_ _08764_ _09015_ _08882_ VGND VGND VPWR VPWR _09016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17549_ _07861_ VGND VGND VPWR VPWR _07862_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_127_Left_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19219_ clknet_4_5_0_clock _00101_ VGND VGND VPWR VPWR prev_error\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_136_Left_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout202 kd_1\[17\] VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__buf_2
Xfanout213 net215 VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__buf_2
XFILLER_0_10_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout224 net225 VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__clkbuf_4
Xfanout235 kd_1\[8\] VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__clkbuf_2
Xfanout246 net247 VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__clkbuf_4
X_09805_ net369 net364 _04885_ net539 VGND VGND VPWR VPWR _05204_ sky130_fd_sc_hd__and4_1
Xfanout257 kd_1\[3\] VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__clkbuf_2
Xfanout268 net269 VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__clkbuf_4
Xfanout279 net280 VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__buf_2
XFILLER_0_157_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09736_ net15 net73 VGND VGND VPWR VPWR _04445_ sky130_fd_sc_hd__and2b_1
X_09667_ net54 _03625_ _03658_ net313 VGND VGND VPWR VPWR _00052_ sky130_fd_sc_hd__a22o_1
X_09598_ net39 net38 net23 net22 VGND VGND VPWR VPWR _03003_ sky130_fd_sc_hd__or4_1
XFILLER_0_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11560_ _01443_ _01444_ VGND VGND VPWR VPWR _01499_ sky130_fd_sc_hd__xor2_1
XFILLER_0_37_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10511_ _00436_ _00448_ VGND VGND VPWR VPWR _00450_ sky130_fd_sc_hd__and2_1
XFILLER_0_108_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11491_ _01391_ _01429_ VGND VGND VPWR VPWR _01430_ sky130_fd_sc_hd__or2_1
X_13230_ net239 _02090_ _03182_ VGND VGND VPWR VPWR _03183_ sky130_fd_sc_hd__nand3_1
XFILLER_0_134_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10442_ _00291_ _00380_ VGND VGND VPWR VPWR _00381_ sky130_fd_sc_hd__xor2_1
XFILLER_0_150_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13161_ net232 _02331_ _02408_ net229 VGND VGND VPWR VPWR _03111_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10373_ _00300_ _00307_ _00311_ VGND VGND VPWR VPWR _00312_ sky130_fd_sc_hd__or3_1
X_12112_ _02046_ _02047_ _02049_ VGND VGND VPWR VPWR _02051_ sky130_fd_sc_hd__nand3_1
X_13092_ _03026_ _03030_ _03034_ VGND VGND VPWR VPWR _03035_ sky130_fd_sc_hd__a21oi_1
X_16920_ _07169_ _07100_ VGND VGND VPWR VPWR _07170_ sky130_fd_sc_hd__xnor2_1
X_12043_ _01972_ _01981_ VGND VGND VPWR VPWR _01982_ sky130_fd_sc_hd__and2_1
X_16851_ _07093_ VGND VGND VPWR VPWR _07094_ sky130_fd_sc_hd__clkbuf_4
X_15802_ _05669_ _05671_ VGND VGND VPWR VPWR _05940_ sky130_fd_sc_hd__and2_1
X_16782_ net320 _06314_ _06318_ VGND VGND VPWR VPWR _07018_ sky130_fd_sc_hd__and3_1
X_13994_ _03963_ _03965_ VGND VGND VPWR VPWR _03966_ sky130_fd_sc_hd__nor2_1
X_18521_ _08792_ _08929_ _08930_ _08796_ VGND VGND VPWR VPWR _08931_ sky130_fd_sc_hd__a22o_1
X_15733_ _05829_ _05863_ VGND VGND VPWR VPWR _05865_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12945_ _02878_ _02883_ VGND VGND VPWR VPWR _02884_ sky130_fd_sc_hd__or2b_1
XFILLER_0_88_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18452_ i_error\[10\] _08589_ VGND VGND VPWR VPWR _08855_ sky130_fd_sc_hd__nand2_1
X_15664_ net455 net195 net191 net457 VGND VGND VPWR VPWR _05789_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_157_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12876_ _02810_ _02811_ _02813_ VGND VGND VPWR VPWR _02815_ sky130_fd_sc_hd__nor3_1
XFILLER_0_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17403_ net566 _06409_ VGND VGND VPWR VPWR _07702_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14615_ _04516_ _04534_ _04524_ _04532_ VGND VGND VPWR VPWR _04635_ sky130_fd_sc_hd__a211o_1
XFILLER_0_56_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11827_ _01763_ _01765_ VGND VGND VPWR VPWR _01766_ sky130_fd_sc_hd__or2_1
X_18383_ _08777_ _08778_ VGND VGND VPWR VPWR _08780_ sky130_fd_sc_hd__or2b_1
X_15595_ _05698_ _05701_ VGND VGND VPWR VPWR _05713_ sky130_fd_sc_hd__or2b_1
XFILLER_0_68_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17334_ _07620_ _07623_ VGND VGND VPWR VPWR _07626_ sky130_fd_sc_hd__and2_1
X_11758_ _00186_ _01696_ _00184_ VGND VGND VPWR VPWR _01697_ sky130_fd_sc_hd__a21bo_1
X_14546_ net429 net160 _04558_ VGND VGND VPWR VPWR _04559_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10709_ _00630_ _00646_ VGND VGND VPWR VPWR _00648_ sky130_fd_sc_hd__or2b_1
XFILLER_0_153_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17265_ net298 _06889_ VGND VGND VPWR VPWR _07550_ sky130_fd_sc_hd__nand2_2
X_14477_ net465 net125 _04482_ VGND VGND VPWR VPWR _04483_ sky130_fd_sc_hd__and3_1
X_11689_ _01595_ _01627_ VGND VGND VPWR VPWR _01628_ sky130_fd_sc_hd__xnor2_1
X_19004_ _09193_ _09086_ VGND VGND VPWR VPWR _09463_ sky130_fd_sc_hd__or2b_1
X_16216_ _06372_ _06375_ _06394_ VGND VGND VPWR VPWR _06396_ sky130_fd_sc_hd__o21a_1
X_13428_ _03368_ _03384_ _03323_ _03385_ VGND VGND VPWR VPWR _03386_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_102_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17196_ net319 _06400_ _07473_ VGND VGND VPWR VPWR _07474_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13359_ _03311_ _03239_ VGND VGND VPWR VPWR _03312_ sky130_fd_sc_hd__xnor2_1
X_16147_ _06319_ VGND VGND VPWR VPWR _06320_ sky130_fd_sc_hd__buf_2
XFILLER_0_140_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16078_ _06231_ _06243_ VGND VGND VPWR VPWR _06244_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15029_ _05064_ _05087_ _05088_ _05089_ VGND VGND VPWR VPWR _05090_ sky130_fd_sc_hd__nand4_2
Xinput2 measurement[0] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_1
XFILLER_0_36_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18719_ _09084_ _09137_ _09147_ VGND VGND VPWR VPWR _09149_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_144_Left_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09719_ net12 net70 VGND VGND VPWR VPWR _04258_ sky130_fd_sc_hd__nor2b_1
XPHY_EDGE_ROW_153_Left_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10991_ net401 _05413_ _00928_ _00929_ VGND VGND VPWR VPWR _00930_ sky130_fd_sc_hd__a31o_1
X_12730_ _02630_ _02631_ _02662_ VGND VGND VPWR VPWR _02669_ sky130_fd_sc_hd__a21o_1
XFILLER_0_139_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12661_ net241 _01835_ _01806_ net245 VGND VGND VPWR VPWR _02600_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14400_ _04396_ _04397_ VGND VGND VPWR VPWR _04398_ sky130_fd_sc_hd__and2_1
X_11612_ _01358_ _01549_ _01550_ _01356_ VGND VGND VPWR VPWR _01551_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12592_ _02421_ _02530_ VGND VGND VPWR VPWR _02531_ sky130_fd_sc_hd__nor2_1
X_15380_ _05471_ _05473_ _05475_ VGND VGND VPWR VPWR _05476_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14331_ _04319_ _04321_ VGND VGND VPWR VPWR _04322_ sky130_fd_sc_hd__nor2_1
X_11543_ _01415_ _01438_ _01439_ _01437_ VGND VGND VPWR VPWR _01482_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14262_ _04223_ _04227_ _04244_ VGND VGND VPWR VPWR _04246_ sky130_fd_sc_hd__nand3_1
X_17050_ _07231_ _07312_ VGND VGND VPWR VPWR _07313_ sky130_fd_sc_hd__or2_1
X_11474_ _06590_ _06601_ _01412_ _00871_ VGND VGND VPWR VPWR _01413_ sky130_fd_sc_hd__a211o_1
XFILLER_0_80_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13213_ _03023_ _03046_ _03045_ VGND VGND VPWR VPWR _03166_ sky130_fd_sc_hd__a21o_1
X_16001_ _06136_ _06138_ _06141_ _06158_ VGND VGND VPWR VPWR _06159_ sky130_fd_sc_hd__or4b_4
X_10425_ net387 _04984_ VGND VGND VPWR VPWR _00364_ sky130_fd_sc_hd__nand2_2
X_14193_ _04167_ _04169_ VGND VGND VPWR VPWR _04171_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13144_ net252 _01852_ _01813_ net267 VGND VGND VPWR VPWR _03093_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_21_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10356_ _00291_ _00292_ _00294_ VGND VGND VPWR VPWR _00295_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_131_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13075_ _03010_ _03016_ VGND VGND VPWR VPWR _03017_ sky130_fd_sc_hd__or2_1
X_17952_ _08256_ _08263_ VGND VGND VPWR VPWR _08305_ sky130_fd_sc_hd__and2b_1
X_10287_ _09558_ _09565_ VGND VGND VPWR VPWR _00226_ sky130_fd_sc_hd__nand2_2
X_16903_ _07114_ _07149_ _07150_ VGND VGND VPWR VPWR _07152_ sky130_fd_sc_hd__o21a_1
X_12026_ _01962_ _01964_ VGND VGND VPWR VPWR _01965_ sky130_fd_sc_hd__xnor2_1
X_17883_ net326 _06890_ _08179_ VGND VGND VPWR VPWR _08230_ sky130_fd_sc_hd__a21oi_1
X_16834_ _07075_ _06983_ VGND VGND VPWR VPWR _07076_ sky130_fd_sc_hd__xor2_1
XFILLER_0_88_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16765_ _06988_ _06999_ VGND VGND VPWR VPWR _07000_ sky130_fd_sc_hd__or2b_1
XFILLER_0_87_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13977_ _03943_ _03948_ VGND VGND VPWR VPWR _03949_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18504_ _08909_ _08833_ _08843_ _08912_ VGND VGND VPWR VPWR _08913_ sky130_fd_sc_hd__o22ai_1
X_15716_ _05838_ _05843_ _05845_ VGND VGND VPWR VPWR _05846_ sky130_fd_sc_hd__o21ai_1
X_12928_ _02775_ _02866_ VGND VGND VPWR VPWR _02867_ sky130_fd_sc_hd__xnor2_1
X_16696_ _06905_ _06922_ VGND VGND VPWR VPWR _06924_ sky130_fd_sc_hd__and2_1
X_18435_ _08836_ _08743_ VGND VGND VPWR VPWR _08837_ sky130_fd_sc_hd__nor2_1
X_15647_ _05697_ _05708_ _05707_ VGND VGND VPWR VPWR _05770_ sky130_fd_sc_hd__a21o_1
X_12859_ _02795_ _02797_ VGND VGND VPWR VPWR _02798_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18366_ _06169_ _08760_ VGND VGND VPWR VPWR _08761_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15578_ _05691_ _05693_ VGND VGND VPWR VPWR _05694_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17317_ net329 _06334_ _07300_ _07299_ VGND VGND VPWR VPWR _07607_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14529_ net413 net417 net175 net170 VGND VGND VPWR VPWR _04540_ sky130_fd_sc_hd__and4_1
XFILLER_0_56_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18297_ i_error\[17\] _08681_ VGND VGND VPWR VPWR _08685_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17248_ _07523_ _07524_ _07528_ _07529_ VGND VGND VPWR VPWR _07531_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17179_ _07430_ _07441_ VGND VGND VPWR VPWR _07455_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10210_ net341 _08207_ _06634_ net345 VGND VGND VPWR VPWR _09589_ sky130_fd_sc_hd__a22oi_1
X_11190_ _01125_ _01128_ VGND VGND VPWR VPWR _01129_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10141_ net349 _05677_ VGND VGND VPWR VPWR _08900_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_0_0_clock clknet_0_clock VGND VGND VPWR VPWR clknet_4_0_0_clock sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10072_ _06568_ _06689_ _06700_ VGND VGND VPWR VPWR _08141_ sky130_fd_sc_hd__nor3_1
XFILLER_0_27_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13900_ _02875_ _02982_ VGND VGND VPWR VPWR _03867_ sky130_fd_sc_hd__or2_1
X_14880_ _04902_ _04909_ _04911_ VGND VGND VPWR VPWR _04926_ sky130_fd_sc_hd__nand3_1
XFILLER_0_89_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13831_ net251 _02934_ _02546_ net268 VGND VGND VPWR VPWR _03797_ sky130_fd_sc_hd__a22o_1
X_16550_ net306 _06311_ _06759_ _06762_ VGND VGND VPWR VPWR _06763_ sky130_fd_sc_hd__a31oi_2
X_13762_ net267 _02330_ _02745_ net251 VGND VGND VPWR VPWR _03728_ sky130_fd_sc_hd__a22o_1
X_10974_ _00902_ _00906_ _00909_ VGND VGND VPWR VPWR _00913_ sky130_fd_sc_hd__nor3_1
XFILLER_0_57_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15501_ _05533_ _05536_ VGND VGND VPWR VPWR _05609_ sky130_fd_sc_hd__and2_1
X_12713_ _02549_ _02548_ VGND VGND VPWR VPWR _02652_ sky130_fd_sc_hd__or2b_1
X_16481_ net296 _06352_ VGND VGND VPWR VPWR _06687_ sky130_fd_sc_hd__nand2_1
X_13693_ _03594_ _03655_ _03650_ _03654_ VGND VGND VPWR VPWR _03659_ sky130_fd_sc_hd__a211o_1
X_18220_ _08587_ _08590_ _08597_ _08598_ _08599_ VGND VGND VPWR VPWR _08600_ sky130_fd_sc_hd__o311a_2
X_15432_ _05532_ VGND VGND VPWR VPWR _05533_ sky130_fd_sc_hd__inv_2
X_12644_ _02580_ _02582_ VGND VGND VPWR VPWR _02583_ sky130_fd_sc_hd__or2b_1
XFILLER_0_150_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18151_ _06836_ _08522_ _08523_ VGND VGND VPWR VPWR _08524_ sky130_fd_sc_hd__a21o_1
X_12575_ _02400_ _02399_ VGND VGND VPWR VPWR _02514_ sky130_fd_sc_hd__and2b_1
X_15363_ _05385_ _05456_ VGND VGND VPWR VPWR _05458_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17102_ _07071_ _07369_ VGND VGND VPWR VPWR _07370_ sky130_fd_sc_hd__or2_1
X_14314_ _04297_ _04303_ VGND VGND VPWR VPWR _04304_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11526_ net381 _00516_ VGND VGND VPWR VPWR _01465_ sky130_fd_sc_hd__nand2_1
X_18082_ _08446_ _08447_ VGND VGND VPWR VPWR _08448_ sky130_fd_sc_hd__or2b_1
XFILLER_0_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15294_ _04016_ net197 _05378_ VGND VGND VPWR VPWR _05382_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17033_ _06364_ _06353_ _07293_ VGND VGND VPWR VPWR _07295_ sky130_fd_sc_hd__a21oi_1
X_14245_ _04218_ _04221_ _04226_ VGND VGND VPWR VPWR _04228_ sky130_fd_sc_hd__or3_1
X_11457_ _01393_ _01395_ VGND VGND VPWR VPWR _01396_ sky130_fd_sc_hd__xor2_1
XFILLER_0_21_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10408_ _00273_ _00314_ VGND VGND VPWR VPWR _00347_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14176_ _04124_ _04125_ _04150_ VGND VGND VPWR VPWR _04152_ sky130_fd_sc_hd__o21ai_2
X_11388_ _01324_ _01285_ _00244_ net382 VGND VGND VPWR VPWR _01327_ sky130_fd_sc_hd__a22oi_1
X_13127_ _02987_ _03049_ VGND VGND VPWR VPWR _03074_ sky130_fd_sc_hd__xor2_1
X_10339_ _00276_ _00277_ VGND VGND VPWR VPWR _00278_ sky130_fd_sc_hd__and2b_1
X_18984_ _08733_ _08730_ VGND VGND VPWR VPWR _09441_ sky130_fd_sc_hd__and2b_1
X_13058_ net261 _01859_ VGND VGND VPWR VPWR _02998_ sky130_fd_sc_hd__nand2_1
X_17935_ net310 _07570_ VGND VGND VPWR VPWR _08287_ sky130_fd_sc_hd__nand2_1
X_12009_ _01929_ _01947_ VGND VGND VPWR VPWR _01948_ sky130_fd_sc_hd__and2b_1
X_17866_ _08205_ _08206_ _08209_ VGND VGND VPWR VPWR _08211_ sky130_fd_sc_hd__nand3_1
X_16817_ ki\[7\] _06345_ VGND VGND VPWR VPWR _07057_ sky130_fd_sc_hd__nand2_2
XFILLER_0_89_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17797_ _08104_ _08116_ VGND VGND VPWR VPWR _08135_ sky130_fd_sc_hd__or2_1
X_16748_ net285 _06468_ _06980_ VGND VGND VPWR VPWR _06981_ sky130_fd_sc_hd__and3_1
XFILLER_0_124_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16679_ _06783_ _06787_ VGND VGND VPWR VPWR _06905_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18418_ _08817_ net571 VGND VGND VPWR VPWR _08818_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18349_ _06261_ _08618_ VGND VGND VPWR VPWR _08742_ sky130_fd_sc_hd__and2b_2
XFILLER_0_32_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput60 target[0] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_1
Xinput71 target[2] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_1
XFILLER_0_142_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09984_ net336 _07008_ _07162_ VGND VGND VPWR VPWR _07173_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10690_ _00594_ _00628_ VGND VGND VPWR VPWR _00629_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12360_ _02283_ _02298_ VGND VGND VPWR VPWR _02299_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11311_ _01185_ _01174_ _01184_ VGND VGND VPWR VPWR _01250_ sky130_fd_sc_hd__nand3_2
X_12291_ _02217_ _02228_ _02229_ VGND VGND VPWR VPWR _02230_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_133_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14030_ _03997_ _04001_ VGND VGND VPWR VPWR _04002_ sky130_fd_sc_hd__and2_1
X_11242_ _01049_ _01180_ VGND VGND VPWR VPWR _01181_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11173_ _01025_ _01028_ _01030_ VGND VGND VPWR VPWR _01112_ sky130_fd_sc_hd__nand3_1
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10124_ _08691_ _08702_ VGND VGND VPWR VPWR _08713_ sky130_fd_sc_hd__xnor2_1
X_15981_ _01134_ _01209_ _01681_ _01686_ VGND VGND VPWR VPWR _06137_ sky130_fd_sc_hd__o31a_2
X_17720_ _08038_ _08044_ _08045_ VGND VGND VPWR VPWR _08050_ sky130_fd_sc_hd__or3_1
X_10055_ _07932_ _07943_ VGND VGND VPWR VPWR _07954_ sky130_fd_sc_hd__or2_1
X_14932_ _04982_ _04980_ VGND VGND VPWR VPWR _04983_ sky130_fd_sc_hd__xnor2_1
X_17651_ _07884_ _07972_ _07973_ VGND VGND VPWR VPWR _07974_ sky130_fd_sc_hd__o21ai_1
X_14863_ _04899_ _04901_ VGND VGND VPWR VPWR _04908_ sky130_fd_sc_hd__xnor2_1
X_16602_ _06398_ _06724_ _06819_ VGND VGND VPWR VPWR _06820_ sky130_fd_sc_hd__or3_1
X_13814_ _03772_ _03777_ _03744_ _03779_ VGND VGND VPWR VPWR _03780_ sky130_fd_sc_hd__o211a_1
X_17582_ net315 _06400_ _07897_ VGND VGND VPWR VPWR _07898_ sky130_fd_sc_hd__and3_1
X_14794_ _04829_ _04831_ net439 net163 VGND VGND VPWR VPWR _04832_ sky130_fd_sc_hd__and4bb_1
X_19321_ clknet_4_1_0_clock _00004_ VGND VGND VPWR VPWR kd_1\[13\] sky130_fd_sc_hd__dfxtp_1
X_16533_ _06707_ _06743_ VGND VGND VPWR VPWR _06745_ sky130_fd_sc_hd__nand2_1
X_13745_ _03705_ _03709_ _03710_ VGND VGND VPWR VPWR _03711_ sky130_fd_sc_hd__or3_1
X_10957_ _00893_ _00895_ VGND VGND VPWR VPWR _00896_ sky130_fd_sc_hd__and2b_1
X_19252_ clknet_4_10_0_clock _00134_ VGND VGND VPWR VPWR prev_d_error\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16464_ _06589_ _06666_ VGND VGND VPWR VPWR _06669_ sky130_fd_sc_hd__and2_1
X_13676_ _03638_ _03639_ VGND VGND VPWR VPWR _03640_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10888_ _00716_ _00797_ _00823_ _00826_ VGND VGND VPWR VPWR _00827_ sky130_fd_sc_hd__a31oi_4
X_18203_ _08499_ _08540_ _08481_ VGND VGND VPWR VPWR _08582_ sky130_fd_sc_hd__o21ai_1
X_15415_ net432 net197 _05514_ VGND VGND VPWR VPWR _05515_ sky130_fd_sc_hd__nand3_1
X_12627_ _02563_ _02565_ VGND VGND VPWR VPWR _02566_ sky130_fd_sc_hd__or2b_1
X_19183_ _09550_ _09004_ _09588_ net492 VGND VGND VPWR VPWR _00146_ sky130_fd_sc_hd__o211a_1
X_16395_ _06342_ _06358_ VGND VGND VPWR VPWR _06593_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18134_ _07446_ _07453_ _07451_ VGND VGND VPWR VPWR _08506_ sky130_fd_sc_hd__a21oi_1
X_15346_ _05434_ _05436_ _05438_ VGND VGND VPWR VPWR _05439_ sky130_fd_sc_hd__a21o_1
X_12558_ _02478_ _02496_ VGND VGND VPWR VPWR _02497_ sky130_fd_sc_hd__xor2_1
XFILLER_0_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11509_ _01442_ _01445_ _01447_ VGND VGND VPWR VPWR _01448_ sky130_fd_sc_hd__o21a_1
X_18065_ _08167_ _08168_ _08429_ VGND VGND VPWR VPWR _08430_ sky130_fd_sc_hd__a21oi_2
X_15277_ _05275_ _05277_ VGND VGND VPWR VPWR _05363_ sky130_fd_sc_hd__or2_1
X_12489_ net254 _01759_ _02427_ VGND VGND VPWR VPWR _02428_ sky130_fd_sc_hd__and3_1
X_17016_ _07246_ _07275_ VGND VGND VPWR VPWR _07276_ sky130_fd_sc_hd__xnor2_2
X_14228_ _04147_ _04151_ _04208_ VGND VGND VPWR VPWR _04209_ sky130_fd_sc_hd__a21oi_2
X_14159_ _04130_ _04132_ VGND VGND VPWR VPWR _04133_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18967_ _09420_ _09421_ VGND VGND VPWR VPWR _09422_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17918_ net326 _07093_ _08267_ VGND VGND VPWR VPWR _08268_ sky130_fd_sc_hd__and3_1
X_18898_ _08886_ VGND VGND VPWR VPWR _09346_ sky130_fd_sc_hd__inv_2
X_17849_ _08190_ _08191_ VGND VGND VPWR VPWR _08192_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09967_ _05633_ _05655_ _06964_ VGND VGND VPWR VPWR _06986_ sky130_fd_sc_hd__o21a_1
X_09898_ net338 _06194_ _06216_ VGND VGND VPWR VPWR _06227_ sky130_fd_sc_hd__and3_1
X_11860_ _01798_ VGND VGND VPWR VPWR _01799_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10811_ _00663_ _00749_ VGND VGND VPWR VPWR _00750_ sky130_fd_sc_hd__xnor2_1
X_11791_ prev_error\[7\] _00226_ VGND VGND VPWR VPWR _01730_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13530_ _03384_ _03485_ _03480_ _03484_ VGND VGND VPWR VPWR _03489_ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10742_ _00590_ _00592_ VGND VGND VPWR VPWR _00681_ sky130_fd_sc_hd__xor2_1
XFILLER_0_82_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13461_ _03303_ _03332_ VGND VGND VPWR VPWR _03420_ sky130_fd_sc_hd__nor2_1
X_10673_ _04225_ _04269_ VGND VGND VPWR VPWR _00612_ sky130_fd_sc_hd__xor2_4
X_15200_ _05275_ _05277_ VGND VGND VPWR VPWR _05278_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12412_ _02349_ _02350_ VGND VGND VPWR VPWR _02351_ sky130_fd_sc_hd__and2b_1
XFILLER_0_35_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16180_ net283 _06346_ _06355_ VGND VGND VPWR VPWR _06356_ sky130_fd_sc_hd__and3_1
X_13392_ net265 _01852_ _03309_ VGND VGND VPWR VPWR _03346_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15131_ _05196_ _05190_ _05194_ VGND VGND VPWR VPWR _05202_ sky130_fd_sc_hd__or3_1
X_12343_ _02199_ _02281_ VGND VGND VPWR VPWR _02282_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12274_ net213 _01854_ _01861_ net217 VGND VGND VPWR VPWR _02213_ sky130_fd_sc_hd__a22o_1
X_15062_ _05013_ _05125_ VGND VGND VPWR VPWR _05126_ sky130_fd_sc_hd__xnor2_1
X_14013_ _03961_ _03962_ VGND VGND VPWR VPWR _03985_ sky130_fd_sc_hd__xnor2_1
X_11225_ _01144_ _01150_ _01151_ VGND VGND VPWR VPWR _01164_ sky130_fd_sc_hd__or3_1
XFILLER_0_120_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18821_ _03916_ _04200_ _09259_ VGND VGND VPWR VPWR _09261_ sky130_fd_sc_hd__or3b_1
X_11156_ _01089_ _01094_ VGND VGND VPWR VPWR _01095_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10107_ _07426_ _07503_ VGND VGND VPWR VPWR _08526_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18752_ _09177_ _09178_ VGND VGND VPWR VPWR _09185_ sky130_fd_sc_hd__and2b_1
X_15964_ _06034_ _06116_ _06118_ VGND VGND VPWR VPWR _06119_ sky130_fd_sc_hd__a21o_1
X_11087_ net565 _00515_ _00614_ net351 VGND VGND VPWR VPWR _01026_ sky130_fd_sc_hd__a22o_1
X_17703_ _08025_ _08030_ VGND VGND VPWR VPWR _08032_ sky130_fd_sc_hd__xnor2_1
X_10038_ _07393_ _07635_ VGND VGND VPWR VPWR _07767_ sky130_fd_sc_hd__xor2_2
X_14915_ _04960_ _04964_ net478 net131 VGND VGND VPWR VPWR _04965_ sky130_fd_sc_hd__and4bb_1
X_18683_ _06089_ _06091_ VGND VGND VPWR VPWR _09110_ sky130_fd_sc_hd__or2_1
X_15895_ _05967_ _06042_ VGND VGND VPWR VPWR _06043_ sky130_fd_sc_hd__and2_1
X_17634_ _07658_ _07663_ VGND VGND VPWR VPWR _07956_ sky130_fd_sc_hd__xnor2_1
X_14846_ _04887_ _04888_ VGND VGND VPWR VPWR _04889_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17565_ _07876_ VGND VGND VPWR VPWR _07880_ sky130_fd_sc_hd__inv_2
X_14777_ _04800_ _04810_ _04812_ VGND VGND VPWR VPWR _04813_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11989_ _01775_ _01927_ VGND VGND VPWR VPWR _01928_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19304_ clknet_4_7_0_clock _00044_ VGND VGND VPWR VPWR ki\[15\] sky130_fd_sc_hd__dfxtp_1
X_16516_ net279 net275 _06470_ _06621_ VGND VGND VPWR VPWR _06726_ sky130_fd_sc_hd__and4_1
XFILLER_0_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13728_ _03692_ _03693_ VGND VGND VPWR VPWR _03694_ sky130_fd_sc_hd__xnor2_1
X_17496_ net311 _06723_ _07802_ _07803_ VGND VGND VPWR VPWR _07804_ sky130_fd_sc_hd__a31o_1
XFILLER_0_85_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19235_ clknet_4_9_0_clock _00117_ VGND VGND VPWR VPWR i_error\[3\] sky130_fd_sc_hd__dfxtp_1
X_16447_ _06374_ _06591_ VGND VGND VPWR VPWR _06650_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_129_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13659_ _03616_ _03619_ VGND VGND VPWR VPWR _03621_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_140_Right_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19166_ net501 net464 VGND VGND VPWR VPWR _09579_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16378_ _06549_ _06558_ _06573_ VGND VGND VPWR VPWR _06574_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18117_ _08470_ _08474_ _08473_ VGND VGND VPWR VPWR _08487_ sky130_fd_sc_hd__a21o_1
XFILLER_0_26_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15329_ net441 net446 net189 net185 VGND VGND VPWR VPWR _05420_ sky130_fd_sc_hd__and4_1
X_19097_ net563 VGND VGND VPWR VPWR _09536_ sky130_fd_sc_hd__buf_4
XFILLER_0_124_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18048_ _08407_ _08408_ net110 _08409_ VGND VGND VPWR VPWR _08411_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_112_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout406 kp\[0\] VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__buf_4
Xfanout417 prev_d_error\[15\] VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__clkbuf_4
X_09821_ net356 net509 _05369_ VGND VGND VPWR VPWR _05380_ sky130_fd_sc_hd__and3_1
Xfanout428 net429 VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__clkbuf_4
Xfanout439 net440 VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__buf_2
X_09752_ net19 net77 VGND VGND VPWR VPWR _04621_ sky130_fd_sc_hd__nor2b_2
X_09683_ _03870_ VGND VGND VPWR VPWR _03881_ sky130_fd_sc_hd__buf_2
XFILLER_0_65_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout13 net335 VGND VGND VPWR VPWR net568 sky130_fd_sc_hd__buf_4
XFILLER_0_9_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11010_ _00919_ _00917_ VGND VGND VPWR VPWR _00949_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12961_ net228 _02090_ _02896_ _02899_ VGND VGND VPWR VPWR _02900_ sky130_fd_sc_hd__a31o_1
X_14700_ _04725_ _04727_ VGND VGND VPWR VPWR _04728_ sky130_fd_sc_hd__and2b_1
X_11912_ _01849_ _01850_ VGND VGND VPWR VPWR _01851_ sky130_fd_sc_hd__xnor2_4
X_15680_ _05794_ _05805_ VGND VGND VPWR VPWR _05806_ sky130_fd_sc_hd__nor2_1
X_12892_ _02816_ _02830_ VGND VGND VPWR VPWR _02831_ sky130_fd_sc_hd__xnor2_1
X_14631_ _04650_ _04651_ VGND VGND VPWR VPWR _04652_ sky130_fd_sc_hd__xnor2_1
X_11843_ _01777_ _01781_ VGND VGND VPWR VPWR _01782_ sky130_fd_sc_hd__or2b_1
XFILLER_0_157_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17350_ _07639_ _07642_ VGND VGND VPWR VPWR _07643_ sky130_fd_sc_hd__xor2_1
XFILLER_0_28_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14562_ _04564_ _04573_ _04575_ VGND VGND VPWR VPWR _04576_ sky130_fd_sc_hd__a21oi_1
X_11774_ prev_error\[3\] _00600_ VGND VGND VPWR VPWR _01713_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16301_ net292 _06377_ VGND VGND VPWR VPWR _06489_ sky130_fd_sc_hd__xor2_1
XFILLER_0_27_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13513_ _03469_ _03471_ VGND VGND VPWR VPWR _03472_ sky130_fd_sc_hd__and2b_1
XFILLER_0_153_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17281_ _02928_ _01717_ VGND VGND VPWR VPWR _07567_ sky130_fd_sc_hd__xor2_4
X_10725_ net387 net509 _05369_ VGND VGND VPWR VPWR _00664_ sky130_fd_sc_hd__and3_2
XFILLER_0_27_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14493_ _04494_ _04499_ VGND VGND VPWR VPWR _04501_ sky130_fd_sc_hd__and2_1
X_19020_ _09222_ _09479_ _09215_ VGND VGND VPWR VPWR _09480_ sky130_fd_sc_hd__and3b_1
XFILLER_0_83_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16232_ _06406_ _06411_ VGND VGND VPWR VPWR _06413_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13444_ net220 _02935_ VGND VGND VPWR VPWR _03403_ sky130_fd_sc_hd__nand2_1
X_10656_ _08086_ _00410_ _00524_ VGND VGND VPWR VPWR _00595_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_152_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16163_ net296 _06310_ _06320_ net300 VGND VGND VPWR VPWR _06338_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13375_ _03325_ _03326_ _03327_ VGND VGND VPWR VPWR _03328_ sky130_fd_sc_hd__nor3_1
X_10587_ _00502_ _00523_ _00525_ VGND VGND VPWR VPWR _00526_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_23_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15114_ _05181_ _05183_ VGND VGND VPWR VPWR _05184_ sky130_fd_sc_hd__nor2_1
X_12326_ net238 _01798_ VGND VGND VPWR VPWR _02265_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16094_ _06168_ _06131_ _06133_ _06170_ VGND VGND VPWR VPWR _06262_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15045_ _05106_ _05107_ net479 net139 VGND VGND VPWR VPWR _05108_ sky130_fd_sc_hd__and4bb_1
X_12257_ _02192_ _02195_ VGND VGND VPWR VPWR _02196_ sky130_fd_sc_hd__xnor2_1
X_11208_ net373 _00324_ _01146_ VGND VGND VPWR VPWR _01147_ sky130_fd_sc_hd__and3_1
X_12188_ net201 _01808_ VGND VGND VPWR VPWR _02127_ sky130_fd_sc_hd__nand2_1
X_18804_ _04172_ _04175_ _09240_ VGND VGND VPWR VPWR _09243_ sky130_fd_sc_hd__and3_1
X_11139_ _01062_ _01077_ VGND VGND VPWR VPWR _01078_ sky130_fd_sc_hd__nand2_1
X_16996_ net285 _06993_ VGND VGND VPWR VPWR _07254_ sky130_fd_sc_hd__nand2_1
X_15947_ _06067_ _06069_ VGND VGND VPWR VPWR _06100_ sky130_fd_sc_hd__xnor2_1
X_18735_ _06100_ _06075_ _06099_ VGND VGND VPWR VPWR _09167_ sky130_fd_sc_hd__nand3_1
X_18666_ _08936_ _09090_ _08963_ VGND VGND VPWR VPWR _09091_ sky130_fd_sc_hd__mux2_2
X_15878_ _03882_ _06023_ VGND VGND VPWR VPWR _06024_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14829_ net421 net186 _04565_ VGND VGND VPWR VPWR _04870_ sky130_fd_sc_hd__and3_1
X_17617_ net287 _02933_ VGND VGND VPWR VPWR _07937_ sky130_fd_sc_hd__nand2_1
X_18597_ _08762_ VGND VGND VPWR VPWR _09015_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17548_ _07854_ _07859_ _07515_ _07860_ VGND VGND VPWR VPWR _07861_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_86_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17479_ _07267_ _07269_ VGND VGND VPWR VPWR _07785_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19218_ clknet_4_4_0_clock _00100_ VGND VGND VPWR VPWR prev_error\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19149_ net507 net550 net495 _09568_ VGND VGND VPWR VPWR _00129_ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout203 net204 VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_4
Xfanout214 net215 VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout225 kd_1\[11\] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__buf_2
Xfanout236 net237 VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__clkbuf_4
X_09804_ _05182_ VGND VGND VPWR VPWR _05193_ sky130_fd_sc_hd__clkbuf_4
Xfanout247 kd_1\[5\] VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__clkbuf_4
Xfanout258 kd_1\[3\] VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout269 kd_1\[0\] VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__clkbuf_4
X_09735_ net16 net74 VGND VGND VPWR VPWR _04434_ sky130_fd_sc_hd__and2b_1
X_09666_ net53 _03625_ _03658_ ki\[4\] VGND VGND VPWR VPWR _00051_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09597_ net31 VGND VGND VPWR VPWR _02992_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10510_ _00436_ _00448_ VGND VGND VPWR VPWR _00449_ sky130_fd_sc_hd__or2_1
X_11490_ _01388_ _01390_ VGND VGND VPWR VPWR _01429_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10441_ _00294_ _00292_ VGND VGND VPWR VPWR _00380_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13160_ _03029_ _03109_ VGND VGND VPWR VPWR _03110_ sky130_fd_sc_hd__nor2_1
X_10372_ _00309_ _00310_ VGND VGND VPWR VPWR _00311_ sky130_fd_sc_hd__and2_1
X_12111_ _02046_ _02047_ _02049_ VGND VGND VPWR VPWR _02050_ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13091_ _03031_ _03033_ VGND VGND VPWR VPWR _03034_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12042_ _01980_ _01977_ _01975_ VGND VGND VPWR VPWR _01981_ sky130_fd_sc_hd__and3b_1
X_16850_ _02541_ _06280_ VGND VGND VPWR VPWR _07093_ sky130_fd_sc_hd__xnor2_4
X_15801_ _05785_ _05937_ _05676_ _05938_ VGND VGND VPWR VPWR _05939_ sky130_fd_sc_hd__o2bb2a_1
X_16781_ net324 _01755_ _06314_ VGND VGND VPWR VPWR _07017_ sky130_fd_sc_hd__and3_1
X_13993_ _03963_ _03964_ net434 net136 VGND VGND VPWR VPWR _03965_ sky130_fd_sc_hd__and4bb_1
X_18520_ _06265_ _06146_ VGND VGND VPWR VPWR _08930_ sky130_fd_sc_hd__and2b_1
X_15732_ _05830_ _05858_ _05862_ VGND VGND VPWR VPWR _05863_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12944_ net246 _01860_ _02882_ _02881_ VGND VGND VPWR VPWR _02883_ sky130_fd_sc_hd__a31o_1
XFILLER_0_153_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18451_ _08851_ _08853_ _08837_ _08833_ VGND VGND VPWR VPWR _08854_ sky130_fd_sc_hd__a22o_1
X_15663_ _05779_ _05786_ VGND VGND VPWR VPWR _05788_ sky130_fd_sc_hd__nand2_1
X_12875_ _02810_ _02811_ _02813_ VGND VGND VPWR VPWR _02814_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17402_ net317 _06309_ VGND VGND VPWR VPWR _07700_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14614_ _04612_ _04633_ VGND VGND VPWR VPWR _04634_ sky130_fd_sc_hd__or2_1
X_11826_ net268 net250 _01764_ _01762_ VGND VGND VPWR VPWR _01765_ sky130_fd_sc_hd__o211ai_4
X_18382_ _08776_ _06138_ VGND VGND VPWR VPWR _08778_ sky130_fd_sc_hd__nand2_1
X_15594_ _05679_ _05711_ VGND VGND VPWR VPWR _05712_ sky130_fd_sc_hd__or2b_1
XFILLER_0_96_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17333_ _07620_ _07623_ VGND VGND VPWR VPWR _07625_ sky130_fd_sc_hd__nor2_1
X_14545_ net567 net169 VGND VGND VPWR VPWR _04558_ sky130_fd_sc_hd__and2_1
X_11757_ _00268_ _00358_ _01694_ _01695_ VGND VGND VPWR VPWR _01696_ sky130_fd_sc_hd__a31o_4
X_17264_ _07545_ _07546_ _07499_ _07515_ VGND VGND VPWR VPWR _07549_ sky130_fd_sc_hd__a211oi_4
X_10708_ _00630_ _00646_ VGND VGND VPWR VPWR _00647_ sky130_fd_sc_hd__xnor2_2
X_14476_ _04481_ VGND VGND VPWR VPWR _04482_ sky130_fd_sc_hd__clkbuf_2
X_11688_ _01601_ _01600_ VGND VGND VPWR VPWR _01627_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19003_ _09183_ _09460_ VGND VGND VPWR VPWR _09462_ sky130_fd_sc_hd__xor2_2
XFILLER_0_141_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16215_ _06376_ _06394_ VGND VGND VPWR VPWR _06395_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13427_ _03320_ _03322_ _03321_ VGND VGND VPWR VPWR _03385_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17195_ net324 _06431_ _06434_ VGND VGND VPWR VPWR _07473_ sky130_fd_sc_hd__and3_1
X_10639_ _00492_ _00494_ VGND VGND VPWR VPWR _00578_ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16146_ _06316_ _06318_ VGND VGND VPWR VPWR _06319_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13358_ net265 _01859_ VGND VGND VPWR VPWR _03311_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12309_ _02237_ _02240_ _02246_ _02247_ VGND VGND VPWR VPWR _02248_ sky130_fd_sc_hd__o211a_1
X_16077_ _06240_ _06242_ VGND VGND VPWR VPWR _06243_ sky130_fd_sc_hd__xnor2_1
X_13289_ _03191_ _03241_ VGND VGND VPWR VPWR _03242_ sky130_fd_sc_hd__nand2_1
X_15028_ _04985_ _05003_ _05063_ VGND VGND VPWR VPWR _05089_ sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16979_ _07232_ _07234_ VGND VGND VPWR VPWR _07235_ sky130_fd_sc_hd__xor2_1
Xinput3 measurement[10] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
X_18718_ _09084_ _09137_ _09147_ VGND VGND VPWR VPWR _09148_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18649_ _09069_ _09071_ VGND VGND VPWR VPWR _09072_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09718_ net12 net70 VGND VGND VPWR VPWR _04247_ sky130_fd_sc_hd__xnor2_4
X_10990_ _00927_ _00834_ VGND VGND VPWR VPWR _00929_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09649_ net44 _03347_ _03380_ net215 VGND VGND VPWR VPWR _00004_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12660_ net234 _01860_ VGND VGND VPWR VPWR _02599_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11611_ net564 _00612_ VGND VGND VPWR VPWR _01550_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12591_ net199 _02419_ _02420_ VGND VGND VPWR VPWR _02530_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14330_ _04319_ _04320_ net434 net141 VGND VGND VPWR VPWR _04321_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_9_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11542_ _01453_ _01480_ VGND VGND VPWR VPWR _01481_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14261_ _04223_ _04227_ _04244_ VGND VGND VPWR VPWR _04245_ sky130_fd_sc_hd__a21o_1
X_11473_ net386 _00323_ VGND VGND VPWR VPWR _01412_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16000_ _06154_ _06157_ VGND VGND VPWR VPWR _06158_ sky130_fd_sc_hd__and2_1
X_13212_ _03163_ _03164_ VGND VGND VPWR VPWR _03165_ sky130_fd_sc_hd__and2_1
XFILLER_0_150_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10424_ _00362_ VGND VGND VPWR VPWR _00363_ sky130_fd_sc_hd__clkbuf_4
X_14192_ net408 net134 _04168_ _04165_ VGND VGND VPWR VPWR _04169_ sky130_fd_sc_hd__o2bb2a_1
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13143_ _03051_ _03082_ _03090_ VGND VGND VPWR VPWR _03092_ sky130_fd_sc_hd__and3_1
X_10355_ net364 _05325_ _00293_ VGND VGND VPWR VPWR _00294_ sky130_fd_sc_hd__and3_1
XFILLER_0_148_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13074_ _03011_ _02887_ _03012_ _03015_ VGND VGND VPWR VPWR _03016_ sky130_fd_sc_hd__o22a_1
X_17951_ _08212_ _08213_ VGND VGND VPWR VPWR _08304_ sky130_fd_sc_hd__xnor2_2
X_10286_ _00223_ _00224_ VGND VGND VPWR VPWR _00225_ sky130_fd_sc_hd__xnor2_1
X_16902_ _07148_ _07147_ VGND VGND VPWR VPWR _07150_ sky130_fd_sc_hd__or2b_1
X_12025_ _01881_ _01887_ _01963_ VGND VGND VPWR VPWR _01964_ sky130_fd_sc_hd__a21bo_1
X_17882_ _08224_ _08225_ _08227_ VGND VGND VPWR VPWR _08228_ sky130_fd_sc_hd__o21ba_1
X_16833_ net282 _06724_ VGND VGND VPWR VPWR _07075_ sky130_fd_sc_hd__nand2_1
X_16764_ _06990_ _06998_ VGND VGND VPWR VPWR _06999_ sky130_fd_sc_hd__nand2_1
X_13976_ _03944_ _03947_ VGND VGND VPWR VPWR _03948_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15715_ _05803_ _05844_ VGND VGND VPWR VPWR _05845_ sky130_fd_sc_hd__nor2_1
X_18503_ _06266_ _08840_ VGND VGND VPWR VPWR _08912_ sky130_fd_sc_hd__nor2_1
X_12927_ _02835_ _02865_ VGND VGND VPWR VPWR _02866_ sky130_fd_sc_hd__and2_1
X_16695_ _06905_ _06922_ VGND VGND VPWR VPWR _06923_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15646_ _05756_ _05767_ _05768_ VGND VGND VPWR VPWR _05769_ sky130_fd_sc_hd__nand3_1
X_18434_ _06163_ _08835_ VGND VGND VPWR VPWR _08836_ sky130_fd_sc_hd__nand2_1
X_12858_ _02796_ _02704_ VGND VGND VPWR VPWR _02797_ sky130_fd_sc_hd__xor2_2
XFILLER_0_56_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18365_ _06166_ _06168_ VGND VGND VPWR VPWR _08760_ sky130_fd_sc_hd__nor2_1
X_11809_ _01745_ _01746_ _01747_ VGND VGND VPWR VPWR _01748_ sky130_fd_sc_hd__a21oi_4
X_15577_ _05685_ _05692_ VGND VGND VPWR VPWR _05693_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12789_ _02718_ _02727_ VGND VGND VPWR VPWR _02728_ sky130_fd_sc_hd__xor2_1
XFILLER_0_138_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17316_ _07519_ _07521_ VGND VGND VPWR VPWR _07606_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14528_ _04527_ _04529_ _04538_ VGND VGND VPWR VPWR _04539_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18296_ _08529_ _08534_ _08611_ _08612_ _08527_ VGND VGND VPWR VPWR _08684_ sky130_fd_sc_hd__a311o_1
XFILLER_0_22_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17247_ _07523_ _07524_ _07528_ _07529_ VGND VGND VPWR VPWR _07530_ sky130_fd_sc_hd__nand4_1
XFILLER_0_141_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14459_ _04441_ _04462_ VGND VGND VPWR VPWR _04463_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17178_ _07446_ _07453_ VGND VGND VPWR VPWR _07454_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16129_ _06298_ _01742_ _06299_ _01811_ VGND VGND VPWR VPWR _06300_ sky130_fd_sc_hd__and4_1
XFILLER_0_110_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_30 kp\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10140_ _08878_ VGND VGND VPWR VPWR _08889_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10071_ _08075_ _08119_ VGND VGND VPWR VPWR _08130_ sky130_fd_sc_hd__xnor2_1
X_13830_ _03762_ _03792_ _03793_ _03795_ VGND VGND VPWR VPWR _03796_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_43_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13761_ _03723_ _03726_ VGND VGND VPWR VPWR _03727_ sky130_fd_sc_hd__nor2_1
X_10973_ _00911_ _00816_ VGND VGND VPWR VPWR _00912_ sky130_fd_sc_hd__or2_1
X_15500_ _05591_ _05598_ _05607_ VGND VGND VPWR VPWR _05608_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12712_ net202 _02546_ VGND VGND VPWR VPWR _02651_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16480_ _06685_ _06602_ VGND VGND VPWR VPWR _06686_ sky130_fd_sc_hd__xnor2_2
X_13692_ _03628_ _03630_ VGND VGND VPWR VPWR _03657_ sky130_fd_sc_hd__xor2_1
X_15431_ _05530_ _05531_ VGND VGND VPWR VPWR _05532_ sky130_fd_sc_hd__and2_1
X_12643_ _02429_ _02581_ VGND VGND VPWR VPWR _02582_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18150_ _06751_ _06835_ VGND VGND VPWR VPWR _08523_ sky130_fd_sc_hd__and2b_1
X_15362_ _05387_ _05448_ _05455_ VGND VGND VPWR VPWR _05456_ sky130_fd_sc_hd__o21ai_1
X_12574_ net209 _02091_ VGND VGND VPWR VPWR _02513_ sky130_fd_sc_hd__nand2_1
X_17101_ net294 _06468_ _07070_ VGND VGND VPWR VPWR _07369_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_136_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14313_ _04296_ _04289_ _04294_ VGND VGND VPWR VPWR _04303_ sky130_fd_sc_hd__nor3_1
XFILLER_0_136_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11525_ _01462_ _01463_ VGND VGND VPWR VPWR _01464_ sky130_fd_sc_hd__xnor2_1
X_18081_ _08443_ _08445_ VGND VGND VPWR VPWR _08447_ sky130_fd_sc_hd__xor2_2
XFILLER_0_151_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15293_ _05299_ _05377_ _05379_ VGND VGND VPWR VPWR _05381_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17032_ _07291_ _06321_ _06322_ _07292_ VGND VGND VPWR VPWR _07293_ sky130_fd_sc_hd__o31a_1
X_14244_ _04218_ _04221_ _04226_ VGND VGND VPWR VPWR _04227_ sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_12_Left_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11456_ _01237_ _01394_ VGND VGND VPWR VPWR _01395_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10407_ _00344_ _00345_ VGND VGND VPWR VPWR _00346_ sky130_fd_sc_hd__and2_1
X_14175_ _04124_ _04125_ _04150_ VGND VGND VPWR VPWR _04151_ sky130_fd_sc_hd__or3_2
XFILLER_0_1_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11387_ _01260_ _01318_ _01322_ VGND VGND VPWR VPWR _01326_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13126_ _03053_ _03072_ VGND VGND VPWR VPWR _03073_ sky130_fd_sc_hd__xnor2_1
X_10338_ net384 _07294_ net539 _05534_ VGND VGND VPWR VPWR _00277_ sky130_fd_sc_hd__a31o_1
X_18983_ _08885_ VGND VGND VPWR VPWR _09440_ sky130_fd_sc_hd__inv_2
X_13057_ net256 _01859_ _01834_ net260 VGND VGND VPWR VPWR _02997_ sky130_fd_sc_hd__a22o_1
X_17934_ _06544_ _08285_ _08276_ VGND VGND VPWR VPWR _08286_ sky130_fd_sc_hd__o21ai_1
X_10269_ net365 _05325_ _05424_ net368 VGND VGND VPWR VPWR _00208_ sky130_fd_sc_hd__a22oi_1
X_12008_ _01945_ _01946_ VGND VGND VPWR VPWR _01947_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17865_ _08205_ _08206_ _08209_ VGND VGND VPWR VPWR _08210_ sky130_fd_sc_hd__a21o_1
X_16816_ net309 _06352_ VGND VGND VPWR VPWR _07056_ sky130_fd_sc_hd__nand2_1
X_17796_ _08117_ _08133_ VGND VGND VPWR VPWR _08134_ sky130_fd_sc_hd__nor2_1
X_16747_ net288 _06620_ VGND VGND VPWR VPWR _06980_ sky130_fd_sc_hd__and2_1
X_13959_ net426 net567 net133 net128 VGND VGND VPWR VPWR _03931_ sky130_fd_sc_hd__and4_1
XFILLER_0_88_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16678_ _06878_ _06903_ VGND VGND VPWR VPWR _06904_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_29_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18417_ _06158_ _08816_ VGND VGND VPWR VPWR _08817_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15629_ _05742_ _05738_ _05740_ VGND VGND VPWR VPWR _05750_ sky130_fd_sc_hd__or3_1
XFILLER_0_57_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18348_ _06131_ _08740_ VGND VGND VPWR VPWR _08741_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18279_ _08663_ _08664_ VGND VGND VPWR VPWR _08665_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput50 reg_data[1] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput61 target[10] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_1
Xinput72 target[3] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09983_ _07140_ _07151_ VGND VGND VPWR VPWR _07162_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_149_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_154_Right_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11310_ _01188_ _01189_ _01187_ VGND VGND VPWR VPWR _01249_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_132_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12290_ _02215_ _02216_ VGND VGND VPWR VPWR _02229_ sky130_fd_sc_hd__xor2_1
XFILLER_0_121_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11241_ net392 _01178_ _01179_ VGND VGND VPWR VPWR _01180_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11172_ net343 _00812_ _01110_ VGND VGND VPWR VPWR _01111_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10123_ _07019_ _07129_ _07107_ VGND VGND VPWR VPWR _08702_ sky130_fd_sc_hd__a21oi_1
X_15980_ _00959_ net103 VGND VGND VPWR VPWR _06136_ sky130_fd_sc_hd__xor2_4
X_10054_ _06469_ _06491_ VGND VGND VPWR VPWR _07943_ sky130_fd_sc_hd__xnor2_1
X_14931_ _04826_ _04957_ VGND VGND VPWR VPWR _04982_ sky130_fd_sc_hd__nand2_1
X_14862_ _04903_ _04904_ _04905_ VGND VGND VPWR VPWR _04906_ sky130_fd_sc_hd__o21ba_1
X_17650_ _07798_ _07883_ VGND VGND VPWR VPWR _07973_ sky130_fd_sc_hd__nand2_1
X_16601_ _06797_ _06818_ VGND VGND VPWR VPWR _06819_ sky130_fd_sc_hd__xnor2_1
X_13813_ _03778_ VGND VGND VPWR VPWR _03779_ sky130_fd_sc_hd__inv_2
X_17581_ net332 _06718_ _06719_ VGND VGND VPWR VPWR _07897_ sky130_fd_sc_hd__and3_1
X_14793_ net445 net159 net154 net449 VGND VGND VPWR VPWR _04831_ sky130_fd_sc_hd__a22oi_1
XPHY_EDGE_ROW_121_Right_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16532_ _06735_ _06709_ VGND VGND VPWR VPWR _06743_ sky130_fd_sc_hd__or2b_1
X_19320_ clknet_4_1_0_clock _00003_ VGND VGND VPWR VPWR kd_1\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13744_ _03653_ _03704_ _03690_ _03703_ VGND VGND VPWR VPWR _03710_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_98_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10956_ _00884_ _00894_ VGND VGND VPWR VPWR _00895_ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19251_ clknet_4_11_0_clock _00133_ VGND VGND VPWR VPWR prev_d_error\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16463_ _06589_ _06666_ VGND VGND VPWR VPWR _06668_ sky130_fd_sc_hd__nor2_1
X_13675_ net256 _02543_ _02407_ net260 VGND VGND VPWR VPWR _03639_ sky130_fd_sc_hd__a22oi_1
X_10887_ _00818_ _00825_ net568 VGND VGND VPWR VPWR _00826_ sky130_fd_sc_hd__and3b_2
X_15414_ _05511_ _05513_ VGND VGND VPWR VPWR _05514_ sky130_fd_sc_hd__and2_1
X_18202_ _08499_ _08481_ _08540_ VGND VGND VPWR VPWR _08580_ sky130_fd_sc_hd__or3_1
X_12626_ _02421_ _02529_ _02530_ _02564_ VGND VGND VPWR VPWR _02565_ sky130_fd_sc_hd__o31ai_2
X_19182_ net507 net427 VGND VGND VPWR VPWR _09588_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16394_ _06591_ _06374_ VGND VGND VPWR VPWR _06592_ sky130_fd_sc_hd__and2b_1
X_18133_ _08503_ _07149_ VGND VGND VPWR VPWR _08505_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15345_ _05350_ _05437_ VGND VGND VPWR VPWR _05438_ sky130_fd_sc_hd__or2_1
X_12557_ net246 _01799_ VGND VGND VPWR VPWR _02496_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18064_ _08162_ _08223_ _08426_ _08428_ VGND VGND VPWR VPWR _08429_ sky130_fd_sc_hd__o22a_1
X_11508_ _01369_ _01446_ VGND VGND VPWR VPWR _01447_ sky130_fd_sc_hd__xnor2_1
X_15276_ _05301_ _05361_ VGND VGND VPWR VPWR _05362_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12488_ net259 net111 VGND VGND VPWR VPWR _02427_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17015_ _07192_ _07247_ VGND VGND VPWR VPWR _07275_ sky130_fd_sc_hd__nor2_1
X_14227_ _04206_ _04207_ VGND VGND VPWR VPWR _04208_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11439_ net395 _09558_ _09565_ _01376_ VGND VGND VPWR VPWR _01378_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14158_ net122 _04131_ VGND VGND VPWR VPWR _04132_ sky130_fd_sc_hd__and2_1
X_13109_ _02927_ _02937_ _02938_ VGND VGND VPWR VPWR _03054_ sky130_fd_sc_hd__and3_1
X_18966_ prev_d_error\[18\] _04961_ _09244_ _09242_ VGND VGND VPWR VPWR _09421_ sky130_fd_sc_hd__a31o_1
X_14089_ _04059_ _04060_ VGND VGND VPWR VPWR _04061_ sky130_fd_sc_hd__nor2_1
X_17917_ _08226_ _08266_ VGND VGND VPWR VPWR _08267_ sky130_fd_sc_hd__xor2_1
X_18897_ _09343_ _09344_ VGND VGND VPWR VPWR _09345_ sky130_fd_sc_hd__xnor2_4
X_17848_ _08085_ _08087_ _08084_ VGND VGND VPWR VPWR _08191_ sky130_fd_sc_hd__o21a_1
X_17779_ _08104_ _08105_ _08114_ VGND VGND VPWR VPWR _08115_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09966_ _05666_ _06964_ VGND VGND VPWR VPWR _06975_ sky130_fd_sc_hd__xnor2_1
X_09897_ _06139_ _06205_ VGND VGND VPWR VPWR _06216_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10810_ _00720_ _00747_ _00748_ VGND VGND VPWR VPWR _00749_ sky130_fd_sc_hd__a21oi_1
X_11790_ prev_error\[7\] _00226_ VGND VGND VPWR VPWR _01729_ sky130_fd_sc_hd__nand2_2
XFILLER_0_156_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10741_ _00672_ _00678_ _00679_ VGND VGND VPWR VPWR _00680_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_149_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13460_ _03411_ _03413_ _03418_ VGND VGND VPWR VPWR _03419_ sky130_fd_sc_hd__or3_1
X_10672_ _00604_ _00607_ _00610_ VGND VGND VPWR VPWR _00611_ sky130_fd_sc_hd__o21a_1
XFILLER_0_137_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12411_ _02307_ _02309_ _02341_ VGND VGND VPWR VPWR _02350_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_153_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13391_ _03325_ _03326_ _03327_ VGND VGND VPWR VPWR _03345_ sky130_fd_sc_hd__o21a_1
XFILLER_0_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15130_ _05190_ _05194_ _05196_ VGND VGND VPWR VPWR _05201_ sky130_fd_sc_hd__o21ai_1
X_12342_ _02196_ _02198_ VGND VGND VPWR VPWR _02281_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15061_ _05015_ _05014_ VGND VGND VPWR VPWR _05125_ sky130_fd_sc_hd__nor2_1
X_12273_ _02097_ _02211_ VGND VGND VPWR VPWR _02212_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14012_ _03982_ _03970_ _03977_ VGND VGND VPWR VPWR _03984_ sky130_fd_sc_hd__nor3_1
XFILLER_0_121_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11224_ _01160_ _01162_ _01158_ VGND VGND VPWR VPWR _01163_ sky130_fd_sc_hd__a21oi_4
X_18820_ _03916_ _04200_ _09259_ VGND VGND VPWR VPWR _09260_ sky130_fd_sc_hd__o21ba_1
X_11155_ _01090_ _01093_ _01091_ VGND VGND VPWR VPWR _01094_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_156_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10106_ _06997_ _07195_ _07228_ VGND VGND VPWR VPWR _08515_ sky130_fd_sc_hd__a21bo_1
X_18751_ _09150_ _09165_ _09179_ _09183_ VGND VGND VPWR VPWR _09184_ sky130_fd_sc_hd__nand4bb_2
X_15963_ _06024_ _06027_ VGND VGND VPWR VPWR _06118_ sky130_fd_sc_hd__xnor2_1
X_11086_ _01024_ _00903_ VGND VGND VPWR VPWR _01025_ sky130_fd_sc_hd__or2_1
X_17702_ _08028_ _08029_ VGND VGND VPWR VPWR _08030_ sky130_fd_sc_hd__nor2_1
X_10037_ _07745_ VGND VGND VPWR VPWR _07756_ sky130_fd_sc_hd__inv_2
X_14914_ net469 net138 _04961_ _04963_ VGND VGND VPWR VPWR _04964_ sky130_fd_sc_hd__o2bb2a_1
X_15894_ _05966_ _05960_ _05964_ VGND VGND VPWR VPWR _06042_ sky130_fd_sc_hd__nand3_1
X_18682_ _06148_ VGND VGND VPWR VPWR _09108_ sky130_fd_sc_hd__inv_2
X_17633_ _07945_ _07953_ VGND VGND VPWR VPWR _07955_ sky130_fd_sc_hd__nor2_1
X_14845_ _04886_ _04854_ _04883_ VGND VGND VPWR VPWR _04888_ sky130_fd_sc_hd__or3_1
X_14776_ _04696_ _04811_ VGND VGND VPWR VPWR _04812_ sky130_fd_sc_hd__nand2_1
X_17564_ _07839_ _07876_ _07878_ VGND VGND VPWR VPWR _07879_ sky130_fd_sc_hd__and3_1
X_11988_ _01777_ _01926_ VGND VGND VPWR VPWR _01927_ sky130_fd_sc_hd__or2b_1
XFILLER_0_129_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19303_ clknet_4_7_0_clock _00043_ VGND VGND VPWR VPWR ki\[14\] sky130_fd_sc_hd__dfxtp_2
X_16515_ net279 _06470_ _06621_ net276 VGND VGND VPWR VPWR _06725_ sky130_fd_sc_hd__a22o_1
X_13727_ _03566_ _03624_ _03623_ VGND VGND VPWR VPWR _03693_ sky130_fd_sc_hd__o21a_1
XFILLER_0_156_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10939_ _00874_ _00876_ VGND VGND VPWR VPWR _00878_ sky130_fd_sc_hd__xnor2_1
X_17495_ net332 net315 _06408_ _06619_ VGND VGND VPWR VPWR _07803_ sky130_fd_sc_hd__and4_1
XFILLER_0_129_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19234_ clknet_4_9_0_clock _00116_ VGND VGND VPWR VPWR i_error\[2\] sky130_fd_sc_hd__dfxtp_1
X_13658_ _03616_ _03619_ VGND VGND VPWR VPWR _03620_ sky130_fd_sc_hd__nand2_1
X_16446_ _06542_ _06547_ net106 VGND VGND VPWR VPWR _06649_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_116_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12609_ _02404_ _02547_ VGND VGND VPWR VPWR _02548_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19165_ _09559_ _09168_ _09578_ net490 VGND VGND VPWR VPWR _00137_ sky130_fd_sc_hd__o211a_1
X_16377_ _06555_ _06572_ VGND VGND VPWR VPWR _06573_ sky130_fd_sc_hd__xor2_1
XFILLER_0_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13589_ _03523_ _03546_ _03547_ VGND VGND VPWR VPWR _03548_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15328_ _05401_ _05417_ _05418_ VGND VGND VPWR VPWR _05419_ sky130_fd_sc_hd__a21bo_1
X_18116_ _07796_ _07766_ VGND VGND VPWR VPWR _08486_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19096_ _09523_ _06645_ _09535_ net488 VGND VGND VPWR VPWR _00104_ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15259_ _05241_ _05342_ VGND VGND VPWR VPWR _05343_ sky130_fd_sc_hd__xnor2_1
X_18047_ _08407_ _08408_ net110 _08409_ VGND VGND VPWR VPWR _08410_ sky130_fd_sc_hd__a211o_1
XFILLER_0_41_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout407 net410 VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__buf_2
XFILLER_0_1_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09820_ _04709_ _04731_ _04753_ _05358_ _04720_ VGND VGND VPWR VPWR _05369_ sky130_fd_sc_hd__o2111ai_4
Xfanout418 net419 VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__buf_2
XFILLER_0_39_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout429 prev_d_error\[13\] VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__buf_2
XFILLER_0_10_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09751_ _04566_ _04599_ VGND VGND VPWR VPWR _04610_ sky130_fd_sc_hd__or2_1
X_18949_ _09381_ _09401_ VGND VGND VPWR VPWR _09402_ sky130_fd_sc_hd__xnor2_1
X_09682_ net79 _03859_ VGND VGND VPWR VPWR _03870_ sky130_fd_sc_hd__nor2_4
XFILLER_0_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09949_ _05875_ _06436_ _06777_ VGND VGND VPWR VPWR _06788_ sky130_fd_sc_hd__a21bo_1
X_12960_ net224 _02331_ _02898_ VGND VGND VPWR VPWR _02899_ sky130_fd_sc_hd__and3_1
X_11911_ _01707_ _01734_ _01735_ VGND VGND VPWR VPWR _01850_ sky130_fd_sc_hd__o21ai_2
X_12891_ _02827_ _02829_ _02825_ VGND VGND VPWR VPWR _02830_ sky130_fd_sc_hd__a21oi_1
X_14630_ _04606_ _04609_ VGND VGND VPWR VPWR _04651_ sky130_fd_sc_hd__nor2_1
X_11842_ _01769_ _01780_ VGND VGND VPWR VPWR _01781_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14561_ _04546_ _04574_ VGND VGND VPWR VPWR _04575_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11773_ _00406_ _00407_ _01711_ VGND VGND VPWR VPWR _01712_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13512_ _03470_ _03351_ VGND VGND VPWR VPWR _03471_ sky130_fd_sc_hd__xnor2_1
X_16300_ _06384_ _06393_ _06383_ VGND VGND VPWR VPWR _06488_ sky130_fd_sc_hd__a21bo_1
X_17280_ _07563_ _07564_ VGND VGND VPWR VPWR _07566_ sky130_fd_sc_hd__nand2_1
X_10724_ _00626_ _00652_ VGND VGND VPWR VPWR _00663_ sky130_fd_sc_hd__xnor2_1
X_14492_ _04483_ _04486_ _04493_ VGND VGND VPWR VPWR _04499_ sky130_fd_sc_hd__or3_1
XFILLER_0_82_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16231_ _06406_ _06411_ VGND VGND VPWR VPWR _06412_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13443_ _03400_ _03401_ VGND VGND VPWR VPWR _03402_ sky130_fd_sc_hd__nor2_1
X_10655_ _00580_ _00593_ VGND VGND VPWR VPWR _00594_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16162_ _06335_ VGND VGND VPWR VPWR _06336_ sky130_fd_sc_hd__buf_2
XFILLER_0_23_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13374_ _03297_ _03299_ VGND VGND VPWR VPWR _03327_ sky130_fd_sc_hd__xnor2_1
X_10586_ _00410_ _00524_ net568 VGND VGND VPWR VPWR _00525_ sky130_fd_sc_hd__and3b_1
X_15113_ _05158_ _05162_ _05180_ VGND VGND VPWR VPWR _05183_ sky130_fd_sc_hd__nor3_1
XFILLER_0_134_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12325_ _02262_ _02263_ VGND VGND VPWR VPWR _02264_ sky130_fd_sc_hd__nor2_1
X_16093_ _06229_ _06259_ VGND VGND VPWR VPWR _06261_ sky130_fd_sc_hd__xnor2_4
X_15044_ net471 net149 net143 net476 VGND VGND VPWR VPWR _05107_ sky130_fd_sc_hd__a22oi_1
X_12256_ net221 _01836_ _02193_ _02194_ VGND VGND VPWR VPWR _02195_ sky130_fd_sc_hd__a31o_1
X_11207_ _01145_ _01065_ VGND VGND VPWR VPWR _01146_ sky130_fd_sc_hd__xor2_1
X_12187_ net200 _01836_ _01959_ _02125_ VGND VGND VPWR VPWR _02126_ sky130_fd_sc_hd__a31o_1
X_18803_ _04172_ _04175_ _09240_ VGND VGND VPWR VPWR _09242_ sky130_fd_sc_hd__a21oi_1
X_11138_ _01075_ _01076_ VGND VGND VPWR VPWR _01077_ sky130_fd_sc_hd__nor2_2
X_16995_ _07174_ _07252_ VGND VGND VPWR VPWR _07253_ sky130_fd_sc_hd__nor2_1
X_18734_ _06155_ _06156_ VGND VGND VPWR VPWR _09166_ sky130_fd_sc_hd__xor2_4
X_15946_ _06080_ _06096_ _06098_ VGND VGND VPWR VPWR _06099_ sky130_fd_sc_hd__a21o_1
X_11069_ _00906_ _01007_ VGND VGND VPWR VPWR _01008_ sky130_fd_sc_hd__nor2_1
X_18665_ _08811_ _08815_ _08881_ VGND VGND VPWR VPWR _09090_ sky130_fd_sc_hd__mux2_1
X_15877_ _03880_ _02673_ _03879_ VGND VGND VPWR VPWR _06023_ sky130_fd_sc_hd__and3_1
XFILLER_0_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17616_ _07934_ _07935_ VGND VGND VPWR VPWR _07936_ sky130_fd_sc_hd__nor2_1
X_14828_ net417 net186 net182 net424 VGND VGND VPWR VPWR _04869_ sky130_fd_sc_hd__a22o_1
X_18596_ _08899_ VGND VGND VPWR VPWR _09014_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17547_ _07499_ _07513_ _07512_ VGND VGND VPWR VPWR _07860_ sky130_fd_sc_hd__o21a_1
X_14759_ net475 net124 _04683_ _04684_ VGND VGND VPWR VPWR _04793_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_46_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17478_ _07715_ _07728_ _07783_ VGND VGND VPWR VPWR _07784_ sky130_fd_sc_hd__a21oi_2
X_19217_ clknet_4_4_0_clock _00099_ VGND VGND VPWR VPWR prev_error\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16429_ _06453_ _06627_ VGND VGND VPWR VPWR _06630_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_4_Left_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19148_ net507 _08976_ VGND VGND VPWR VPWR _09568_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19079_ net498 prev_error\[1\] VGND VGND VPWR VPWR _09525_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout204 kd_1\[16\] VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_4
Xfanout215 kd_1\[13\] VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_4
Xfanout226 net227 VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__buf_2
X_09803_ _05171_ VGND VGND VPWR VPWR _05182_ sky130_fd_sc_hd__clkbuf_4
Xfanout237 kd_1\[8\] VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__clkbuf_4
Xfanout248 net249 VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout259 net261 VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__buf_2
X_09734_ _04192_ _04313_ _04346_ _04379_ _04412_ VGND VGND VPWR VPWR _04423_ sky130_fd_sc_hd__a2111o_4
XFILLER_0_97_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09665_ net52 _03625_ _03658_ net321 VGND VGND VPWR VPWR _00050_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10440_ _00375_ _00377_ VGND VGND VPWR VPWR _00379_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10371_ _00305_ _00306_ VGND VGND VPWR VPWR _00310_ sky130_fd_sc_hd__xor2_1
XFILLER_0_33_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12110_ _01843_ _02048_ VGND VGND VPWR VPWR _02049_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13090_ _02922_ _03032_ VGND VGND VPWR VPWR _03033_ sky130_fd_sc_hd__nor2_1
X_12041_ net264 net259 net254 _01764_ VGND VGND VPWR VPWR _01980_ sky130_fd_sc_hd__o31a_1
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15800_ _05730_ _05784_ _05734_ VGND VGND VPWR VPWR _05938_ sky130_fd_sc_hd__or3_1
X_13992_ net438 net132 net127 net443 VGND VGND VPWR VPWR _03964_ sky130_fd_sc_hd__a22oi_1
X_16780_ _07014_ net329 _07015_ VGND VGND VPWR VPWR _07016_ sky130_fd_sc_hd__mux2_1
X_15731_ _05860_ _05861_ VGND VGND VPWR VPWR _05862_ sky130_fd_sc_hd__nor2_1
X_12943_ _02879_ _02881_ VGND VGND VPWR VPWR _02882_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18450_ _08852_ _08743_ VGND VGND VPWR VPWR _08853_ sky130_fd_sc_hd__nor2_1
X_15662_ _05772_ _05778_ _05777_ VGND VGND VPWR VPWR _05786_ sky130_fd_sc_hd__o21ai_1
X_12874_ _02812_ _02725_ VGND VGND VPWR VPWR _02813_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17401_ _07621_ _07622_ _07625_ VGND VGND VPWR VPWR _07699_ sky130_fd_sc_hd__o21bai_2
X_11825_ _01759_ VGND VGND VPWR VPWR _01764_ sky130_fd_sc_hd__clkbuf_4
X_14613_ _04613_ _04631_ _04629_ VGND VGND VPWR VPWR _04633_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15593_ _05697_ _05709_ VGND VGND VPWR VPWR _05711_ sky130_fd_sc_hd__nand2_1
X_18381_ _08776_ _06138_ VGND VGND VPWR VPWR _08777_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14544_ _04016_ net182 VGND VGND VPWR VPWR _04557_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17332_ _07621_ _07622_ VGND VGND VPWR VPWR _07623_ sky130_fd_sc_hd__xnor2_1
X_11756_ _00265_ _00356_ _00267_ VGND VGND VPWR VPWR _01695_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10707_ _00632_ _00644_ _00645_ VGND VGND VPWR VPWR _00646_ sky130_fd_sc_hd__a21o_1
X_14475_ net485 net117 VGND VGND VPWR VPWR _04481_ sky130_fd_sc_hd__and2_1
X_17263_ _07499_ _07515_ _07545_ _07546_ VGND VGND VPWR VPWR _07548_ sky130_fd_sc_hd__o211a_4
X_11687_ _01617_ _01621_ _01625_ VGND VGND VPWR VPWR _01626_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19002_ _09185_ _09453_ VGND VGND VPWR VPWR _09460_ sky130_fd_sc_hd__nor2_1
X_13426_ _03368_ _03382_ _03383_ VGND VGND VPWR VPWR _03384_ sky130_fd_sc_hd__nor3_2
X_16214_ _06385_ _06393_ VGND VGND VPWR VPWR _06394_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17194_ net323 _06400_ _06435_ net319 VGND VGND VPWR VPWR _07472_ sky130_fd_sc_hd__a22o_1
X_10638_ _00569_ _00571_ _00576_ VGND VGND VPWR VPWR _00577_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16145_ _06317_ VGND VGND VPWR VPWR _06318_ sky130_fd_sc_hd__clkbuf_4
X_13357_ net265 _01852_ _03309_ VGND VGND VPWR VPWR _03310_ sky130_fd_sc_hd__and3_1
XFILLER_0_106_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10569_ net337 _00410_ VGND VGND VPWR VPWR _00508_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12308_ _02111_ _02245_ _02209_ _02244_ VGND VGND VPWR VPWR _02247_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_87_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16076_ _05666_ _06204_ _06241_ VGND VGND VPWR VPWR _06242_ sky130_fd_sc_hd__o21a_1
X_13288_ net248 _01908_ _03190_ VGND VGND VPWR VPWR _03241_ sky130_fd_sc_hd__a21o_1
XFILLER_0_122_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15027_ _05086_ _05078_ _05081_ VGND VGND VPWR VPWR _05088_ sky130_fd_sc_hd__or3_1
X_12239_ _02175_ _02176_ _02177_ VGND VGND VPWR VPWR _02178_ sky130_fd_sc_hd__o21ba_1
X_16978_ _07069_ _07193_ _07233_ VGND VGND VPWR VPWR _07234_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput4 measurement[11] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
X_18717_ _06138_ _09145_ _09146_ VGND VGND VPWR VPWR _09147_ sky130_fd_sc_hd__a21bo_1
X_15929_ _06077_ _06079_ VGND VGND VPWR VPWR _06080_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18648_ _06162_ _09068_ VGND VGND VPWR VPWR _09071_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18579_ _08992_ _08994_ VGND VGND VPWR VPWR _08995_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_49_Left_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_58_Left_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09717_ net60 net2 VGND VGND VPWR VPWR _04236_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_97_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09648_ net43 _03347_ _03380_ net218 VGND VGND VPWR VPWR _00003_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_67_Left_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11610_ net385 _00613_ VGND VGND VPWR VPWR _01549_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12590_ _02520_ _02523_ VGND VGND VPWR VPWR _02529_ sky130_fd_sc_hd__nor2_2
XFILLER_0_107_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11541_ _01450_ _01452_ VGND VGND VPWR VPWR _01480_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14260_ _03977_ _04243_ VGND VGND VPWR VPWR _04244_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11472_ _01354_ _01406_ VGND VGND VPWR VPWR _01411_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13211_ _03142_ _03160_ VGND VGND VPWR VPWR _03164_ sky130_fd_sc_hd__xor2_1
X_10423_ net405 _05512_ _05523_ VGND VGND VPWR VPWR _00362_ sky130_fd_sc_hd__and3_1
X_14191_ _04166_ VGND VGND VPWR VPWR _04168_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13142_ _03083_ VGND VGND VPWR VPWR _03090_ sky130_fd_sc_hd__inv_2
X_10354_ net368 net510 _06029_ VGND VGND VPWR VPWR _00293_ sky130_fd_sc_hd__and3_1
XFILLER_0_104_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_76_Left_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13073_ _03011_ _02887_ _03013_ VGND VGND VPWR VPWR _03015_ sky130_fd_sc_hd__o21ai_1
X_17950_ net298 _02933_ _08259_ VGND VGND VPWR VPWR _08303_ sky130_fd_sc_hd__and3_1
X_10285_ _09483_ _00159_ VGND VGND VPWR VPWR _00224_ sky130_fd_sc_hd__xor2_1
X_16901_ _07147_ _07148_ VGND VGND VPWR VPWR _07149_ sky130_fd_sc_hd__xor2_1
X_12024_ _01880_ _01888_ VGND VGND VPWR VPWR _01963_ sky130_fd_sc_hd__or2b_1
X_17881_ _08178_ _08226_ VGND VGND VPWR VPWR _08227_ sky130_fd_sc_hd__nor2_1
X_16832_ _07068_ _07072_ VGND VGND VPWR VPWR _07073_ sky130_fd_sc_hd__xnor2_1
X_16763_ _06994_ _06996_ VGND VGND VPWR VPWR _06998_ sky130_fd_sc_hd__or2b_1
X_13975_ _03945_ _03946_ VGND VGND VPWR VPWR _03947_ sky130_fd_sc_hd__nor2_1
X_18502_ _08851_ _08907_ _08909_ _08833_ VGND VGND VPWR VPWR _08910_ sky130_fd_sc_hd__a22o_1
X_15714_ net478 net179 _05801_ _05802_ VGND VGND VPWR VPWR _05844_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12926_ _02835_ _02863_ _02864_ VGND VGND VPWR VPWR _02865_ sky130_fd_sc_hd__nand3_1
X_16694_ _06907_ _06919_ _06921_ VGND VGND VPWR VPWR _06922_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_85_Left_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18433_ _06159_ _06162_ _06135_ VGND VGND VPWR VPWR _08835_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15645_ _05755_ _05744_ _05752_ VGND VGND VPWR VPWR _05768_ sky130_fd_sc_hd__nand3_1
X_12857_ net235 _01853_ VGND VGND VPWR VPWR _02796_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18364_ _08754_ _08755_ _08758_ VGND VGND VPWR VPWR _08759_ sky130_fd_sc_hd__a21oi_1
X_11808_ _05754_ prev_error\[14\] VGND VGND VPWR VPWR _01747_ sky130_fd_sc_hd__and2b_1
X_15576_ _05684_ _05680_ _05682_ VGND VGND VPWR VPWR _05692_ sky130_fd_sc_hd__or3_1
X_12788_ _02724_ _02725_ _02726_ VGND VGND VPWR VPWR _02727_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17315_ _07300_ _07298_ _07299_ VGND VGND VPWR VPWR _07605_ sky130_fd_sc_hd__nand3_1
XFILLER_0_126_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14527_ _04452_ _04537_ VGND VGND VPWR VPWR _04538_ sky130_fd_sc_hd__nor2_1
X_11739_ _01212_ _01278_ VGND VGND VPWR VPWR _01678_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18295_ i_error\[16\] _08525_ VGND VGND VPWR VPWR _08683_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17246_ _07526_ _07527_ net311 _06437_ VGND VGND VPWR VPWR _07529_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_142_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14458_ _04442_ _04461_ _04459_ VGND VGND VPWR VPWR _04462_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13409_ _03362_ _03364_ VGND VGND VPWR VPWR _03365_ sky130_fd_sc_hd__nor2_1
X_17177_ _07451_ _07452_ VGND VGND VPWR VPWR _07453_ sky130_fd_sc_hd__nor2_1
X_14389_ net451 net456 net128 net125 VGND VGND VPWR VPWR _04386_ sky130_fd_sc_hd__and4_1
XFILLER_0_4_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_94_Left_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16128_ _01805_ VGND VGND VPWR VPWR _06299_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16059_ _09098_ _06222_ VGND VGND VPWR VPWR _06223_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_135_Right_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_20 net347 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_31 net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10070_ _06755_ _08108_ VGND VGND VPWR VPWR _08119_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_102_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13760_ net263 _02543_ _03725_ VGND VGND VPWR VPWR _03726_ sky130_fd_sc_hd__and3_1
X_10972_ net343 _00811_ VGND VGND VPWR VPWR _00911_ sky130_fd_sc_hd__nand2_1
X_12711_ _02647_ _02649_ VGND VGND VPWR VPWR _02650_ sky130_fd_sc_hd__or2b_1
X_13691_ _03650_ _03654_ _03594_ _03655_ VGND VGND VPWR VPWR _03656_ sky130_fd_sc_hd__o211ai_2
Xmax_cap99 net536 VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12642_ _02493_ _02492_ VGND VGND VPWR VPWR _02581_ sky130_fd_sc_hd__and2b_1
X_15430_ _05429_ _05519_ _05521_ VGND VGND VPWR VPWR _05531_ sky130_fd_sc_hd__or3_1
XFILLER_0_66_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15361_ _05449_ _05454_ VGND VGND VPWR VPWR _05455_ sky130_fd_sc_hd__or2b_1
X_12573_ _02511_ VGND VGND VPWR VPWR _02512_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17100_ _07334_ _07342_ _07367_ VGND VGND VPWR VPWR _07368_ sky130_fd_sc_hd__a21o_1
X_14312_ _04158_ _04298_ _04297_ VGND VGND VPWR VPWR _04301_ sky130_fd_sc_hd__a21o_1
X_11524_ net385 _00798_ VGND VGND VPWR VPWR _01463_ sky130_fd_sc_hd__nand2_1
X_15292_ _04016_ net197 _05378_ VGND VGND VPWR VPWR _05379_ sky130_fd_sc_hd__nor3_1
XFILLER_0_124_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18080_ _07786_ _07787_ _07790_ VGND VGND VPWR VPWR _08446_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_80_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14243_ _04223_ _04224_ VGND VGND VPWR VPWR _04226_ sky130_fd_sc_hd__and2_1
X_17031_ net315 _06352_ VGND VGND VPWR VPWR _07292_ sky130_fd_sc_hd__nand2_1
X_11455_ _01308_ _01307_ VGND VGND VPWR VPWR _01394_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10406_ _00318_ _00343_ VGND VGND VPWR VPWR _00345_ sky130_fd_sc_hd__nand2_1
X_14174_ _04147_ _04149_ VGND VGND VPWR VPWR _04150_ sky130_fd_sc_hd__nand2_1
X_11386_ net382 _01324_ _01285_ _00244_ VGND VGND VPWR VPWR _01325_ sky130_fd_sc_hd__and4_1
XFILLER_0_104_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13125_ _03055_ _03068_ _03071_ VGND VGND VPWR VPWR _03072_ sky130_fd_sc_hd__o21ba_1
X_10337_ _00274_ _00275_ VGND VGND VPWR VPWR _00276_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18982_ _09360_ _09437_ VGND VGND VPWR VPWR _09438_ sky130_fd_sc_hd__xnor2_4
X_13056_ _02952_ _02995_ VGND VGND VPWR VPWR _02996_ sky130_fd_sc_hd__or2_1
X_17933_ _07570_ _08277_ VGND VGND VPWR VPWR _08285_ sky130_fd_sc_hd__nand2_1
X_10268_ net360 _06073_ VGND VGND VPWR VPWR _00207_ sky130_fd_sc_hd__nand2_1
X_12007_ _01938_ _01944_ VGND VGND VPWR VPWR _01946_ sky130_fd_sc_hd__and2_1
X_17864_ _08018_ _08208_ _08125_ VGND VGND VPWR VPWR _08209_ sky130_fd_sc_hd__a21o_1
X_10199_ net350 _06194_ _09514_ VGND VGND VPWR VPWR _09521_ sky130_fd_sc_hd__and3_1
X_16815_ _07051_ _07054_ VGND VGND VPWR VPWR _07055_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17795_ _08117_ _08118_ _08132_ VGND VGND VPWR VPWR _08133_ sky130_fd_sc_hd__nor3_1
X_16746_ _06888_ _06894_ _06895_ VGND VGND VPWR VPWR _06979_ sky130_fd_sc_hd__or3_2
X_13958_ _03926_ _03929_ VGND VGND VPWR VPWR _03930_ sky130_fd_sc_hd__xor2_1
X_12909_ _02846_ _02847_ VGND VGND VPWR VPWR _02848_ sky130_fd_sc_hd__xnor2_1
X_16677_ _06899_ _06902_ VGND VGND VPWR VPWR _06903_ sky130_fd_sc_hd__nor2_1
X_13889_ _03425_ _03854_ VGND VGND VPWR VPWR _03855_ sky130_fd_sc_hd__or2b_1
XFILLER_0_146_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18416_ _06154_ _06157_ VGND VGND VPWR VPWR _08816_ sky130_fd_sc_hd__nor2_1
X_15628_ _05747_ _05748_ VGND VGND VPWR VPWR _05749_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18347_ _06133_ _08616_ VGND VGND VPWR VPWR _08740_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15559_ _05548_ _05672_ VGND VGND VPWR VPWR _05673_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18278_ _06567_ _08655_ _08662_ VGND VGND VPWR VPWR _08664_ sky130_fd_sc_hd__or3_1
XFILLER_0_71_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput40 reg_data[0] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_4
X_17229_ _07508_ _07509_ VGND VGND VPWR VPWR _07510_ sky130_fd_sc_hd__xor2_1
XFILLER_0_31_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput51 reg_data[2] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput62 target[11] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput73 target[4] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_1
XFILLER_0_3_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09982_ _06282_ _06381_ _06359_ VGND VGND VPWR VPWR _07151_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_58_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11240_ _04621_ _06579_ _04533_ VGND VGND VPWR VPWR _01179_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_132_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11171_ net346 _00812_ _01109_ _01107_ VGND VGND VPWR VPWR _01110_ sky130_fd_sc_hd__a31o_1
X_10122_ _08669_ _08680_ VGND VGND VPWR VPWR _08691_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10053_ _07844_ _07910_ VGND VGND VPWR VPWR _07932_ sky130_fd_sc_hd__xnor2_1
X_14930_ _04912_ _04926_ _04920_ _04925_ VGND VGND VPWR VPWR _04981_ sky130_fd_sc_hd__a211o_1
X_14861_ net454 net459 net154 net148 VGND VGND VPWR VPWR _04905_ sky130_fd_sc_hd__and4_1
XFILLER_0_54_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16600_ _06806_ _06816_ _06817_ VGND VGND VPWR VPWR _06818_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13812_ _03738_ _03743_ _03742_ VGND VGND VPWR VPWR _03778_ sky130_fd_sc_hd__a21oi_1
X_17580_ net332 _06400_ _07895_ VGND VGND VPWR VPWR _07896_ sky130_fd_sc_hd__a21oi_1
X_14792_ net449 net155 _04517_ VGND VGND VPWR VPWR _04829_ sky130_fd_sc_hd__and3_1
X_16531_ _06740_ _06739_ VGND VGND VPWR VPWR _06742_ sky130_fd_sc_hd__xor2_1
X_13743_ _03707_ _03708_ VGND VGND VPWR VPWR _03709_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10955_ _00877_ _00882_ _00883_ VGND VGND VPWR VPWR _00894_ sky130_fd_sc_hd__nor3_1
XFILLER_0_85_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19250_ clknet_4_13_0_clock _00132_ VGND VGND VPWR VPWR i_error\[18\] sky130_fd_sc_hd__dfxtp_1
X_16462_ _06646_ _06664_ _06665_ VGND VGND VPWR VPWR _06666_ sky130_fd_sc_hd__a21oi_1
X_13674_ net256 _02407_ _03637_ VGND VGND VPWR VPWR _03638_ sky130_fd_sc_hd__and3_1
X_10886_ _00824_ _00823_ VGND VGND VPWR VPWR _00825_ sky130_fd_sc_hd__xnor2_1
X_18201_ _08544_ _08571_ _08576_ _08577_ _08578_ VGND VGND VPWR VPWR _08579_ sky130_fd_sc_hd__o311a_4
X_15413_ _05510_ _05506_ _05508_ VGND VGND VPWR VPWR _05513_ sky130_fd_sc_hd__or3_1
XFILLER_0_156_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12625_ _02558_ _02532_ VGND VGND VPWR VPWR _02564_ sky130_fd_sc_hd__or2b_1
X_19181_ _09550_ _09013_ _09587_ net490 VGND VGND VPWR VPWR _00145_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16393_ _06368_ _06379_ _06366_ VGND VGND VPWR VPWR _06591_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_54_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18132_ _07084_ _07113_ VGND VGND VPWR VPWR _08503_ sky130_fd_sc_hd__nand2_1
X_12556_ _02491_ _02494_ VGND VGND VPWR VPWR _02495_ sky130_fd_sc_hd__nand2_1
X_15344_ _05345_ _05349_ VGND VGND VPWR VPWR _05437_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11507_ _01371_ _01383_ VGND VGND VPWR VPWR _01446_ sky130_fd_sc_hd__xnor2_1
X_18063_ _08158_ _08162_ VGND VGND VPWR VPWR _08428_ sky130_fd_sc_hd__and2_1
X_12487_ _02425_ VGND VGND VPWR VPWR _02426_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15275_ _05239_ _05302_ _05334_ _05360_ VGND VGND VPWR VPWR _05361_ sky130_fd_sc_hd__a31oi_1
X_17014_ _07248_ _07271_ _07273_ VGND VGND VPWR VPWR _07274_ sky130_fd_sc_hd__o21ba_1
X_14226_ _04186_ _04187_ _04205_ VGND VGND VPWR VPWR _04207_ sky130_fd_sc_hd__o21ai_1
X_11438_ net395 _09558_ _09565_ _01376_ VGND VGND VPWR VPWR _01377_ sky130_fd_sc_hd__nand4_2
XFILLER_0_110_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14157_ net428 net433 net117 VGND VGND VPWR VPWR _04131_ sky130_fd_sc_hd__and3_1
X_11369_ _01303_ _01306_ _01302_ VGND VGND VPWR VPWR _01308_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13108_ _03051_ _03052_ VGND VGND VPWR VPWR _03053_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14088_ _04058_ _04029_ _04032_ VGND VGND VPWR VPWR _04060_ sky130_fd_sc_hd__and3_1
X_18965_ _03916_ _09258_ _03920_ VGND VGND VPWR VPWR _09420_ sky130_fd_sc_hd__o21ba_1
X_13039_ _02865_ _02876_ _02974_ VGND VGND VPWR VPWR _02978_ sky130_fd_sc_hd__a21o_1
X_17916_ net318 _07181_ VGND VGND VPWR VPWR _08266_ sky130_fd_sc_hd__nand2_1
X_18896_ _03891_ _06006_ _06127_ VGND VGND VPWR VPWR _09344_ sky130_fd_sc_hd__o21ba_2
X_17847_ net301 _07568_ VGND VGND VPWR VPWR _08190_ sky130_fd_sc_hd__nand2_1
X_17778_ _08106_ _08113_ VGND VGND VPWR VPWR _08114_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16729_ net299 _06401_ VGND VGND VPWR VPWR _06960_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09965_ _06876_ _06953_ VGND VGND VPWR VPWR _06964_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_31_Left_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09896_ net341 _06007_ _06073_ net344 VGND VGND VPWR VPWR _06205_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_79_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10740_ _00668_ _00671_ VGND VGND VPWR VPWR _00679_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_40_Left_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10671_ _00608_ _00609_ VGND VGND VPWR VPWR _00610_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12410_ _02347_ _02348_ VGND VGND VPWR VPWR _02349_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13390_ _03342_ _03343_ VGND VGND VPWR VPWR _03344_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12341_ _02264_ _02268_ _02262_ VGND VGND VPWR VPWR _02280_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_106_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15060_ _05114_ _05118_ _05115_ VGND VGND VPWR VPWR _05124_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_121_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12272_ _02084_ _02095_ _02096_ VGND VGND VPWR VPWR _02211_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14011_ _03970_ _03977_ _03982_ VGND VGND VPWR VPWR _03983_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11223_ _01161_ _01109_ VGND VGND VPWR VPWR _01162_ sky130_fd_sc_hd__xnor2_2
X_11154_ _01091_ _01092_ VGND VGND VPWR VPWR _01093_ sky130_fd_sc_hd__nand2_1
X_10105_ _07734_ _08493_ VGND VGND VPWR VPWR _08504_ sky130_fd_sc_hd__or2_2
X_18750_ _09181_ _09182_ VGND VGND VPWR VPWR _09183_ sky130_fd_sc_hd__xnor2_4
X_15962_ _06041_ _06114_ _06115_ VGND VGND VPWR VPWR _06116_ sky130_fd_sc_hd__a21o_2
X_11085_ net565 _00613_ VGND VGND VPWR VPWR _01024_ sky130_fd_sc_hd__nand2_1
X_17701_ _08026_ _08007_ _08027_ VGND VGND VPWR VPWR _08029_ sky130_fd_sc_hd__and3_1
X_10036_ _07613_ _07679_ VGND VGND VPWR VPWR _07745_ sky130_fd_sc_hd__xor2_1
X_14913_ net473 VGND VGND VPWR VPWR _04963_ sky130_fd_sc_hd__inv_2
X_18681_ _09101_ _09103_ _09102_ VGND VGND VPWR VPWR _09107_ sky130_fd_sc_hd__o21ai_1
X_15893_ _06036_ _06039_ VGND VGND VPWR VPWR _06041_ sky130_fd_sc_hd__nand2_1
X_17632_ _07940_ _07947_ VGND VGND VPWR VPWR _07953_ sky130_fd_sc_hd__and2b_1
X_14844_ _04854_ _04883_ _04886_ VGND VGND VPWR VPWR _04887_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17563_ _07875_ _07874_ _07873_ _07868_ VGND VGND VPWR VPWR _07878_ sky130_fd_sc_hd__a211o_1
X_14775_ _04693_ _04695_ VGND VGND VPWR VPWR _04811_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11987_ net242 net238 _01772_ _01771_ VGND VGND VPWR VPWR _01926_ sky130_fd_sc_hd__a31o_1
X_19302_ clknet_4_7_0_clock _00042_ VGND VGND VPWR VPWR ki\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16514_ _06723_ VGND VGND VPWR VPWR _06724_ sky130_fd_sc_hd__clkbuf_4
X_13726_ net237 _02934_ VGND VGND VPWR VPWR _03692_ sky130_fd_sc_hd__nand2_1
X_10938_ _00874_ _00876_ VGND VGND VPWR VPWR _00877_ sky130_fd_sc_hd__and2_1
X_17494_ net332 net514 _06619_ net315 VGND VGND VPWR VPWR _07802_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19233_ clknet_4_9_0_clock _00115_ VGND VGND VPWR VPWR i_error\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16445_ _06616_ _06643_ VGND VGND VPWR VPWR _06648_ sky130_fd_sc_hd__xor2_2
X_13657_ _03617_ _03618_ VGND VGND VPWR VPWR _03619_ sky130_fd_sc_hd__xnor2_1
X_10869_ net2 net60 VGND VGND VPWR VPWR _00808_ sky130_fd_sc_hd__or2b_2
XFILLER_0_156_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12608_ net204 _02410_ VGND VGND VPWR VPWR _02547_ sky130_fd_sc_hd__nand2_1
X_19164_ net501 net468 VGND VGND VPWR VPWR _09578_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16376_ _06560_ _06571_ VGND VGND VPWR VPWR _06572_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13588_ _03541_ _03545_ _03490_ _03524_ VGND VGND VPWR VPWR _03547_ sky130_fd_sc_hd__a211o_1
X_18115_ _07795_ _07768_ VGND VGND VPWR VPWR _08485_ sky130_fd_sc_hd__and2b_1
XFILLER_0_14_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15327_ _05410_ _05416_ _05404_ VGND VGND VPWR VPWR _05418_ sky130_fd_sc_hd__a21o_1
XFILLER_0_81_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12539_ _02476_ _02477_ VGND VGND VPWR VPWR _02478_ sky130_fd_sc_hd__nor2_1
X_19095_ net499 prev_error\[9\] VGND VGND VPWR VPWR _09535_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18046_ _08296_ _08298_ _08297_ VGND VGND VPWR VPWR _08409_ sky130_fd_sc_hd__o21a_1
X_15258_ _05243_ _05242_ VGND VGND VPWR VPWR _05342_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14209_ _04136_ _04138_ _04128_ VGND VGND VPWR VPWR _04188_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_100_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15189_ _05075_ _05178_ VGND VGND VPWR VPWR _05266_ sky130_fd_sc_hd__nor2_1
Xfanout408 net410 VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__buf_2
Xfanout419 prev_d_error\[15\] VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__buf_2
X_09750_ _04577_ _04588_ VGND VGND VPWR VPWR _04599_ sky130_fd_sc_hd__nand2_1
X_18948_ _09388_ _09400_ VGND VGND VPWR VPWR _09401_ sky130_fd_sc_hd__xnor2_1
X_09681_ net21 net33 net32 _03592_ VGND VGND VPWR VPWR _03859_ sky130_fd_sc_hd__or4b_4
XFILLER_0_146_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18879_ _02145_ _02162_ _02160_ VGND VGND VPWR VPWR _09325_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09948_ _06447_ _06766_ VGND VGND VPWR VPWR _06777_ sky130_fd_sc_hd__or2_1
X_09879_ net338 _06007_ VGND VGND VPWR VPWR _06018_ sky130_fd_sc_hd__nand2_1
X_11910_ _01705_ _01736_ VGND VGND VPWR VPWR _01849_ sky130_fd_sc_hd__nand2_4
XFILLER_0_99_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12890_ _02828_ _02740_ VGND VGND VPWR VPWR _02829_ sky130_fd_sc_hd__xnor2_1
X_11841_ _01771_ _01779_ VGND VGND VPWR VPWR _01780_ sky130_fd_sc_hd__nand2_1
X_14560_ _04540_ _04542_ _04545_ VGND VGND VPWR VPWR _04574_ sky130_fd_sc_hd__or3_1
X_11772_ prev_error\[4\] VGND VGND VPWR VPWR _01711_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13511_ net265 _01874_ VGND VGND VPWR VPWR _03470_ sky130_fd_sc_hd__nand2_1
X_10723_ _00656_ _00654_ VGND VGND VPWR VPWR _00662_ sky130_fd_sc_hd__xor2_4
X_14491_ _04490_ _04495_ _04496_ _04497_ VGND VGND VPWR VPWR _04498_ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16230_ net275 _06410_ VGND VGND VPWR VPWR _06411_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13442_ _03399_ _03394_ _03397_ VGND VGND VPWR VPWR _03401_ sky130_fd_sc_hd__nor3_1
X_10654_ _00590_ _00592_ _00588_ VGND VGND VPWR VPWR _00593_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13373_ _03249_ _03324_ _03320_ _03323_ VGND VGND VPWR VPWR _03326_ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16161_ _06334_ VGND VGND VPWR VPWR _06335_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10585_ _00502_ _00522_ VGND VGND VPWR VPWR _00524_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15112_ _05158_ _05162_ _05180_ VGND VGND VPWR VPWR _05181_ sky130_fd_sc_hd__o21a_1
X_12324_ _02259_ _02261_ VGND VGND VPWR VPWR _02263_ sky130_fd_sc_hd__nor2_1
X_16092_ _06250_ _06258_ VGND VGND VPWR VPWR _06259_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_23_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15043_ net471 net476 net149 net143 VGND VGND VPWR VPWR _05106_ sky130_fd_sc_hd__and4_1
X_12255_ net230 net226 _01807_ _01814_ VGND VGND VPWR VPWR _02194_ sky130_fd_sc_hd__and4_1
XFILLER_0_32_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11206_ net374 _00242_ VGND VGND VPWR VPWR _01145_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12186_ _01883_ _01958_ VGND VGND VPWR VPWR _02125_ sky130_fd_sc_hd__nor2_1
X_18802_ _09231_ _09239_ VGND VGND VPWR VPWR _09240_ sky130_fd_sc_hd__xnor2_1
X_11137_ _01073_ _01074_ _01066_ VGND VGND VPWR VPWR _01076_ sky130_fd_sc_hd__a21oi_1
X_16994_ net294 _06802_ VGND VGND VPWR VPWR _07252_ sky130_fd_sc_hd__nand2_1
X_18733_ _09162_ _09163_ VGND VGND VPWR VPWR _09165_ sky130_fd_sc_hd__or2_4
X_15945_ _06075_ _06097_ VGND VGND VPWR VPWR _06098_ sky130_fd_sc_hd__nand2_1
X_11068_ net346 _00615_ _00905_ VGND VGND VPWR VPWR _01007_ sky130_fd_sc_hd__a21oi_1
X_10019_ _07360_ _07415_ _07547_ VGND VGND VPWR VPWR _07558_ sky130_fd_sc_hd__a21oi_1
X_18664_ _06099_ _09088_ VGND VGND VPWR VPWR _09089_ sky130_fd_sc_hd__and2_1
X_15876_ _02466_ _03883_ VGND VGND VPWR VPWR _06022_ sky130_fd_sc_hd__xor2_4
X_17615_ _07933_ _07927_ _07930_ VGND VGND VPWR VPWR _07935_ sky130_fd_sc_hd__nor3_1
XFILLER_0_25_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14827_ _04864_ _04867_ VGND VGND VPWR VPWR _04868_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18595_ _06119_ _09012_ VGND VGND VPWR VPWR _09013_ sky130_fd_sc_hd__and2_2
XFILLER_0_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17546_ _07856_ _07858_ VGND VGND VPWR VPWR _07859_ sky130_fd_sc_hd__nand2_1
X_14758_ _04715_ _04717_ VGND VGND VPWR VPWR _04792_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13709_ _03673_ _03674_ VGND VGND VPWR VPWR _03675_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17477_ _07717_ _07727_ VGND VGND VPWR VPWR _07783_ sky130_fd_sc_hd__and2_1
X_14689_ _04699_ _04688_ _04696_ VGND VGND VPWR VPWR _04716_ sky130_fd_sc_hd__nand3_1
XFILLER_0_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19216_ clknet_4_4_0_clock _00098_ VGND VGND VPWR VPWR prev_error\[3\] sky130_fd_sc_hd__dfxtp_2
X_16428_ net283 _06404_ VGND VGND VPWR VPWR _06629_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19147_ _09559_ _08991_ _09567_ net495 VGND VGND VPWR VPWR _00128_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16359_ _06542_ _06547_ _06552_ VGND VGND VPWR VPWR _06553_ sky130_fd_sc_hd__nor3_1
X_19078_ _09523_ _00812_ _09524_ net487 VGND VGND VPWR VPWR _00095_ sky130_fd_sc_hd__o211a_1
XFILLER_0_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18029_ _08385_ _08389_ VGND VGND VPWR VPWR _08390_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout205 net207 VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout216 kd_1\[13\] VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__buf_2
Xfanout227 kd_1\[10\] VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__clkbuf_4
X_09802_ _05160_ VGND VGND VPWR VPWR _05171_ sky130_fd_sc_hd__buf_8
XFILLER_0_10_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout238 net241 VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__clkbuf_4
Xfanout249 kd_1\[5\] VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_66_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09733_ _04390_ _04401_ VGND VGND VPWR VPWR _04412_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_105_Left_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09664_ net51 _03625_ _03658_ net325 VGND VGND VPWR VPWR _00049_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_114_Left_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_149_Right_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10370_ _00284_ _00308_ VGND VGND VPWR VPWR _00309_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12040_ _01972_ _01978_ VGND VGND VPWR VPWR _01979_ sky130_fd_sc_hd__nor2b_4
XFILLER_0_103_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_123_Left_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13991_ net438 net443 net132 net127 VGND VGND VPWR VPWR _03963_ sky130_fd_sc_hd__and4_1
X_15730_ _05830_ _05858_ VGND VGND VPWR VPWR _05861_ sky130_fd_sc_hd__xnor2_1
X_12942_ net252 _02880_ _01785_ VGND VGND VPWR VPWR _02881_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15661_ _05730_ _05734_ _05784_ VGND VGND VPWR VPWR _05785_ sky130_fd_sc_hd__o21ai_1
X_12873_ _02726_ _02724_ VGND VGND VPWR VPWR _02812_ sky130_fd_sc_hd__or2b_1
X_17400_ _07308_ _07696_ _07695_ VGND VGND VPWR VPWR _07698_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_157_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14612_ _04629_ _04630_ VGND VGND VPWR VPWR _04631_ sky130_fd_sc_hd__nor2_1
X_11824_ net246 VGND VGND VPWR VPWR _01763_ sky130_fd_sc_hd__inv_2
X_18380_ _06141_ _06158_ VGND VGND VPWR VPWR _08776_ sky130_fd_sc_hd__or2b_1
X_15592_ _05697_ _05707_ _05708_ VGND VGND VPWR VPWR _05709_ sky130_fd_sc_hd__nand3_1
XFILLER_0_157_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17331_ net308 _06437_ VGND VGND VPWR VPWR _07622_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14543_ _04553_ _04554_ VGND VGND VPWR VPWR _04556_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11755_ _00464_ _00563_ _01692_ _01693_ _00463_ VGND VGND VPWR VPWR _01694_ sky130_fd_sc_hd__a32o_2
XPHY_EDGE_ROW_132_Left_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17262_ _07532_ _07533_ _07544_ VGND VGND VPWR VPWR _07546_ sky130_fd_sc_hd__o21ai_1
X_10706_ _00633_ _00643_ VGND VGND VPWR VPWR _00645_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14474_ _04476_ _04479_ VGND VGND VPWR VPWR _04480_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11686_ _01623_ _01624_ VGND VGND VPWR VPWR _01625_ sky130_fd_sc_hd__and2b_1
XFILLER_0_153_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19001_ _09165_ _09454_ VGND VGND VPWR VPWR _09459_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_36_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16213_ _06387_ _06391_ VGND VGND VPWR VPWR _06393_ sky130_fd_sc_hd__xnor2_1
X_13425_ _03367_ _03354_ _03365_ VGND VGND VPWR VPWR _03383_ sky130_fd_sc_hd__nor3_1
X_17193_ _07466_ _07467_ _07468_ VGND VGND VPWR VPWR _07471_ sky130_fd_sc_hd__a21o_1
X_10637_ _00574_ _00575_ VGND VGND VPWR VPWR _00576_ sky130_fd_sc_hd__and2b_1
XFILLER_0_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16144_ _06313_ _06307_ _01757_ VGND VGND VPWR VPWR _06317_ sky130_fd_sc_hd__nand3_1
XFILLER_0_134_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13356_ _03307_ _03308_ VGND VGND VPWR VPWR _03309_ sky130_fd_sc_hd__nor2_1
X_10568_ net352 _09583_ _00398_ _00506_ VGND VGND VPWR VPWR _00507_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_116_Right_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12307_ _02209_ _02244_ _02111_ _02245_ VGND VGND VPWR VPWR _02246_ sky130_fd_sc_hd__a211o_1
XFILLER_0_133_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16075_ _05666_ _06204_ _06201_ VGND VGND VPWR VPWR _06241_ sky130_fd_sc_hd__a21o_1
X_13287_ net265 _01859_ _03239_ _03237_ VGND VGND VPWR VPWR _03240_ sky130_fd_sc_hd__a31o_1
X_10499_ net401 _05061_ VGND VGND VPWR VPWR _00438_ sky130_fd_sc_hd__nand2_2
X_15026_ _05078_ _05081_ _05086_ VGND VGND VPWR VPWR _05087_ sky130_fd_sc_hd__o21ai_2
X_12238_ net242 net238 net111 _01786_ VGND VGND VPWR VPWR _02177_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12169_ _02106_ _02102_ VGND VGND VPWR VPWR _02108_ sky130_fd_sc_hd__or2b_1
XFILLER_0_127_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16977_ net299 _06437_ _06467_ net297 VGND VGND VPWR VPWR _07233_ sky130_fd_sc_hd__a22oi_2
Xinput5 measurement[12] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_1
XFILLER_0_36_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15928_ _03853_ _06078_ VGND VGND VPWR VPWR _06079_ sky130_fd_sc_hd__nor2_1
X_18716_ _09144_ _09139_ _09140_ VGND VGND VPWR VPWR _09146_ sky130_fd_sc_hd__nand3_1
X_18647_ _09060_ _09067_ _09069_ VGND VGND VPWR VPWR _09070_ sky130_fd_sc_hd__or3_1
X_15859_ _04300_ _04301_ _05999_ _06002_ VGND VGND VPWR VPWR _06003_ sky130_fd_sc_hd__and4_1
XFILLER_0_148_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18578_ _06133_ _08993_ VGND VGND VPWR VPWR _08994_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17529_ _07488_ _07496_ VGND VGND VPWR VPWR _07840_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09716_ _04203_ _04214_ VGND VGND VPWR VPWR _04225_ sky130_fd_sc_hd__nand2_4
X_09647_ net42 _03347_ _03380_ net223 VGND VGND VPWR VPWR _00002_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11540_ _01476_ _01478_ VGND VGND VPWR VPWR _01479_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11471_ _01350_ _01351_ _01409_ VGND VGND VPWR VPWR _01410_ sky130_fd_sc_hd__a21o_1
XFILLER_0_107_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10422_ _00280_ _00360_ VGND VGND VPWR VPWR _00361_ sky130_fd_sc_hd__xor2_2
X_13210_ _03122_ _03162_ VGND VGND VPWR VPWR _03163_ sky130_fd_sc_hd__nor2_1
X_14190_ _04165_ net134 net408 _04166_ VGND VGND VPWR VPWR _04167_ sky130_fd_sc_hd__and4b_1
XFILLER_0_104_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13141_ _03086_ _03088_ VGND VGND VPWR VPWR _03089_ sky130_fd_sc_hd__or2_1
X_10353_ net364 _06062_ _00209_ VGND VGND VPWR VPWR _00292_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13072_ net239 _01908_ _01874_ net244 VGND VGND VPWR VPWR _03013_ sky130_fd_sc_hd__a22o_1
X_10284_ _00201_ _00203_ _00222_ VGND VGND VPWR VPWR _00223_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_57_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16900_ _07006_ _07034_ VGND VGND VPWR VPWR _07148_ sky130_fd_sc_hd__xnor2_1
X_12023_ _01955_ _01961_ VGND VGND VPWR VPWR _01962_ sky130_fd_sc_hd__xor2_1
X_17880_ net322 _07155_ VGND VGND VPWR VPWR _08226_ sky130_fd_sc_hd__nand2_1
X_16831_ net299 _06402_ _07069_ _07071_ VGND VGND VPWR VPWR _07072_ sky130_fd_sc_hd__a31oi_2
X_16762_ _06990_ _06995_ VGND VGND VPWR VPWR _06996_ sky130_fd_sc_hd__and2_1
X_13974_ net426 net128 net126 net567 VGND VGND VPWR VPWR _03946_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_88_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18501_ _08908_ VGND VGND VPWR VPWR _08909_ sky130_fd_sc_hd__inv_2
X_15713_ _05839_ _05841_ VGND VGND VPWR VPWR _05843_ sky130_fd_sc_hd__nor2_1
X_12925_ _02730_ _02834_ _02809_ _02833_ VGND VGND VPWR VPWR _02864_ sky130_fd_sc_hd__a211o_1
X_16693_ _06908_ _06918_ VGND VGND VPWR VPWR _06921_ sky130_fd_sc_hd__nor2_1
X_18432_ _08595_ _08832_ VGND VGND VPWR VPWR _08833_ sky130_fd_sc_hd__xnor2_2
X_15644_ _05764_ _05766_ VGND VGND VPWR VPWR _05767_ sky130_fd_sc_hd__nor2_1
X_12856_ _02779_ _02780_ _02794_ VGND VGND VPWR VPWR _02795_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_146_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18363_ _08756_ _08620_ VGND VGND VPWR VPWR _08758_ sky130_fd_sc_hd__nand2_1
X_11807_ prev_error\[14\] _05754_ VGND VGND VPWR VPWR _01746_ sky130_fd_sc_hd__or2b_1
XFILLER_0_28_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15575_ _05689_ _05690_ VGND VGND VPWR VPWR _05691_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12787_ _02720_ _02723_ VGND VGND VPWR VPWR _02726_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17314_ _07523_ _07530_ VGND VGND VPWR VPWR _07604_ sky130_fd_sc_hd__nand2_1
X_14526_ net409 net175 _04450_ _04451_ VGND VGND VPWR VPWR _04537_ sky130_fd_sc_hd__o2bb2a_1
X_11738_ _01410_ _01675_ _01676_ VGND VGND VPWR VPWR _01677_ sky130_fd_sc_hd__a21oi_2
X_18294_ i_error\[17\] _08681_ VGND VGND VPWR VPWR _08682_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17245_ _06544_ _06452_ _07526_ _07527_ VGND VGND VPWR VPWR _07528_ sky130_fd_sc_hd__or4_4
X_14457_ _04459_ _04460_ VGND VGND VPWR VPWR _04461_ sky130_fd_sc_hd__nor2_1
X_11669_ _01592_ _01607_ VGND VGND VPWR VPWR _01608_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13408_ _03354_ _03363_ VGND VGND VPWR VPWR _03364_ sky130_fd_sc_hd__or2_1
X_17176_ _07447_ _07449_ _07450_ VGND VGND VPWR VPWR _07452_ sky130_fd_sc_hd__and3_1
X_14388_ _03955_ _04316_ VGND VGND VPWR VPWR _04385_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16127_ _01706_ VGND VGND VPWR VPWR _06298_ sky130_fd_sc_hd__inv_2
X_13339_ _03289_ _03290_ _03291_ VGND VGND VPWR VPWR _03292_ sky130_fd_sc_hd__o21ba_1
X_16058_ _06220_ _06221_ VGND VGND VPWR VPWR _06222_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15009_ net427 net432 net184 net181 VGND VGND VPWR VPWR _05068_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_10 ki\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_21 net355 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_32 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10971_ _00902_ _00906_ _00909_ VGND VGND VPWR VPWR _00910_ sky130_fd_sc_hd__o21ai_1
X_12710_ _02646_ _02648_ VGND VGND VPWR VPWR _02649_ sky130_fd_sc_hd__and2_1
X_13690_ _03589_ _03593_ _03591_ VGND VGND VPWR VPWR _03655_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12641_ _02577_ _02578_ _02579_ VGND VGND VPWR VPWR _02580_ sky130_fd_sc_hd__o21ba_1
X_15360_ _05452_ _05453_ VGND VGND VPWR VPWR _05454_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12572_ _02506_ _02510_ VGND VGND VPWR VPWR _02511_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14311_ _04299_ VGND VGND VPWR VPWR _04300_ sky130_fd_sc_hd__inv_2
X_11523_ _00871_ _06579_ _08163_ VGND VGND VPWR VPWR _01462_ sky130_fd_sc_hd__or3_1
X_15291_ _05299_ _05377_ VGND VGND VPWR VPWR _05378_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17030_ net332 VGND VGND VPWR VPWR _07291_ sky130_fd_sc_hd__inv_2
X_14242_ _03896_ _04222_ VGND VGND VPWR VPWR _04224_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11454_ _01364_ _01368_ _01392_ VGND VGND VPWR VPWR _01393_ sky130_fd_sc_hd__a21bo_1
X_10405_ _00318_ _00343_ VGND VGND VPWR VPWR _00344_ sky130_fd_sc_hd__or2_1
X_14173_ _03916_ _04146_ _04088_ VGND VGND VPWR VPWR _04149_ sky130_fd_sc_hd__or3_1
X_11385_ net386 _01286_ _05963_ _05974_ VGND VGND VPWR VPWR _01324_ sky130_fd_sc_hd__nand4_1
XFILLER_0_0_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13124_ net202 _02915_ _03070_ VGND VGND VPWR VPWR _03071_ sky130_fd_sc_hd__and3_1
X_10336_ _00192_ _00191_ VGND VGND VPWR VPWR _00275_ sky130_fd_sc_hd__or2b_1
X_18981_ _09365_ _09436_ VGND VGND VPWR VPWR _09437_ sky130_fd_sc_hd__xnor2_2
X_10267_ _00205_ _09318_ VGND VGND VPWR VPWR _00206_ sky130_fd_sc_hd__xor2_1
X_13055_ net264 _01813_ _02951_ VGND VGND VPWR VPWR _02995_ sky130_fd_sc_hd__a21oi_1
X_17932_ _08272_ _08281_ _08282_ VGND VGND VPWR VPWR _08283_ sky130_fd_sc_hd__o21a_1
X_12006_ _01938_ _01944_ VGND VGND VPWR VPWR _01945_ sky130_fd_sc_hd__nor2_1
X_17863_ net295 _02933_ VGND VGND VPWR VPWR _08208_ sky130_fd_sc_hd__nand2_1
X_10198_ _09499_ _09507_ VGND VGND VPWR VPWR _09514_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16814_ _07053_ _06949_ VGND VGND VPWR VPWR _07054_ sky130_fd_sc_hd__xnor2_1
X_17794_ _08129_ _08131_ VGND VGND VPWR VPWR _08132_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16745_ _06974_ _06977_ VGND VGND VPWR VPWR _06978_ sky130_fd_sc_hd__xnor2_1
X_13957_ net434 net128 _03927_ _03928_ VGND VGND VPWR VPWR _03929_ sky130_fd_sc_hd__a31o_1
X_12908_ _02751_ _02749_ VGND VGND VPWR VPWR _02847_ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16676_ net270 _06900_ _06901_ VGND VGND VPWR VPWR _06902_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13888_ _03427_ _03499_ _03853_ VGND VGND VPWR VPWR _03854_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_57_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15627_ net462 net187 VGND VGND VPWR VPWR _05748_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18415_ _08808_ _08743_ VGND VGND VPWR VPWR _08815_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12839_ net250 _01806_ VGND VGND VPWR VPWR _02778_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18346_ _08737_ net534 VGND VGND VPWR VPWR _08739_ sky130_fd_sc_hd__nor2_2
X_15558_ _05669_ _05671_ VGND VGND VPWR VPWR _05672_ sky130_fd_sc_hd__or2_1
XFILLER_0_139_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14509_ net439 net147 _04517_ VGND VGND VPWR VPWR _04518_ sky130_fd_sc_hd__and3_1
XFILLER_0_142_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18277_ _06567_ _08655_ _08662_ VGND VGND VPWR VPWR _08663_ sky130_fd_sc_hd__o21ai_1
X_15489_ net442 net447 net196 net192 VGND VGND VPWR VPWR _05596_ sky130_fd_sc_hd__and4_1
X_17228_ net302 _06802_ VGND VGND VPWR VPWR _07509_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput30 reg_addr[18] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
Xinput41 reg_data[10] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput52 reg_data[3] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_4
XFILLER_0_24_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput63 target[12] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_1
XFILLER_0_52_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17159_ _07117_ _07141_ VGND VGND VPWR VPWR _07433_ sky130_fd_sc_hd__xor2_1
XFILLER_0_142_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput74 target[5] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_141_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09981_ _07019_ _07129_ VGND VGND VPWR VPWR _07140_ sky130_fd_sc_hd__xor2_1
XFILLER_0_149_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11170_ _01107_ _01108_ VGND VGND VPWR VPWR _01109_ sky130_fd_sc_hd__nor2_1
X_10121_ _08548_ _08658_ VGND VGND VPWR VPWR _08680_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10052_ _07844_ _07910_ VGND VGND VPWR VPWR _07921_ sky130_fd_sc_hd__or2_1
X_14860_ net454 net154 net148 net459 VGND VGND VPWR VPWR _04904_ sky130_fd_sc_hd__a22oi_2
X_13811_ _03776_ VGND VGND VPWR VPWR _03777_ sky130_fd_sc_hd__inv_2
X_14791_ _04718_ _04792_ _04827_ VGND VGND VPWR VPWR _04828_ sky130_fd_sc_hd__and3_1
X_16530_ _06739_ _06740_ VGND VGND VPWR VPWR _06741_ sky130_fd_sc_hd__and2b_1
X_13742_ _03706_ _03695_ _03699_ VGND VGND VPWR VPWR _03708_ sky130_fd_sc_hd__nand3_1
X_10954_ _00802_ _00891_ _00892_ _00886_ _00890_ VGND VGND VPWR VPWR _00893_ sky130_fd_sc_hd__o32a_1
XFILLER_0_39_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16461_ _06647_ _06663_ VGND VGND VPWR VPWR _06665_ sky130_fd_sc_hd__nor2_1
X_13673_ net260 _02543_ VGND VGND VPWR VPWR _03637_ sky130_fd_sc_hd__and2_1
X_10885_ _00716_ _00797_ VGND VGND VPWR VPWR _00824_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18200_ _08540_ _08541_ i_error\[7\] VGND VGND VPWR VPWR _08578_ sky130_fd_sc_hd__or3b_4
X_15412_ _05506_ _05508_ _05510_ VGND VGND VPWR VPWR _05511_ sky130_fd_sc_hd__o21ai_2
X_12624_ _02471_ _02562_ VGND VGND VPWR VPWR _02563_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19180_ net502 net567 VGND VGND VPWR VPWR _09587_ sky130_fd_sc_hd__or2_1
X_16392_ _06487_ _06588_ VGND VGND VPWR VPWR _06589_ sky130_fd_sc_hd__xor2_1
X_18131_ _07454_ _07457_ VGND VGND VPWR VPWR _08502_ sky130_fd_sc_hd__or2_4
XFILLER_0_26_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15343_ _05400_ _05396_ VGND VGND VPWR VPWR _05436_ sky130_fd_sc_hd__or2b_1
XFILLER_0_136_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12555_ _02430_ _02492_ _02493_ VGND VGND VPWR VPWR _02494_ sky130_fd_sc_hd__a21o_1
XFILLER_0_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18062_ _08316_ _08424_ _08425_ VGND VGND VPWR VPWR _08426_ sky130_fd_sc_hd__or3_1
X_11506_ _01443_ _01444_ VGND VGND VPWR VPWR _01445_ sky130_fd_sc_hd__nor2_1
X_15274_ _05337_ _05357_ _05359_ VGND VGND VPWR VPWR _05360_ sky130_fd_sc_hd__and3_1
X_12486_ _02424_ _02363_ VGND VGND VPWR VPWR _02425_ sky130_fd_sc_hd__xor2_1
XFILLER_0_151_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17013_ _07260_ _07270_ _07251_ VGND VGND VPWR VPWR _07273_ sky130_fd_sc_hd__a21oi_1
X_14225_ _04186_ _04187_ _04205_ VGND VGND VPWR VPWR _04206_ sky130_fd_sc_hd__or3_1
XFILLER_0_124_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11437_ net391 _09552_ _04478_ _00241_ VGND VGND VPWR VPWR _01376_ sky130_fd_sc_hd__and4_1
X_14156_ net428 net119 net118 net433 VGND VGND VPWR VPWR _04130_ sky130_fd_sc_hd__a22oi_1
X_11368_ _01302_ _01303_ _01306_ VGND VGND VPWR VPWR _01307_ sky130_fd_sc_hd__nor3_1
X_13107_ _03040_ _03043_ _03050_ VGND VGND VPWR VPWR _03052_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10319_ _00188_ _00221_ _00257_ VGND VGND VPWR VPWR _00258_ sky130_fd_sc_hd__o21ba_1
X_14087_ _04029_ _04032_ _04058_ VGND VGND VPWR VPWR _04059_ sky130_fd_sc_hd__a21oi_2
X_18964_ _09410_ _09418_ VGND VGND VPWR VPWR _09419_ sky130_fd_sc_hd__xnor2_1
X_11299_ net351 _00811_ _00818_ net565 VGND VGND VPWR VPWR _01238_ sky130_fd_sc_hd__a22o_1
X_13038_ _02910_ _02976_ VGND VGND VPWR VPWR _02977_ sky130_fd_sc_hd__nand2_1
X_17915_ _08263_ _08264_ VGND VGND VPWR VPWR _08265_ sky130_fd_sc_hd__nand2_1
X_18895_ _09341_ _09342_ VGND VGND VPWR VPWR _09343_ sky130_fd_sc_hd__nand2_4
XFILLER_0_28_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17846_ _07895_ _08188_ _08171_ _08172_ VGND VGND VPWR VPWR _08189_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_0_89_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14989_ _04932_ VGND VGND VPWR VPWR _05046_ sky130_fd_sc_hd__inv_2
X_17777_ _08109_ _08112_ VGND VGND VPWR VPWR _08113_ sky130_fd_sc_hd__xor2_1
XFILLER_0_77_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16728_ _06958_ _06864_ VGND VGND VPWR VPWR _06959_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16659_ net286 _06470_ _06807_ _06882_ VGND VGND VPWR VPWR _06883_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18329_ _08653_ _08667_ VGND VGND VPWR VPWR _08720_ sky130_fd_sc_hd__and2b_1
XFILLER_0_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09964_ _06920_ _06942_ VGND VGND VPWR VPWR _06953_ sky130_fd_sc_hd__nand2_1
X_09895_ _06183_ VGND VGND VPWR VPWR _06194_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10670_ _00519_ _00518_ _00517_ VGND VGND VPWR VPWR _00609_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12340_ _02257_ _02278_ VGND VGND VPWR VPWR _02279_ sky130_fd_sc_hd__or2_2
XFILLER_0_35_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12271_ _02089_ VGND VGND VPWR VPWR _02210_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14010_ _03980_ _03981_ VGND VGND VPWR VPWR _03982_ sky130_fd_sc_hd__and2_1
X_11222_ net346 _00811_ VGND VGND VPWR VPWR _01161_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11153_ net363 _00798_ _01001_ net367 VGND VGND VPWR VPWR _01092_ sky130_fd_sc_hd__a22o_1
X_10104_ _07756_ _08438_ _08482_ VGND VGND VPWR VPWR _08493_ sky130_fd_sc_hd__o21a_1
X_15961_ _06031_ _06033_ VGND VGND VPWR VPWR _06115_ sky130_fd_sc_hd__xnor2_1
X_11084_ _01021_ _01022_ VGND VGND VPWR VPWR _01023_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10035_ _06788_ _07723_ VGND VGND VPWR VPWR _07734_ sky130_fd_sc_hd__xnor2_2
X_14912_ net134 VGND VGND VPWR VPWR _04961_ sky130_fd_sc_hd__inv_2
X_17700_ _08026_ _08007_ _08027_ VGND VGND VPWR VPWR _08028_ sky130_fd_sc_hd__a21oi_2
X_15892_ _05982_ _06038_ VGND VGND VPWR VPWR _06039_ sky130_fd_sc_hd__and2b_1
X_18680_ _09093_ _09105_ VGND VGND VPWR VPWR _09106_ sky130_fd_sc_hd__or2_4
X_14843_ _04777_ _04884_ VGND VGND VPWR VPWR _04886_ sky130_fd_sc_hd__nor2_1
X_17631_ _07923_ _07949_ _07950_ _07951_ VGND VGND VPWR VPWR _07952_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_59_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17562_ _07868_ _07873_ _07874_ _07875_ VGND VGND VPWR VPWR _07876_ sky130_fd_sc_hd__o211ai_2
X_14774_ _04807_ _04809_ VGND VGND VPWR VPWR _04810_ sky130_fd_sc_hd__nand2_1
X_11986_ _01894_ _01924_ VGND VGND VPWR VPWR _01925_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19301_ clknet_4_7_0_clock _00041_ VGND VGND VPWR VPWR ki\[12\] sky130_fd_sc_hd__dfxtp_1
X_16513_ _06721_ VGND VGND VPWR VPWR _06723_ sky130_fd_sc_hd__clkbuf_4
X_13725_ _03431_ _03680_ _03682_ _03683_ VGND VGND VPWR VPWR _03691_ sky130_fd_sc_hd__o22ai_1
X_17493_ _07760_ _07762_ _07687_ _07761_ VGND VGND VPWR VPWR _07801_ sky130_fd_sc_hd__a211o_1
X_10937_ _00769_ _00875_ VGND VGND VPWR VPWR _00876_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19232_ clknet_4_9_0_clock _00114_ VGND VGND VPWR VPWR i_error\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16444_ _06580_ _06586_ VGND VGND VPWR VPWR _06647_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_128_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13656_ _03568_ _03567_ VGND VGND VPWR VPWR _03618_ sky130_fd_sc_hd__and2b_1
XFILLER_0_73_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10868_ _00803_ _00806_ VGND VGND VPWR VPWR _00807_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_144_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12607_ _02545_ VGND VGND VPWR VPWR _02546_ sky130_fd_sc_hd__clkbuf_4
X_19163_ _09559_ _09089_ _09576_ net490 VGND VGND VPWR VPWR _00136_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16375_ _06376_ _06570_ VGND VGND VPWR VPWR _06571_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13587_ _03490_ _03524_ _03541_ _03545_ VGND VGND VPWR VPWR _03546_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_30_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10799_ _00731_ _00737_ VGND VGND VPWR VPWR _00738_ sky130_fd_sc_hd__nand2_1
X_18114_ _07797_ _07764_ VGND VGND VPWR VPWR _08484_ sky130_fd_sc_hd__and2b_1
X_15326_ _05404_ _05410_ _05416_ VGND VGND VPWR VPWR _05417_ sky130_fd_sc_hd__nand3_1
X_12538_ _02364_ _01786_ VGND VGND VPWR VPWR _02477_ sky130_fd_sc_hd__and2_1
X_19094_ _09523_ _08207_ _09534_ net488 VGND VGND VPWR VPWR _00103_ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18045_ _08345_ _08346_ _08323_ VGND VGND VPWR VPWR _08408_ sky130_fd_sc_hd__or3b_1
X_15257_ _05338_ _05339_ _05340_ VGND VGND VPWR VPWR _05341_ sky130_fd_sc_hd__o21ba_1
X_12469_ _02407_ VGND VGND VPWR VPWR _02408_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_151_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14208_ _04118_ _04162_ _04185_ VGND VGND VPWR VPWR _04187_ sky130_fd_sc_hd__and3_1
X_15188_ _05165_ _05206_ _05264_ VGND VGND VPWR VPWR _05265_ sky130_fd_sc_hd__or3_2
X_14139_ net408 net138 _04107_ _04110_ VGND VGND VPWR VPWR _04111_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_10_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout409 net410 VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__buf_2
X_18947_ _09390_ _09399_ VGND VGND VPWR VPWR _09400_ sky130_fd_sc_hd__xnor2_1
X_09680_ net49 _03614_ _03647_ ki\[18\] VGND VGND VPWR VPWR _00047_ sky130_fd_sc_hd__a22o_1
X_18878_ _09306_ _09323_ VGND VGND VPWR VPWR _09324_ sky130_fd_sc_hd__xnor2_1
X_17829_ ki\[4\] _07094_ VGND VGND VPWR VPWR _08170_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09947_ _06458_ _06733_ _06755_ VGND VGND VPWR VPWR _06766_ sky130_fd_sc_hd__a21oi_1
X_09878_ _05996_ VGND VGND VPWR VPWR _06007_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11840_ net111 VGND VGND VPWR VPWR _01779_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11771_ _00242_ prev_error\[6\] VGND VGND VPWR VPWR _01710_ sky130_fd_sc_hd__or2b_2
XFILLER_0_95_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13510_ _03465_ _03468_ VGND VGND VPWR VPWR _03469_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10722_ _00659_ _00660_ VGND VGND VPWR VPWR _00661_ sky130_fd_sc_hd__xnor2_4
X_14490_ net451 net139 net133 net458 VGND VGND VPWR VPWR _04497_ sky130_fd_sc_hd__a22oi_2
X_13441_ _03394_ _03397_ _03399_ VGND VGND VPWR VPWR _03400_ sky130_fd_sc_hd__o21a_1
X_10653_ _00506_ _00591_ VGND VGND VPWR VPWR _00592_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16160_ _06306_ _06333_ VGND VGND VPWR VPWR _06334_ sky130_fd_sc_hd__nor2_8
X_13372_ _03320_ _03323_ _03249_ _03324_ VGND VGND VPWR VPWR _03325_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_24_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10584_ _00522_ VGND VGND VPWR VPWR _00523_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15111_ _05081_ _05179_ VGND VGND VPWR VPWR _05180_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12323_ _02259_ _02261_ VGND VGND VPWR VPWR _02262_ sky130_fd_sc_hd__and2_1
X_16091_ _06220_ _06257_ VGND VGND VPWR VPWR _06258_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15042_ _05099_ _05103_ VGND VGND VPWR VPWR _05104_ sky130_fd_sc_hd__nor2_1
X_12254_ net226 _01807_ _01814_ net230 VGND VGND VPWR VPWR _02193_ sky130_fd_sc_hd__a22o_1
X_11205_ _01139_ _01143_ VGND VGND VPWR VPWR _01144_ sky130_fd_sc_hd__and2b_1
X_12185_ _01961_ _01955_ VGND VGND VPWR VPWR _02124_ sky130_fd_sc_hd__or2b_1
XFILLER_0_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18801_ _09237_ _09238_ VGND VGND VPWR VPWR _09239_ sky130_fd_sc_hd__nor2_1
X_11136_ _01066_ _01073_ _01074_ VGND VGND VPWR VPWR _01075_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16993_ _07189_ _07249_ VGND VGND VPWR VPWR _07251_ sky130_fd_sc_hd__nand2_1
X_18732_ _09151_ _09152_ _09161_ VGND VGND VPWR VPWR _09163_ sky130_fd_sc_hd__a21oi_1
X_15944_ _06072_ _06074_ VGND VGND VPWR VPWR _06097_ sky130_fd_sc_hd__or2_1
X_11067_ _01000_ _01005_ VGND VGND VPWR VPWR _01006_ sky130_fd_sc_hd__xor2_1
X_10018_ _07525_ _07536_ VGND VGND VPWR VPWR _07547_ sky130_fd_sc_hd__or2_1
X_15875_ _05998_ _06020_ VGND VGND VPWR VPWR _06021_ sky130_fd_sc_hd__nor2_2
X_18663_ _06098_ _06080_ _06096_ VGND VGND VPWR VPWR _09088_ sky130_fd_sc_hd__nand3_1
XFILLER_0_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14826_ _04762_ _04866_ VGND VGND VPWR VPWR _04867_ sky130_fd_sc_hd__nor2_1
X_17614_ _07927_ _07930_ _07933_ VGND VGND VPWR VPWR _07934_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18594_ _06118_ _06034_ _06116_ VGND VGND VPWR VPWR _09012_ sky130_fd_sc_hd__nand3_1
X_14757_ _04744_ _04790_ VGND VGND VPWR VPWR _04791_ sky130_fd_sc_hd__nand2_1
X_17545_ _07817_ _07857_ VGND VGND VPWR VPWR _07858_ sky130_fd_sc_hd__and2_1
XFILLER_0_157_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11969_ _01907_ VGND VGND VPWR VPWR _01908_ sky130_fd_sc_hd__buf_2
XFILLER_0_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13708_ net256 _02639_ _03637_ VGND VGND VPWR VPWR _03674_ sky130_fd_sc_hd__a21oi_1
X_17476_ _07737_ _07751_ _07750_ VGND VGND VPWR VPWR _07782_ sky130_fd_sc_hd__o21ba_1
X_14688_ _04713_ _04714_ VGND VGND VPWR VPWR _04715_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19215_ clknet_4_4_0_clock _00097_ VGND VGND VPWR VPWR prev_error\[2\] sky130_fd_sc_hd__dfxtp_2
X_16427_ _06453_ _06627_ VGND VGND VPWR VPWR _06628_ sky130_fd_sc_hd__or2_1
X_13639_ _03539_ _03595_ _03589_ _03594_ VGND VGND VPWR VPWR _03599_ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19146_ net504 i_error\[14\] VGND VGND VPWR VPWR _09567_ sky130_fd_sc_hd__or2_1
X_16358_ _06551_ VGND VGND VPWR VPWR _06552_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15309_ net453 net178 net172 net459 VGND VGND VPWR VPWR _05398_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19077_ net498 prev_error\[0\] VGND VGND VPWR VPWR _09524_ sky130_fd_sc_hd__or2_1
X_16289_ _06454_ _06459_ _06461_ VGND VGND VPWR VPWR _06476_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18028_ _08381_ _08384_ VGND VGND VPWR VPWR _08389_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout206 net207 VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout217 net219 VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__buf_2
X_09801_ _05138_ _05149_ VGND VGND VPWR VPWR _05160_ sky130_fd_sc_hd__and2_4
XFILLER_0_5_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout228 net229 VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout239 net240 VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__buf_2
X_09732_ net76 net18 VGND VGND VPWR VPWR _04401_ sky130_fd_sc_hd__or2b_1
X_09663_ net50 _03625_ _03658_ net330 VGND VGND VPWR VPWR _00048_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13990_ _03909_ _03955_ VGND VGND VPWR VPWR _03962_ sky130_fd_sc_hd__xnor2_1
X_12941_ net267 _01834_ VGND VGND VPWR VPWR _02880_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15660_ _05736_ _05783_ VGND VGND VPWR VPWR _05784_ sky130_fd_sc_hd__nand2_1
X_12872_ _02803_ _02798_ VGND VGND VPWR VPWR _02811_ sky130_fd_sc_hd__and2b_1
X_14611_ _04628_ _04620_ _04626_ VGND VGND VPWR VPWR _04630_ sky130_fd_sc_hd__nor3_1
X_11823_ net250 _01761_ VGND VGND VPWR VPWR _01762_ sky130_fd_sc_hd__nand2_1
X_15591_ _05696_ _05685_ _05694_ VGND VGND VPWR VPWR _05708_ sky130_fd_sc_hd__nand3_1
XFILLER_0_139_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17330_ net306 _06467_ VGND VGND VPWR VPWR _07621_ sky130_fd_sc_hd__nand2_1
X_14542_ _04516_ _04535_ _04552_ VGND VGND VPWR VPWR _04554_ sky130_fd_sc_hd__nand3_1
XFILLER_0_96_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11754_ _00462_ _00561_ VGND VGND VPWR VPWR _01693_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17261_ _07532_ _07533_ _07544_ VGND VGND VPWR VPWR _07545_ sky130_fd_sc_hd__or3_4
X_10705_ _00633_ _00643_ VGND VGND VPWR VPWR _00644_ sky130_fd_sc_hd__xor2_4
XFILLER_0_153_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14473_ _04475_ _04470_ _04474_ VGND VGND VPWR VPWR _04479_ sky130_fd_sc_hd__nor3_1
XFILLER_0_83_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11685_ _01617_ _01621_ VGND VGND VPWR VPWR _01624_ sky130_fd_sc_hd__xor2_1
X_19000_ _09194_ _09457_ VGND VGND VPWR VPWR _09458_ sky130_fd_sc_hd__xnor2_1
X_16212_ _06388_ _06390_ VGND VGND VPWR VPWR _06391_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13424_ _03379_ _03381_ VGND VGND VPWR VPWR _03382_ sky130_fd_sc_hd__nand2_1
X_17192_ _07466_ _07467_ _07468_ VGND VGND VPWR VPWR _07469_ sky130_fd_sc_hd__nand3_1
X_10636_ _00569_ _00571_ VGND VGND VPWR VPWR _00575_ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16143_ _06314_ VGND VGND VPWR VPWR _06316_ sky130_fd_sc_hd__buf_2
XFILLER_0_3_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13355_ net258 _01907_ _01872_ kd_1\[2\] VGND VGND VPWR VPWR _03308_ sky130_fd_sc_hd__a22oi_1
X_10567_ net347 _00245_ _00505_ VGND VGND VPWR VPWR _00506_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12306_ _02073_ _02110_ _02109_ VGND VGND VPWR VPWR _02245_ sky130_fd_sc_hd__o21a_1
XFILLER_0_121_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16074_ _06234_ _06239_ VGND VGND VPWR VPWR _06240_ sky130_fd_sc_hd__xnor2_1
X_13286_ _03237_ _03238_ VGND VGND VPWR VPWR _03239_ sky130_fd_sc_hd__nor2_1
X_10498_ _00365_ _00366_ VGND VGND VPWR VPWR _00437_ sky130_fd_sc_hd__xnor2_4
X_15025_ _05084_ _05085_ VGND VGND VPWR VPWR _05086_ sky130_fd_sc_hd__nor2_1
X_12237_ net242 _01779_ _01786_ net238 VGND VGND VPWR VPWR _02176_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_20_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12168_ _02102_ _02106_ VGND VGND VPWR VPWR _02107_ sky130_fd_sc_hd__or2b_1
X_11119_ _00966_ _01046_ _01051_ VGND VGND VPWR VPWR _01058_ sky130_fd_sc_hd__a21o_1
X_16976_ net294 _06620_ VGND VGND VPWR VPWR _07232_ sky130_fd_sc_hd__nand2_1
X_12099_ _01769_ _01779_ VGND VGND VPWR VPWR _02038_ sky130_fd_sc_hd__and2b_1
X_18715_ _09139_ _09140_ _09144_ VGND VGND VPWR VPWR _09145_ sky130_fd_sc_hd__a21o_1
X_15927_ _03852_ _03553_ _03851_ VGND VGND VPWR VPWR _06078_ sky130_fd_sc_hd__nor3_1
Xinput6 measurement[13] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
X_18646_ _06162_ _09068_ VGND VGND VPWR VPWR _09069_ sky130_fd_sc_hd__and2_1
X_15858_ _04304_ _06001_ _04382_ VGND VGND VPWR VPWR _06002_ sky130_fd_sc_hd__a21o_1
XFILLER_0_149_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14809_ _04845_ _04846_ _04836_ _04840_ VGND VGND VPWR VPWR _04848_ sky130_fd_sc_hd__a211o_1
X_18577_ _08987_ _08991_ VGND VGND VPWR VPWR _08993_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_143_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15789_ _05868_ _05912_ _05905_ _05910_ VGND VGND VPWR VPWR _05926_ sky130_fd_sc_hd__or4_1
XFILLER_0_87_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17528_ _07820_ _07836_ _07838_ VGND VGND VPWR VPWR _07839_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17459_ _07687_ _07761_ _07760_ _07762_ VGND VGND VPWR VPWR _07763_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_27_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19129_ _09139_ _09140_ _09550_ VGND VGND VPWR VPWR _09556_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09715_ net71 net13 VGND VGND VPWR VPWR _04214_ sky130_fd_sc_hd__or2b_1
XFILLER_0_93_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09646_ net41 _03347_ _03380_ net227 VGND VGND VPWR VPWR _00001_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11470_ _01407_ _01408_ VGND VGND VPWR VPWR _01409_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10421_ _00190_ _00279_ _00281_ VGND VGND VPWR VPWR _00360_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13140_ _02986_ _03085_ VGND VGND VPWR VPWR _03088_ sky130_fd_sc_hd__and2_1
XFILLER_0_61_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10352_ net361 _06007_ VGND VGND VPWR VPWR _00291_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13071_ net236 _02090_ VGND VGND VPWR VPWR _03012_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10283_ _00204_ _00217_ VGND VGND VPWR VPWR _00222_ sky130_fd_sc_hd__or2_1
X_12022_ _01956_ _01960_ VGND VGND VPWR VPWR _01961_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16830_ net294 _06468_ _07070_ VGND VGND VPWR VPWR _07071_ sky130_fd_sc_hd__and3_1
X_16761_ net278 _06802_ _06891_ net274 VGND VGND VPWR VPWR _06995_ sky130_fd_sc_hd__a22o_1
X_13973_ net426 net567 net128 net126 VGND VGND VPWR VPWR _03945_ sky130_fd_sc_hd__and4_1
X_18500_ _06265_ _08836_ VGND VGND VPWR VPWR _08908_ sky130_fd_sc_hd__or2_1
X_15712_ _05838_ _05840_ VGND VGND VPWR VPWR _05841_ sky130_fd_sc_hd__or2_1
X_12924_ _02840_ _02862_ VGND VGND VPWR VPWR _02863_ sky130_fd_sc_hd__xnor2_1
X_16692_ _06908_ _06918_ VGND VGND VPWR VPWR _06919_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18431_ _08831_ _08585_ VGND VGND VPWR VPWR _08832_ sky130_fd_sc_hd__and2_1
X_15643_ _05762_ _05763_ VGND VGND VPWR VPWR _05766_ sky130_fd_sc_hd__nor2_1
X_12855_ _02778_ _02781_ VGND VGND VPWR VPWR _02794_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11806_ _01739_ _01743_ _01744_ VGND VGND VPWR VPWR _01745_ sky130_fd_sc_hd__a21oi_4
X_15574_ net462 net183 VGND VGND VPWR VPWR _05690_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18362_ _06171_ _08616_ VGND VGND VPWR VPWR _08756_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12786_ _02647_ _02649_ VGND VGND VPWR VPWR _02725_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14525_ _04016_ net175 VGND VGND VPWR VPWR _04536_ sky130_fd_sc_hd__nor2_1
X_17313_ _07532_ _07533_ _07544_ VGND VGND VPWR VPWR _07603_ sky130_fd_sc_hd__nor3_1
X_11737_ _01409_ _01350_ _01351_ VGND VGND VPWR VPWR _01676_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18293_ _08678_ _08679_ VGND VGND VPWR VPWR _08681_ sky130_fd_sc_hd__xor2_2
XFILLER_0_22_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14456_ _04458_ _04449_ _04455_ VGND VGND VPWR VPWR _04460_ sky130_fd_sc_hd__and3_1
XFILLER_0_83_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17244_ net566 net316 _06334_ _06401_ VGND VGND VPWR VPWR _07527_ sky130_fd_sc_hd__and4_1
XFILLER_0_154_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11668_ _01593_ _01602_ _01606_ VGND VGND VPWR VPWR _01607_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13407_ _03353_ _03348_ VGND VGND VPWR VPWR _03363_ sky130_fd_sc_hd__and2b_1
X_17175_ _07447_ _07449_ _07450_ VGND VGND VPWR VPWR _07451_ sky130_fd_sc_hd__a21oi_1
X_10619_ _00466_ _00553_ _00557_ VGND VGND VPWR VPWR _00558_ sky130_fd_sc_hd__o21a_2
X_14387_ _04382_ _04383_ VGND VGND VPWR VPWR _04384_ sky130_fd_sc_hd__or2b_1
X_11599_ _01535_ _01536_ _01537_ VGND VGND VPWR VPWR _01538_ sky130_fd_sc_hd__nand3_1
XFILLER_0_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16126_ net115 _06289_ _06296_ VGND VGND VPWR VPWR _06297_ sky130_fd_sc_hd__a21o_2
X_13338_ net233 net228 _02544_ _02640_ VGND VGND VPWR VPWR _03291_ sky130_fd_sc_hd__and4_1
XFILLER_0_51_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16057_ _09043_ _06176_ _06219_ VGND VGND VPWR VPWR _06221_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13269_ _03221_ _03129_ VGND VGND VPWR VPWR _03222_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15008_ net427 net184 net181 net432 VGND VGND VPWR VPWR _05067_ sky130_fd_sc_hd__a22o_1
X_16959_ net305 _06401_ VGND VGND VPWR VPWR _07213_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18629_ _08833_ _09049_ _08882_ VGND VGND VPWR VPWR _09050_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_11 kp\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_22 net369 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_33 net335 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10970_ _00907_ _00908_ VGND VGND VPWR VPWR _00909_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09629_ net49 _03091_ _03124_ net553 VGND VGND VPWR VPWR _00028_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12640_ net259 net255 _01785_ _01798_ VGND VGND VPWR VPWR _02579_ sky130_fd_sc_hd__and4_1
XFILLER_0_77_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12571_ _02380_ _02507_ _02509_ VGND VGND VPWR VPWR _02510_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_66_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14310_ _04297_ _04158_ _04298_ VGND VGND VPWR VPWR _04299_ sky130_fd_sc_hd__and3_1
X_11522_ _01459_ _01460_ VGND VGND VPWR VPWR _01461_ sky130_fd_sc_hd__and2_1
XFILLER_0_136_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15290_ _05374_ _05376_ VGND VGND VPWR VPWR _05377_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14241_ _03896_ _04222_ VGND VGND VPWR VPWR _04223_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11453_ _01360_ _01363_ VGND VGND VPWR VPWR _01392_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10404_ _00319_ _00340_ _00342_ VGND VGND VPWR VPWR _00343_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14172_ _03916_ _04088_ _04146_ VGND VGND VPWR VPWR _04147_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11384_ _01260_ _01318_ _01322_ VGND VGND VPWR VPWR _01323_ sky130_fd_sc_hd__nand3_1
XFILLER_0_110_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13123_ _03055_ _03068_ VGND VGND VPWR VPWR _03070_ sky130_fd_sc_hd__xor2_1
X_10335_ net372 _05182_ VGND VGND VPWR VPWR _00274_ sky130_fd_sc_hd__nand2_1
X_18980_ _09367_ _09435_ VGND VGND VPWR VPWR _09436_ sky130_fd_sc_hd__xnor2_1
X_13054_ _02991_ _02993_ VGND VGND VPWR VPWR _02994_ sky130_fd_sc_hd__xnor2_1
X_17931_ _08239_ _08241_ VGND VGND VPWR VPWR _08282_ sky130_fd_sc_hd__xnor2_1
X_10266_ net360 _05325_ VGND VGND VPWR VPWR _00205_ sky130_fd_sc_hd__nand2_1
X_12005_ _01939_ _01943_ VGND VGND VPWR VPWR _01944_ sky130_fd_sc_hd__xor2_1
X_17862_ _08193_ _08198_ VGND VGND VPWR VPWR _08206_ sky130_fd_sc_hd__or2_1
X_10197_ net354 _05996_ _08273_ VGND VGND VPWR VPWR _09507_ sky130_fd_sc_hd__a21oi_1
X_16813_ net304 _06345_ VGND VGND VPWR VPWR _07053_ sky130_fd_sc_hd__nand2_1
X_17793_ _08120_ _08121_ _08128_ VGND VGND VPWR VPWR _08131_ sky130_fd_sc_hd__and3_1
X_16744_ _06902_ _06976_ VGND VGND VPWR VPWR _06977_ sky130_fd_sc_hd__nor2_1
X_13956_ net438 net444 net123 net120 VGND VGND VPWR VPWR _03928_ sky130_fd_sc_hd__and4_1
XFILLER_0_88_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12907_ net202 _02747_ VGND VGND VPWR VPWR _02846_ sky130_fd_sc_hd__nand2_1
X_16675_ _06879_ _06897_ VGND VGND VPWR VPWR _06901_ sky130_fd_sc_hd__xnor2_1
X_13887_ _03553_ _03851_ _03852_ VGND VGND VPWR VPWR _03853_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18414_ _08797_ _08804_ _08805_ _08806_ _08813_ VGND VGND VPWR VPWR _08814_ sky130_fd_sc_hd__a311o_1
X_15626_ _05745_ _05746_ VGND VGND VPWR VPWR _05747_ sky130_fd_sc_hd__and2b_1
X_12838_ _02694_ _02776_ VGND VGND VPWR VPWR _02777_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18345_ _08534_ _08611_ _08736_ VGND VGND VPWR VPWR _08738_ sky130_fd_sc_hd__and3_1
X_12769_ _02695_ _02681_ VGND VGND VPWR VPWR _02708_ sky130_fd_sc_hd__or2b_1
X_15557_ _05612_ _05670_ VGND VGND VPWR VPWR _05671_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14508_ net445 net152 VGND VGND VPWR VPWR _04517_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15488_ _05508_ _05594_ VGND VGND VPWR VPWR _05595_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18276_ _06376_ _08661_ VGND VGND VPWR VPWR _08662_ sky130_fd_sc_hd__xor2_1
XFILLER_0_127_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput20 measurement[9] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
X_17227_ _07506_ _07507_ VGND VGND VPWR VPWR _07508_ sky130_fd_sc_hd__or2b_1
XFILLER_0_141_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14439_ _04439_ _04440_ VGND VGND VPWR VPWR _04441_ sky130_fd_sc_hd__nor2_1
Xinput31 reg_addr[1] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_1
XFILLER_0_142_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput42 reg_data[11] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_4
Xinput53 reg_data[4] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput64 target[13] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_1
X_17158_ _07392_ _07402_ _07431_ VGND VGND VPWR VPWR _07432_ sky130_fd_sc_hd__a21o_1
Xinput75 target[6] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_1
XFILLER_0_40_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16109_ _02744_ _06276_ _06277_ VGND VGND VPWR VPWR _06278_ sky130_fd_sc_hd__a21o_2
X_09980_ _07107_ _07118_ VGND VGND VPWR VPWR _07129_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17089_ _07355_ _07127_ VGND VGND VPWR VPWR _07356_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_149_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_150_Left_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10120_ _08548_ _08658_ VGND VGND VPWR VPWR _08669_ sky130_fd_sc_hd__and2_1
XFILLER_0_101_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10051_ _07866_ _07899_ VGND VGND VPWR VPWR _07910_ sky130_fd_sc_hd__nor2_1
X_13810_ _03772_ _03774_ _03775_ VGND VGND VPWR VPWR _03776_ sky130_fd_sc_hd__or3_1
X_14790_ _04813_ _04826_ VGND VGND VPWR VPWR _04827_ sky130_fd_sc_hd__nand2_1
X_13741_ _03695_ _03699_ _03706_ VGND VGND VPWR VPWR _03707_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10953_ net346 _00516_ _00801_ VGND VGND VPWR VPWR _00892_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13672_ _03577_ _03634_ VGND VGND VPWR VPWR _03635_ sky130_fd_sc_hd__or2_1
X_16460_ _06647_ _06663_ VGND VGND VPWR VPWR _06664_ sky130_fd_sc_hd__xor2_2
X_10884_ _00803_ _00806_ _00822_ VGND VGND VPWR VPWR _00823_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_39_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12623_ _02473_ _02528_ _02561_ VGND VGND VPWR VPWR _02562_ sky130_fd_sc_hd__o21a_1
X_15411_ _05422_ _05509_ VGND VGND VPWR VPWR _05510_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16391_ _06577_ _06587_ VGND VGND VPWR VPWR _06588_ sky130_fd_sc_hd__xnor2_1
X_15342_ _05393_ _05395_ VGND VGND VPWR VPWR _05434_ sky130_fd_sc_hd__or2b_1
X_18130_ _08441_ _08483_ _08495_ _08498_ _08500_ VGND VGND VPWR VPWR _08501_ sky130_fd_sc_hd__a311o_2
X_12554_ net254 _01785_ _02427_ VGND VGND VPWR VPWR _02493_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11505_ _01432_ _01441_ VGND VGND VPWR VPWR _01444_ sky130_fd_sc_hd__xor2_1
X_15273_ _05355_ _05356_ _05344_ _05350_ VGND VGND VPWR VPWR _05359_ sky130_fd_sc_hd__a211o_1
X_18061_ _08158_ _08169_ _08222_ VGND VGND VPWR VPWR _08425_ sky130_fd_sc_hd__a21oi_1
X_12485_ _02362_ _02365_ VGND VGND VPWR VPWR _02424_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14224_ _04202_ _04204_ VGND VGND VPWR VPWR _04205_ sky130_fd_sc_hd__xnor2_1
X_17012_ _07251_ _07260_ _07270_ VGND VGND VPWR VPWR _07271_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11436_ _01374_ _01320_ VGND VGND VPWR VPWR _01375_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14155_ _03902_ _03907_ VGND VGND VPWR VPWR _04129_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11367_ net358 _00810_ _01305_ VGND VGND VPWR VPWR _01306_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13106_ _03040_ _03043_ _03050_ VGND VGND VPWR VPWR _03051_ sky130_fd_sc_hd__o21ai_1
X_10318_ _00255_ _00256_ VGND VGND VPWR VPWR _00257_ sky130_fd_sc_hd__nor2_1
X_14086_ _04056_ _04057_ VGND VGND VPWR VPWR _04058_ sky130_fd_sc_hd__nand2_1
X_18963_ _09413_ _09416_ VGND VGND VPWR VPWR _09418_ sky130_fd_sc_hd__xnor2_1
X_11298_ net565 _00811_ VGND VGND VPWR VPWR _01237_ sky130_fd_sc_hd__nand2_2
XFILLER_0_28_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13037_ _02944_ _02912_ VGND VGND VPWR VPWR _02976_ sky130_fd_sc_hd__or2b_1
X_17914_ _08256_ _08261_ _08260_ VGND VGND VPWR VPWR _08264_ sky130_fd_sc_hd__o21ai_1
X_10249_ _00166_ _00168_ VGND VGND VPWR VPWR _00188_ sky130_fd_sc_hd__xnor2_1
X_18894_ _09278_ _09339_ VGND VGND VPWR VPWR _09342_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17845_ net331 _07094_ VGND VGND VPWR VPWR _08188_ sky130_fd_sc_hd__and2_1
X_17776_ _08110_ _08111_ VGND VGND VPWR VPWR _08112_ sky130_fd_sc_hd__xnor2_1
X_14988_ _05043_ _05041_ VGND VGND VPWR VPWR _05045_ sky130_fd_sc_hd__xnor2_1
X_16727_ net293 _06402_ VGND VGND VPWR VPWR _06958_ sky130_fd_sc_hd__nand2_1
X_13939_ _03895_ _03893_ VGND VGND VPWR VPWR _03910_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16658_ net284 _06621_ _06881_ VGND VGND VPWR VPWR _06882_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15609_ _05634_ _05667_ _05665_ VGND VGND VPWR VPWR _05728_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16589_ net271 _06803_ _06804_ _06805_ VGND VGND VPWR VPWR _06806_ sky130_fd_sc_hd__a31o_1
XFILLER_0_84_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18328_ ki\[14\] _06328_ VGND VGND VPWR VPWR _08719_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18259_ _06519_ _06522_ _08642_ VGND VGND VPWR VPWR _08643_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09963_ _06931_ _05677_ _05710_ VGND VGND VPWR VPWR _06942_ sky130_fd_sc_hd__or3b_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09894_ _06172_ VGND VGND VPWR VPWR _06183_ sky130_fd_sc_hd__buf_4
XFILLER_0_68_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12270_ _02186_ _02207_ _02071_ _02208_ VGND VGND VPWR VPWR _02209_ sky130_fd_sc_hd__a211o_2
X_11221_ _01158_ _01159_ VGND VGND VPWR VPWR _01160_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11152_ net367 net362 _00409_ _01001_ VGND VGND VPWR VPWR _01091_ sky130_fd_sc_hd__nand4_1
XFILLER_0_101_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10103_ _08449_ _08471_ VGND VGND VPWR VPWR _08482_ sky130_fd_sc_hd__or2b_1
X_15960_ _06046_ _06112_ _06113_ VGND VGND VPWR VPWR _06114_ sky130_fd_sc_hd__a21o_1
X_11083_ _00996_ _01018_ _01020_ VGND VGND VPWR VPWR _01022_ sky130_fd_sc_hd__nor3_1
X_10034_ _07701_ _07712_ VGND VGND VPWR VPWR _07723_ sky130_fd_sc_hd__and2b_1
X_14911_ net472 net474 net138 net134 VGND VGND VPWR VPWR _04960_ sky130_fd_sc_hd__and4_1
X_15891_ _05981_ _06037_ _04787_ VGND VGND VPWR VPWR _06038_ sky130_fd_sc_hd__o21ai_1
X_17630_ _07861_ _07864_ _07863_ VGND VGND VPWR VPWR _07951_ sky130_fd_sc_hd__o21a_1
X_14842_ _04773_ _04776_ VGND VGND VPWR VPWR _04884_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17561_ _07655_ _07656_ _07691_ VGND VGND VPWR VPWR _07875_ sky130_fd_sc_hd__or3_1
X_14773_ _04794_ _04799_ VGND VGND VPWR VPWR _04809_ sky130_fd_sc_hd__xor2_1
X_11985_ _01921_ _01923_ VGND VGND VPWR VPWR _01924_ sky130_fd_sc_hd__or2b_1
X_19300_ clknet_4_8_0_clock _00040_ VGND VGND VPWR VPWR ki\[11\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_98_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16512_ _06720_ VGND VGND VPWR VPWR _06721_ sky130_fd_sc_hd__buf_2
X_13724_ _03679_ _03687_ _03689_ VGND VGND VPWR VPWR _03690_ sky130_fd_sc_hd__o21a_1
X_10936_ _00771_ _00770_ VGND VGND VPWR VPWR _00875_ sky130_fd_sc_hd__nor2_1
X_17492_ _06399_ _03220_ VGND VGND VPWR VPWR _07799_ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19231_ clknet_4_5_0_clock _00113_ VGND VGND VPWR VPWR prev_error\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16443_ _06613_ _06615_ _06644_ VGND VGND VPWR VPWR _06646_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_129_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13655_ net237 _02914_ VGND VGND VPWR VPWR _03617_ sky130_fd_sc_hd__nand2_1
X_10867_ _00804_ _00805_ VGND VGND VPWR VPWR _00806_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12606_ _02544_ VGND VGND VPWR VPWR _02545_ sky130_fd_sc_hd__buf_2
XFILLER_0_54_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19162_ net501 prev_d_error\[3\] VGND VGND VPWR VPWR _09576_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13586_ _03541_ _03543_ _03544_ VGND VGND VPWR VPWR _03545_ sky130_fd_sc_hd__nand3_2
X_16374_ _06567_ _06569_ VGND VGND VPWR VPWR _06570_ sky130_fd_sc_hd__or2_1
X_10798_ _00732_ _00733_ _00736_ VGND VGND VPWR VPWR _00737_ sky130_fd_sc_hd__a21boi_2
X_18113_ _08478_ _08481_ VGND VGND VPWR VPWR _08483_ sky130_fd_sc_hd__and2_1
X_12537_ net250 _01786_ _01761_ VGND VGND VPWR VPWR _02476_ sky130_fd_sc_hd__a21oi_1
X_15325_ _05412_ _05415_ VGND VGND VPWR VPWR _05416_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19093_ net499 prev_error\[8\] VGND VGND VPWR VPWR _09534_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18044_ _08338_ _08343_ _08292_ _08344_ VGND VGND VPWR VPWR _08407_ sky130_fd_sc_hd__a211o_1
XFILLER_0_81_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15256_ net442 net447 net184 net181 VGND VGND VPWR VPWR _05340_ sky130_fd_sc_hd__and4_1
X_12468_ _01723_ _02406_ VGND VGND VPWR VPWR _02407_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_152_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14207_ _04118_ _04162_ _04185_ VGND VGND VPWR VPWR _04186_ sky130_fd_sc_hd__a21oi_1
X_11419_ net564 _00243_ VGND VGND VPWR VPWR _01358_ sky130_fd_sc_hd__nand2_1
X_15187_ _05135_ _05207_ _05240_ _05263_ VGND VGND VPWR VPWR _05264_ sky130_fd_sc_hd__a31oi_1
X_12399_ _02313_ _02337_ VGND VGND VPWR VPWR _02338_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_111_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14138_ _04108_ VGND VGND VPWR VPWR _04110_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18946_ _09391_ _09398_ VGND VGND VPWR VPWR _09399_ sky130_fd_sc_hd__xnor2_1
X_14069_ _04015_ _04021_ _04039_ _04040_ VGND VGND VPWR VPWR _04041_ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18877_ _09321_ _09322_ VGND VGND VPWR VPWR _09323_ sky130_fd_sc_hd__nor2_1
X_17828_ _08156_ _08157_ _08145_ _08147_ VGND VGND VPWR VPWR _08169_ sky130_fd_sc_hd__a211o_1
XFILLER_0_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17759_ _07999_ _08085_ VGND VGND VPWR VPWR _08093_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09946_ _06194_ _06744_ net568 VGND VGND VPWR VPWR _06755_ sky130_fd_sc_hd__and3b_1
X_09877_ _05985_ VGND VGND VPWR VPWR _05996_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11770_ _06579_ _08163_ prev_error\[8\] VGND VGND VPWR VPWR _01709_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_56_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10721_ _00465_ _00558_ VGND VGND VPWR VPWR _00660_ sky130_fd_sc_hd__xor2_4
X_13440_ _03289_ _03398_ VGND VGND VPWR VPWR _03399_ sky130_fd_sc_hd__xnor2_1
X_10652_ net347 _00245_ _00505_ VGND VGND VPWR VPWR _00591_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13371_ _03246_ _03247_ _03248_ VGND VGND VPWR VPWR _03324_ sky130_fd_sc_hd__o21a_1
X_10583_ _00507_ _00511_ _00521_ VGND VGND VPWR VPWR _00522_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_23_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12322_ _02175_ _02260_ VGND VGND VPWR VPWR _02261_ sky130_fd_sc_hd__xnor2_1
X_15110_ net410 net194 _05080_ VGND VGND VPWR VPWR _05179_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16090_ _06255_ _06256_ VGND VGND VPWR VPWR _06257_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15041_ _05098_ _05092_ _05097_ VGND VGND VPWR VPWR _05103_ sky130_fd_sc_hd__and3_1
X_12253_ _02054_ _02056_ VGND VGND VPWR VPWR _02192_ sky130_fd_sc_hd__xnor2_1
X_11204_ net383 _08196_ _01141_ _01142_ VGND VGND VPWR VPWR _01143_ sky130_fd_sc_hd__a31o_1
X_12184_ _01956_ _01960_ VGND VGND VPWR VPWR _02123_ sky130_fd_sc_hd__nand2_1
X_18800_ _04131_ _04193_ _09236_ VGND VGND VPWR VPWR _09238_ sky130_fd_sc_hd__nor3_1
X_11135_ _01068_ _01069_ _01072_ VGND VGND VPWR VPWR _01074_ sky130_fd_sc_hd__or3_1
X_16992_ _07187_ _07188_ VGND VGND VPWR VPWR _07249_ sky130_fd_sc_hd__or2_1
X_18731_ _09151_ _09152_ _09161_ VGND VGND VPWR VPWR _09162_ sky130_fd_sc_hd__and3_1
X_15943_ _06083_ _06092_ _06094_ VGND VGND VPWR VPWR _06096_ sky130_fd_sc_hd__a21o_1
X_11066_ net358 _00410_ _01004_ _01002_ VGND VGND VPWR VPWR _01005_ sky130_fd_sc_hd__a31o_1
X_10017_ _07393_ _07514_ VGND VGND VPWR VPWR _07536_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18662_ _09072_ _09085_ VGND VGND VPWR VPWR _09086_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15874_ _05994_ _05997_ _04477_ VGND VGND VPWR VPWR _06020_ sky130_fd_sc_hd__a21oi_1
X_17613_ _07824_ _07931_ VGND VGND VPWR VPWR _07933_ sky130_fd_sc_hd__nor2_1
X_14825_ net409 net190 _04760_ _04865_ VGND VGND VPWR VPWR _04866_ sky130_fd_sc_hd__o2bb2a_1
X_18593_ _09006_ _09009_ VGND VGND VPWR VPWR _09011_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17544_ _07815_ _07816_ VGND VGND VPWR VPWR _07857_ sky130_fd_sc_hd__or2_1
X_14756_ _04740_ _04743_ VGND VGND VPWR VPWR _04790_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11968_ _01905_ _01906_ VGND VGND VPWR VPWR _01907_ sky130_fd_sc_hd__xor2_4
XFILLER_0_156_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13707_ net256 _02639_ _03637_ VGND VGND VPWR VPWR _03673_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10919_ _00828_ _00856_ _00857_ VGND VGND VPWR VPWR _00858_ sky130_fd_sc_hd__a21oi_1
X_17475_ _07769_ _07780_ VGND VGND VPWR VPWR _07781_ sky130_fd_sc_hd__xnor2_2
X_11899_ net213 _01808_ _01815_ VGND VGND VPWR VPWR _01838_ sky130_fd_sc_hd__a21oi_1
X_14687_ _04712_ _04705_ VGND VGND VPWR VPWR _04714_ sky130_fd_sc_hd__or2b_1
XFILLER_0_41_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19214_ clknet_4_4_0_clock _00096_ VGND VGND VPWR VPWR prev_error\[1\] sky130_fd_sc_hd__dfxtp_2
X_16426_ net286 _06410_ VGND VGND VPWR VPWR _06627_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13638_ _03573_ _03597_ VGND VGND VPWR VPWR _03598_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19145_ net504 i_error\[13\] net495 _09566_ VGND VGND VPWR VPWR _00127_ sky130_fd_sc_hd__o211a_1
X_16357_ _06541_ _06550_ VGND VGND VPWR VPWR _06551_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13569_ net266 _01909_ _03467_ VGND VGND VPWR VPWR _03528_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15308_ net449 net182 VGND VGND VPWR VPWR _05397_ sky130_fd_sc_hd__nand2_1
X_19076_ net563 VGND VGND VPWR VPWR _09523_ sky130_fd_sc_hd__buf_4
X_16288_ _06471_ _06472_ _06474_ VGND VGND VPWR VPWR _06475_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_30_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18027_ _08385_ _08386_ VGND VGND VPWR VPWR _08388_ sky130_fd_sc_hd__nor2_1
X_15239_ _05309_ _05318_ _05320_ VGND VGND VPWR VPWR _05321_ sky130_fd_sc_hd__a21o_1
XFILLER_0_140_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout207 kd_1\[15\] VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_4
X_09800_ _04170_ _04764_ _05127_ VGND VGND VPWR VPWR _05149_ sky130_fd_sc_hd__nand3_4
Xfanout218 net219 VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__buf_2
Xfanout229 kd_1\[10\] VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__buf_2
XFILLER_0_157_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18929_ _09284_ _09301_ VGND VGND VPWR VPWR _09380_ sky130_fd_sc_hd__and2b_1
X_09731_ net18 net76 VGND VGND VPWR VPWR _04390_ sky130_fd_sc_hd__or2b_1
XFILLER_0_66_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09662_ net40 _03625_ _03658_ net334 VGND VGND VPWR VPWR _00038_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_19_Left_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_28_Left_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09929_ net341 _06007_ _06557_ VGND VGND VPWR VPWR _06568_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_130_Right_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12940_ net250 _01834_ _01785_ net268 VGND VGND VPWR VPWR _02879_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_99_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_37_Left_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12871_ _02797_ _02795_ VGND VGND VPWR VPWR _02810_ sky130_fd_sc_hd__and2b_1
X_14610_ _04620_ _04626_ _04628_ VGND VGND VPWR VPWR _04629_ sky130_fd_sc_hd__o21a_1
X_11822_ _01760_ VGND VGND VPWR VPWR _01761_ sky130_fd_sc_hd__dlymetal6s2s_1
X_15590_ _05702_ _05706_ VGND VGND VPWR VPWR _05707_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14541_ _04516_ _04535_ _04552_ VGND VGND VPWR VPWR _04553_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11753_ _00661_ _00759_ _01690_ _01691_ _00660_ VGND VGND VPWR VPWR _01692_ sky130_fd_sc_hd__a32o_2
XFILLER_0_83_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10704_ _00636_ _00641_ _00642_ VGND VGND VPWR VPWR _00643_ sky130_fd_sc_hd__a21boi_4
X_17260_ _07534_ _07543_ VGND VGND VPWR VPWR _07544_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_154_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14472_ _04384_ _04476_ VGND VGND VPWR VPWR _04477_ sky130_fd_sc_hd__xnor2_1
X_11684_ _01614_ _01622_ VGND VGND VPWR VPWR _01623_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16211_ net289 _06336_ _06389_ VGND VGND VPWR VPWR _06390_ sky130_fd_sc_hd__and3_1
X_13423_ _03378_ _03373_ VGND VGND VPWR VPWR _03381_ sky130_fd_sc_hd__or2b_1
X_10635_ net371 _06007_ _00572_ _00573_ VGND VGND VPWR VPWR _00574_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_107_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17191_ net328 _06344_ VGND VGND VPWR VPWR _07468_ sky130_fd_sc_hd__and2_1
XFILLER_0_153_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13354_ net262 kd_1\[3\] _01907_ _01872_ VGND VGND VPWR VPWR _03307_ sky130_fd_sc_hd__and4_1
X_16142_ _06313_ _06307_ _01757_ VGND VGND VPWR VPWR _06314_ sky130_fd_sc_hd__a21o_2
X_10566_ net352 _08207_ _00503_ _00504_ VGND VGND VPWR VPWR _00505_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_12_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12305_ _02209_ _02242_ _02243_ VGND VGND VPWR VPWR _02244_ sky130_fd_sc_hd__nand3_2
X_16073_ _06235_ _06237_ VGND VGND VPWR VPWR _06239_ sky130_fd_sc_hd__xnor2_1
X_13285_ net262 _01852_ _01873_ net258 VGND VGND VPWR VPWR _03238_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_87_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10497_ _00304_ _00435_ VGND VGND VPWR VPWR _00436_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12236_ net234 _01799_ VGND VGND VPWR VPWR _02175_ sky130_fd_sc_hd__nand2_1
X_15024_ _05055_ _05057_ _05082_ VGND VGND VPWR VPWR _05085_ sky130_fd_sc_hd__and3_1
X_12167_ _02103_ _02105_ VGND VGND VPWR VPWR _02106_ sky130_fd_sc_hd__xnor2_1
X_11118_ _01055_ _01056_ VGND VGND VPWR VPWR _01057_ sky130_fd_sc_hd__xnor2_1
X_12098_ net242 _01764_ _01779_ net238 VGND VGND VPWR VPWR _02037_ sky130_fd_sc_hd__a22oi_1
X_16975_ _07229_ _07230_ VGND VGND VPWR VPWR _07231_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18714_ _09141_ _09143_ VGND VGND VPWR VPWR _09144_ sky130_fd_sc_hd__nor2_1
X_15926_ _06076_ _05947_ VGND VGND VPWR VPWR _06077_ sky130_fd_sc_hd__xnor2_2
X_11049_ _00975_ _00986_ _00987_ VGND VGND VPWR VPWR _00988_ sky130_fd_sc_hd__nand3_1
Xinput7 measurement[14] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
XFILLER_0_79_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18645_ _09062_ _09066_ VGND VGND VPWR VPWR _09068_ sky130_fd_sc_hd__xnor2_1
X_15857_ _06000_ _05998_ VGND VGND VPWR VPWR _06001_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14808_ _04836_ _04840_ _04845_ _04846_ VGND VGND VPWR VPWR _04847_ sky130_fd_sc_hd__o211ai_2
X_18576_ _08987_ _08991_ VGND VGND VPWR VPWR _08992_ sky130_fd_sc_hd__or2b_1
X_15788_ _05921_ _05924_ _05868_ VGND VGND VPWR VPWR _05925_ sky130_fd_sc_hd__o21ba_1
X_17527_ _07673_ _07837_ VGND VGND VPWR VPWR _07838_ sky130_fd_sc_hd__nand2_1
X_14739_ _04769_ _04770_ VGND VGND VPWR VPWR _04771_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17458_ _07758_ _07759_ _07655_ _07692_ VGND VGND VPWR VPWR _07762_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16409_ _06606_ _06607_ _06604_ VGND VGND VPWR VPWR _06608_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17389_ _07684_ _07685_ VGND VGND VPWR VPWR _07686_ sky130_fd_sc_hd__xor2_1
X_19128_ net506 net559 net494 _09555_ VGND VGND VPWR VPWR _00119_ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19059_ _09510_ _09511_ net495 VGND VGND VPWR VPWR _00087_ sky130_fd_sc_hd__o21a_1
XFILLER_0_140_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09714_ net13 net71 VGND VGND VPWR VPWR _04203_ sky130_fd_sc_hd__or2b_2
X_09645_ net58 _03358_ _03391_ net231 VGND VGND VPWR VPWR _00018_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10420_ _00351_ _00350_ VGND VGND VPWR VPWR _00359_ sky130_fd_sc_hd__xor2_1
XFILLER_0_61_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10351_ _00207_ _00289_ VGND VGND VPWR VPWR _00290_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_131_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13070_ net245 _01908_ VGND VGND VPWR VPWR _03011_ sky130_fd_sc_hd__nand2_1
X_10282_ _00199_ _00220_ VGND VGND VPWR VPWR _00221_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12021_ _01957_ _01959_ VGND VGND VPWR VPWR _01960_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_45_Left_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16760_ net271 _06993_ VGND VGND VPWR VPWR _06994_ sky130_fd_sc_hd__nand2_1
X_13972_ net422 net133 VGND VGND VPWR VPWR _03944_ sky130_fd_sc_hd__nand2_1
X_15711_ net469 net191 net187 net473 VGND VGND VPWR VPWR _05840_ sky130_fd_sc_hd__a22oi_1
X_12923_ _02841_ _02861_ _02859_ VGND VGND VPWR VPWR _02862_ sky130_fd_sc_hd__o21a_1
X_16691_ _06914_ _06917_ VGND VGND VPWR VPWR _06918_ sky130_fd_sc_hd__and2_1
X_18430_ i_error\[8\] _08580_ _08582_ VGND VGND VPWR VPWR _08831_ sky130_fd_sc_hd__nand3_1
X_15642_ _05762_ _05763_ VGND VGND VPWR VPWR _05764_ sky130_fd_sc_hd__and2_1
X_12854_ _02777_ _02792_ VGND VGND VPWR VPWR _02793_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18361_ _08601_ _08752_ net519 VGND VGND VPWR VPWR _08755_ sky130_fd_sc_hd__nand3_4
X_11805_ prev_error\[13\] _08735_ VGND VGND VPWR VPWR _01744_ sky130_fd_sc_hd__nor2_1
X_15573_ _05686_ _05687_ VGND VGND VPWR VPWR _05689_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12785_ _02720_ _02723_ VGND VGND VPWR VPWR _02724_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17312_ _07548_ _07549_ _07600_ VGND VGND VPWR VPWR _07601_ sky130_fd_sc_hd__nor3_4
XFILLER_0_28_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14524_ _04524_ _04532_ _04516_ _04534_ VGND VGND VPWR VPWR _04535_ sky130_fd_sc_hd__o211ai_2
X_11736_ _01671_ _01673_ _01674_ VGND VGND VPWR VPWR _01675_ sky130_fd_sc_hd__a21bo_2
X_18292_ _06750_ _08524_ _06748_ VGND VGND VPWR VPWR _08679_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_54_Left_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17243_ net332 _06334_ _06401_ net315 VGND VGND VPWR VPWR _07526_ sky130_fd_sc_hd__a22oi_2
X_14455_ _04449_ _04455_ _04458_ VGND VGND VPWR VPWR _04459_ sky130_fd_sc_hd__a21oi_1
X_11667_ _01604_ _01605_ VGND VGND VPWR VPWR _01606_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13406_ _03360_ _03361_ VGND VGND VPWR VPWR _03362_ sky130_fd_sc_hd__or2_1
X_17174_ _07115_ _07145_ VGND VGND VPWR VPWR _07450_ sky130_fd_sc_hd__xnor2_1
X_10618_ _00554_ _00556_ VGND VGND VPWR VPWR _00557_ sky130_fd_sc_hd__or2b_1
XFILLER_0_24_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14386_ _04381_ _04375_ _04380_ VGND VGND VPWR VPWR _04383_ sky130_fd_sc_hd__or3_1
X_11598_ _01529_ _01530_ _01534_ VGND VGND VPWR VPWR _01537_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16125_ _01849_ _06290_ _06288_ _06294_ _06295_ VGND VGND VPWR VPWR _06296_ sky130_fd_sc_hd__a221o_1
XFILLER_0_52_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13337_ net233 _02545_ _02640_ net228 VGND VGND VPWR VPWR _03290_ sky130_fd_sc_hd__a22oi_2
X_10549_ net369 _05897_ _06150_ VGND VGND VPWR VPWR _00488_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16056_ _09043_ _06176_ _06219_ VGND VGND VPWR VPWR _06220_ sky130_fd_sc_hd__a21oi_1
X_13268_ net216 _02914_ VGND VGND VPWR VPWR _03221_ sky130_fd_sc_hd__nand2_1
X_15007_ _04944_ _05065_ VGND VGND VPWR VPWR _05066_ sky130_fd_sc_hd__nand2_1
X_12219_ _01984_ _02156_ VGND VGND VPWR VPWR _02158_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13199_ net248 _01874_ VGND VGND VPWR VPWR _03152_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_63_Left_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16958_ net309 _06409_ VGND VGND VPWR VPWR _07212_ sky130_fd_sc_hd__nand2_2
XFILLER_0_154_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15909_ _03862_ _03268_ _03860_ VGND VGND VPWR VPWR _06058_ sky130_fd_sc_hd__nand3_1
X_16889_ _07135_ VGND VGND VPWR VPWR _07136_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18628_ _08837_ VGND VGND VPWR VPWR _09049_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18559_ _06124_ _08972_ VGND VGND VPWR VPWR _08973_ sky130_fd_sc_hd__xnor2_4
XPHY_EDGE_ROW_72_Left_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_12 kp\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_23 net382 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 net357 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09628_ net48 _03091_ _03124_ net122 VGND VGND VPWR VPWR _00027_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12570_ net222 _01874_ _02508_ VGND VGND VPWR VPWR _02509_ sky130_fd_sc_hd__nand3_1
XFILLER_0_65_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11521_ _01431_ _01458_ VGND VGND VPWR VPWR _01460_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14240_ _03899_ _03956_ VGND VGND VPWR VPWR _04222_ sky130_fd_sc_hd__xor2_1
X_11452_ _01388_ _01390_ VGND VGND VPWR VPWR _01391_ sky130_fd_sc_hd__and2_1
XFILLER_0_136_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10403_ _00245_ _00341_ net336 VGND VGND VPWR VPWR _00342_ sky130_fd_sc_hd__and3b_1
XFILLER_0_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14171_ _04144_ _04145_ VGND VGND VPWR VPWR _04146_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11383_ net399 _06612_ _01320_ _01321_ VGND VGND VPWR VPWR _01322_ sky130_fd_sc_hd__a31o_1
X_13122_ _03064_ _03066_ _03067_ VGND VGND VPWR VPWR _03068_ sky130_fd_sc_hd__o21a_1
X_10334_ _00220_ _00272_ VGND VGND VPWR VPWR _00273_ sky130_fd_sc_hd__or2_1
X_13053_ net247 _01852_ VGND VGND VPWR VPWR _02993_ sky130_fd_sc_hd__nand2_1
X_17930_ _08279_ _08280_ VGND VGND VPWR VPWR _08281_ sky130_fd_sc_hd__and2b_1
X_10265_ _00201_ _00203_ VGND VGND VPWR VPWR _00204_ sky130_fd_sc_hd__xnor2_1
X_12004_ _01940_ _01942_ VGND VGND VPWR VPWR _01943_ sky130_fd_sc_hd__nor2_1
X_17861_ _08189_ _08192_ VGND VGND VPWR VPWR _08205_ sky130_fd_sc_hd__nand2_1
X_10196_ net354 _05996_ _08273_ VGND VGND VPWR VPWR _09499_ sky130_fd_sc_hd__and3_1
X_16812_ _07049_ _07050_ _06364_ _06310_ VGND VGND VPWR VPWR _07051_ sky130_fd_sc_hd__a2bb2o_1
X_17792_ _08120_ _08121_ _08128_ VGND VGND VPWR VPWR _08129_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout390 net391 VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__clkbuf_4
X_16743_ net270 _06900_ _06901_ VGND VGND VPWR VPWR _06976_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13955_ net438 net123 net120 net444 VGND VGND VPWR VPWR _03927_ sky130_fd_sc_hd__a22o_1
X_12906_ net224 _02223_ _02737_ _02844_ VGND VGND VPWR VPWR _02845_ sky130_fd_sc_hd__a31o_1
X_16674_ _06800_ VGND VGND VPWR VPWR _06900_ sky130_fd_sc_hd__inv_2
X_13886_ _03427_ _03499_ VGND VGND VPWR VPWR _03852_ sky130_fd_sc_hd__xor2_1
X_18413_ _08808_ net571 _08811_ VGND VGND VPWR VPWR _08813_ sky130_fd_sc_hd__o21a_1
X_15625_ net466 net183 net166 net484 VGND VGND VPWR VPWR _05746_ sky130_fd_sc_hd__a22o_1
X_12837_ _02692_ _02693_ VGND VGND VPWR VPWR _02776_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18344_ _08534_ _08611_ _08736_ VGND VGND VPWR VPWR _08737_ sky130_fd_sc_hd__a21oi_2
X_15556_ _05610_ _05605_ _05608_ VGND VGND VPWR VPWR _05670_ sky130_fd_sc_hd__or3_1
X_12768_ _02702_ _02706_ VGND VGND VPWR VPWR _02707_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14507_ _04494_ _04502_ _04515_ VGND VGND VPWR VPWR _04516_ sky130_fd_sc_hd__a21o_1
XFILLER_0_154_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11719_ _01587_ _01610_ VGND VGND VPWR VPWR _01658_ sky130_fd_sc_hd__and2_1
X_18275_ _06566_ _08660_ VGND VGND VPWR VPWR _08661_ sky130_fd_sc_hd__xor2_1
X_15487_ net437 net197 _05506_ _05507_ VGND VGND VPWR VPWR _05594_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_56_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12699_ _02636_ _02637_ VGND VGND VPWR VPWR _02638_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17226_ net308 _06619_ _06721_ net305 VGND VGND VPWR VPWR _07507_ sky130_fd_sc_hd__a22o_1
Xinput10 measurement[17] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
X_14438_ _04425_ _04427_ _04438_ VGND VGND VPWR VPWR _04440_ sky130_fd_sc_hd__and3_1
Xinput21 reg_addr[0] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_1
XFILLER_0_71_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput32 reg_addr[2] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_1
Xinput43 reg_data[12] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput54 reg_data[5] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_4
X_17157_ _07390_ _07391_ VGND VGND VPWR VPWR _07431_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput65 target[14] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_1
X_14369_ _04361_ _04363_ VGND VGND VPWR VPWR _04364_ sky130_fd_sc_hd__and2_1
Xinput76 target[7] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16108_ prev_error\[2\] _00612_ VGND VGND VPWR VPWR _06277_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17088_ _07123_ _07124_ VGND VGND VPWR VPWR _07355_ sky130_fd_sc_hd__xor2_2
X_16039_ _06920_ _08911_ _06887_ VGND VGND VPWR VPWR _06201_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10050_ net360 _05424_ _07888_ VGND VGND VPWR VPWR _07899_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13740_ net232 _03220_ VGND VGND VPWR VPWR _03706_ sky130_fd_sc_hd__nand2_1
X_10952_ _00886_ _00890_ VGND VGND VPWR VPWR _00891_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13671_ net263 _02222_ _03576_ VGND VGND VPWR VPWR _03634_ sky130_fd_sc_hd__a21oi_1
X_10883_ _00807_ _00821_ VGND VGND VPWR VPWR _00822_ sky130_fd_sc_hd__or2b_1
XFILLER_0_85_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15410_ net437 net193 _05420_ _05421_ VGND VGND VPWR VPWR _05509_ sky130_fd_sc_hd__o2bb2a_1
X_12622_ _02559_ _02560_ VGND VGND VPWR VPWR _02561_ sky130_fd_sc_hd__nand2_1
X_16390_ _06580_ _06586_ _06584_ VGND VGND VPWR VPWR _06587_ sky130_fd_sc_hd__a21oi_1
X_15341_ _05428_ _05432_ VGND VGND VPWR VPWR _05433_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12553_ net254 _01786_ _02427_ VGND VGND VPWR VPWR _02492_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18060_ _08315_ _08314_ _08318_ _08423_ VGND VGND VPWR VPWR _08424_ sky130_fd_sc_hd__o31a_1
X_11504_ _01421_ _01427_ VGND VGND VPWR VPWR _01443_ sky130_fd_sc_hd__xnor2_1
X_15272_ _05344_ _05350_ _05355_ _05356_ VGND VGND VPWR VPWR _05357_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_124_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12484_ _02397_ _02422_ VGND VGND VPWR VPWR _02423_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_108_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17011_ _07267_ _07269_ VGND VGND VPWR VPWR _07270_ sky130_fd_sc_hd__nand2_1
X_14223_ _03916_ _04144_ VGND VGND VPWR VPWR _04204_ sky130_fd_sc_hd__nor2_1
X_11435_ _06590_ _06601_ _00964_ VGND VGND VPWR VPWR _01374_ sky130_fd_sc_hd__a21o_1
XFILLER_0_34_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14154_ net435 _03923_ VGND VGND VPWR VPWR _04128_ sky130_fd_sc_hd__and2_1
X_11366_ _01303_ _01304_ VGND VGND VPWR VPWR _01305_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13105_ _02916_ _02943_ VGND VGND VPWR VPWR _03050_ sky130_fd_sc_hd__xor2_1
X_10317_ _00188_ _00221_ VGND VGND VPWR VPWR _00256_ sky130_fd_sc_hd__xnor2_1
X_14085_ _04024_ _04026_ _04055_ VGND VGND VPWR VPWR _04057_ sky130_fd_sc_hd__or3_1
X_18962_ _09414_ _09415_ VGND VGND VPWR VPWR _09416_ sky130_fd_sc_hd__xor2_1
X_11297_ _01231_ _01232_ _01235_ VGND VGND VPWR VPWR _01236_ sky130_fd_sc_hd__or3_1
X_10248_ _00161_ _00173_ VGND VGND VPWR VPWR _00187_ sky130_fd_sc_hd__xnor2_2
X_13036_ _02865_ _02876_ _02974_ VGND VGND VPWR VPWR _02975_ sky130_fd_sc_hd__nand3_1
X_17913_ _08256_ _08260_ _08261_ VGND VGND VPWR VPWR _08263_ sky130_fd_sc_hd__or3_1
X_18893_ _09278_ _09339_ VGND VGND VPWR VPWR _09341_ sky130_fd_sc_hd__nand2_2
XFILLER_0_28_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17844_ _08070_ _08184_ _08186_ VGND VGND VPWR VPWR _08187_ sky130_fd_sc_hd__and3_1
X_10179_ _09296_ _09307_ VGND VGND VPWR VPWR _09318_ sky130_fd_sc_hd__nor2_1
X_17775_ _07907_ _07999_ _07997_ VGND VGND VPWR VPWR _08111_ sky130_fd_sc_hd__o21a_1
X_14987_ _05041_ _05043_ VGND VGND VPWR VPWR _05044_ sky130_fd_sc_hd__and2b_1
XFILLER_0_44_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16726_ _06947_ _06954_ _06956_ VGND VGND VPWR VPWR _06957_ sky130_fd_sc_hd__a21oi_1
X_13938_ _03907_ _03908_ VGND VGND VPWR VPWR _03909_ sky130_fd_sc_hd__or2_2
X_16657_ _06807_ _06880_ VGND VGND VPWR VPWR _06881_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13869_ _03820_ _03821_ _03829_ _03831_ _03834_ VGND VGND VPWR VPWR _03835_ sky130_fd_sc_hd__a221o_1
XFILLER_0_147_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15608_ _05717_ _05725_ _05726_ VGND VGND VPWR VPWR _05727_ sky130_fd_sc_hd__nand3_1
XFILLER_0_146_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16588_ net278 net274 _06620_ _06723_ VGND VGND VPWR VPWR _06805_ sky130_fd_sc_hd__and4_1
XFILLER_0_29_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18327_ _08627_ _08673_ _08671_ VGND VGND VPWR VPWR _08718_ sky130_fd_sc_hd__a21oi_1
X_15539_ _05641_ _05648_ _05650_ VGND VGND VPWR VPWR _05651_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18258_ _08631_ _08641_ VGND VGND VPWR VPWR _08642_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17209_ _07484_ _07487_ VGND VGND VPWR VPWR _07488_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_53_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18189_ _08556_ _08564_ _08565_ VGND VGND VPWR VPWR _08566_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09962_ net360 VGND VGND VPWR VPWR _06931_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09893_ _06161_ VGND VGND VPWR VPWR _06172_ sky130_fd_sc_hd__buf_6
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclone13 _04170_ _04764_ _05127_ VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__a21o_1
XFILLER_0_90_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11220_ _01153_ _01156_ _01157_ VGND VGND VPWR VPWR _01159_ sky130_fd_sc_hd__nor3_1
X_11151_ net358 _00516_ VGND VGND VPWR VPWR _01090_ sky130_fd_sc_hd__nand2_1
X_10102_ _08075_ _08119_ _08460_ VGND VGND VPWR VPWR _08471_ sky130_fd_sc_hd__a21bo_1
X_11082_ _00996_ _01018_ _01020_ VGND VGND VPWR VPWR _01021_ sky130_fd_sc_hd__o21a_1
X_10033_ _07591_ _07690_ VGND VGND VPWR VPWR _07712_ sky130_fd_sc_hd__nand2_1
X_14910_ net479 net124 _04795_ _04958_ VGND VGND VPWR VPWR _04959_ sky130_fd_sc_hd__o2bb2a_1
X_15890_ _05980_ _04894_ _05967_ VGND VGND VPWR VPWR _06037_ sky130_fd_sc_hd__and3_1
X_14841_ _04881_ _04882_ VGND VGND VPWR VPWR _04883_ sky130_fd_sc_hd__nor2_1
X_17560_ _07655_ _07656_ _07691_ VGND VGND VPWR VPWR _07874_ sky130_fd_sc_hd__o21ai_1
X_14772_ _04805_ _04806_ VGND VGND VPWR VPWR _04807_ sky130_fd_sc_hd__nor2_1
X_11984_ _01894_ _01922_ VGND VGND VPWR VPWR _01923_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16511_ _06718_ _06719_ VGND VGND VPWR VPWR _06720_ sky130_fd_sc_hd__and2_1
X_13723_ _03648_ _03688_ VGND VGND VPWR VPWR _03689_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17491_ _07764_ _07797_ VGND VGND VPWR VPWR _07798_ sky130_fd_sc_hd__xor2_2
X_10935_ _00869_ _00870_ _00873_ VGND VGND VPWR VPWR _00874_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19230_ clknet_4_5_0_clock _00112_ VGND VGND VPWR VPWR prev_error\[17\] sky130_fd_sc_hd__dfxtp_1
X_16442_ _06616_ _06643_ VGND VGND VPWR VPWR _06644_ sky130_fd_sc_hd__or2_1
X_13654_ net247 _02641_ _03613_ _03615_ VGND VGND VPWR VPWR _03616_ sky130_fd_sc_hd__a31o_1
XFILLER_0_155_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10866_ _00712_ _00711_ VGND VGND VPWR VPWR _00805_ sky130_fd_sc_hd__and2b_1
XFILLER_0_156_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12605_ _02543_ VGND VGND VPWR VPWR _02544_ sky130_fd_sc_hd__clkbuf_4
X_19161_ _09559_ _09095_ _09575_ net490 VGND VGND VPWR VPWR _00135_ sky130_fd_sc_hd__o211a_1
X_16373_ _06490_ _06493_ _06565_ VGND VGND VPWR VPWR _06569_ sky130_fd_sc_hd__and3_1
X_13585_ _03484_ _03540_ _03536_ net107 VGND VGND VPWR VPWR _03544_ sky130_fd_sc_hd__a211o_1
XFILLER_0_143_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10797_ _00734_ _00735_ VGND VGND VPWR VPWR _00736_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18112_ _08479_ _08480_ VGND VGND VPWR VPWR _08481_ sky130_fd_sc_hd__xor2_2
X_15324_ _05410_ _05414_ VGND VGND VPWR VPWR _05415_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12536_ _02445_ _02474_ VGND VGND VPWR VPWR _02475_ sky130_fd_sc_hd__or2_1
X_19092_ _09523_ _09583_ _09532_ net489 VGND VGND VPWR VPWR _00102_ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18043_ _08265_ _08300_ VGND VGND VPWR VPWR _08406_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_53_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15255_ net441 net184 net182 net446 VGND VGND VPWR VPWR _05339_ sky130_fd_sc_hd__a22oi_1
X_12467_ _01727_ _01725_ VGND VGND VPWR VPWR _02406_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_34_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_144_Right_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14206_ _04163_ _04184_ VGND VGND VPWR VPWR _04185_ sky130_fd_sc_hd__xnor2_1
X_11418_ _01067_ _01356_ VGND VGND VPWR VPWR _01357_ sky130_fd_sc_hd__xor2_1
XFILLER_0_105_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15186_ _05258_ _05260_ _05262_ VGND VGND VPWR VPWR _05263_ sky130_fd_sc_hd__and3_1
X_12398_ _02321_ _02336_ VGND VGND VPWR VPWR _02337_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14137_ _04107_ _04108_ net408 net138 VGND VGND VPWR VPWR _04109_ sky130_fd_sc_hd__and4b_1
X_11349_ net382 _01285_ _00244_ _01287_ VGND VGND VPWR VPWR _01288_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18945_ _09393_ _09397_ VGND VGND VPWR VPWR _09398_ sky130_fd_sc_hd__xnor2_1
X_14068_ _03980_ _04022_ _04038_ VGND VGND VPWR VPWR _04040_ sky130_fd_sc_hd__nand3_1
X_13019_ _02955_ _02957_ VGND VGND VPWR VPWR _02958_ sky130_fd_sc_hd__and2_1
X_18876_ _01979_ _02157_ _09320_ VGND VGND VPWR VPWR _09322_ sky130_fd_sc_hd__nor3_1
XFILLER_0_146_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17827_ _08050_ _08051_ _08166_ VGND VGND VPWR VPWR _08168_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17758_ _07999_ _08085_ VGND VGND VPWR VPWR _08092_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16709_ net312 _06310_ VGND VGND VPWR VPWR _06938_ sky130_fd_sc_hd__nand2_2
XFILLER_0_77_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17689_ _07930_ _08015_ VGND VGND VPWR VPWR _08016_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_111_Right_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_13_0_clock clknet_0_clock VGND VGND VPWR VPWR clknet_4_13_0_clock sky130_fd_sc_hd__clkbuf_8
XFILLER_0_40_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09945_ _06458_ _06722_ VGND VGND VPWR VPWR _06744_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09876_ _05963_ _05974_ VGND VGND VPWR VPWR _05985_ sky130_fd_sc_hd__and2_1
X_10720_ _00564_ _00658_ VGND VGND VPWR VPWR _00659_ sky130_fd_sc_hd__or2_2
XFILLER_0_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10651_ _00588_ _00589_ VGND VGND VPWR VPWR _00590_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13370_ _03321_ _03320_ _03322_ VGND VGND VPWR VPWR _03323_ sky130_fd_sc_hd__nand3_4
X_10582_ _00512_ _00520_ VGND VGND VPWR VPWR _00521_ sky130_fd_sc_hd__and2b_1
XFILLER_0_35_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12321_ _02177_ _02176_ VGND VGND VPWR VPWR _02260_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15040_ _05100_ _05101_ VGND VGND VPWR VPWR _05102_ sky130_fd_sc_hd__nand2_1
X_12252_ _02189_ _02190_ VGND VGND VPWR VPWR _02191_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11203_ net388 _06623_ _00765_ VGND VGND VPWR VPWR _01142_ sky130_fd_sc_hd__and3_1
X_12183_ _01848_ _01836_ VGND VGND VPWR VPWR _02122_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11134_ _01068_ _01069_ _01072_ VGND VGND VPWR VPWR _01073_ sky130_fd_sc_hd__o21ai_1
X_16991_ _06398_ _07183_ VGND VGND VPWR VPWR _07248_ sky130_fd_sc_hd__or2_1
X_15942_ _06080_ _06093_ VGND VGND VPWR VPWR _06094_ sky130_fd_sc_hd__nand2_1
X_18730_ _06141_ _09159_ _09160_ VGND VGND VPWR VPWR _09161_ sky130_fd_sc_hd__a21o_1
X_11065_ _01002_ _01003_ VGND VGND VPWR VPWR _01004_ sky130_fd_sc_hd__nor2_1
X_10016_ _07393_ _07514_ VGND VGND VPWR VPWR _07525_ sky130_fd_sc_hd__nor2_1
X_18661_ _09082_ _09084_ VGND VGND VPWR VPWR _09085_ sky130_fd_sc_hd__and2_1
X_15873_ _06015_ _06017_ VGND VGND VPWR VPWR _06019_ sky130_fd_sc_hd__nor2_1
X_14824_ _04761_ VGND VGND VPWR VPWR _04865_ sky130_fd_sc_hd__inv_2
X_17612_ net291 _07183_ _07823_ VGND VGND VPWR VPWR _07931_ sky130_fd_sc_hd__a21oi_1
X_18592_ _06170_ _09005_ VGND VGND VPWR VPWR _09009_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17543_ _07853_ _07840_ VGND VGND VPWR VPWR _07856_ sky130_fd_sc_hd__xnor2_2
X_14755_ _04787_ _04788_ VGND VGND VPWR VPWR _04789_ sky130_fd_sc_hd__and2_1
X_11967_ prev_error\[9\] _06612_ VGND VGND VPWR VPWR _01906_ sky130_fd_sc_hd__xor2_4
XFILLER_0_129_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13706_ _03660_ _03671_ VGND VGND VPWR VPWR _03672_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10918_ _00829_ _00855_ VGND VGND VPWR VPWR _00857_ sky130_fd_sc_hd__and2b_1
X_17474_ _07772_ _07779_ VGND VGND VPWR VPWR _07780_ sky130_fd_sc_hd__xnor2_2
X_14686_ _04705_ _04712_ VGND VGND VPWR VPWR _04713_ sky130_fd_sc_hd__or2b_1
X_11898_ net213 _01808_ _01815_ VGND VGND VPWR VPWR _01837_ sky130_fd_sc_hd__and3_1
X_16425_ net275 _06473_ _06470_ _06625_ VGND VGND VPWR VPWR _06626_ sky130_fd_sc_hd__a31o_1
XFILLER_0_55_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19213_ clknet_4_4_0_clock _00095_ VGND VGND VPWR VPWR prev_error\[0\] sky130_fd_sc_hd__dfxtp_2
X_13637_ _03564_ _03570_ _03572_ VGND VGND VPWR VPWR _03597_ sky130_fd_sc_hd__and3_1
X_10849_ _00705_ _00787_ VGND VGND VPWR VPWR _00788_ sky130_fd_sc_hd__or2_1
XFILLER_0_156_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19144_ net504 _09003_ VGND VGND VPWR VPWR _09566_ sky130_fd_sc_hd__nand2_1
X_16356_ net329 net324 net320 _06324_ VGND VGND VPWR VPWR _06550_ sky130_fd_sc_hd__o31a_1
XFILLER_0_41_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13568_ net248 _02410_ _03504_ VGND VGND VPWR VPWR _03527_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15307_ _05393_ _05395_ VGND VGND VPWR VPWR _05396_ sky130_fd_sc_hd__xnor2_1
X_12519_ _02423_ _02457_ _02455_ VGND VGND VPWR VPWR _02458_ sky130_fd_sc_hd__a21o_1
X_19075_ _09515_ _09522_ VGND VGND VPWR VPWR _00094_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16287_ net275 _06404_ _06473_ VGND VGND VPWR VPWR _06474_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13499_ _03457_ VGND VGND VPWR VPWR _03458_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18026_ _08385_ _08386_ VGND VGND VPWR VPWR _08387_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15238_ _05222_ _05319_ VGND VGND VPWR VPWR _05320_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15169_ _05241_ _05242_ _05243_ VGND VGND VPWR VPWR _05244_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_157_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout208 net210 VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__buf_2
Xfanout219 kd_1\[12\] VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__buf_2
XFILLER_0_120_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09730_ _04357_ _04368_ VGND VGND VPWR VPWR _04379_ sky130_fd_sc_hd__nand2_1
X_18928_ _09332_ _09378_ VGND VGND VPWR VPWR _09379_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09661_ _03647_ VGND VGND VPWR VPWR _03658_ sky130_fd_sc_hd__buf_2
X_18859_ _09283_ _09302_ VGND VGND VPWR VPWR _09303_ sky130_fd_sc_hd__xor2_1
XFILLER_0_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09928_ net345 _05897_ _06150_ VGND VGND VPWR VPWR _06557_ sky130_fd_sc_hd__and3_1
X_09859_ _05776_ _05787_ VGND VGND VPWR VPWR _05798_ sky130_fd_sc_hd__nor2_1
X_12870_ _02808_ VGND VGND VPWR VPWR _02809_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11821_ net268 _01759_ VGND VGND VPWR VPWR _01760_ sky130_fd_sc_hd__and2_1
XFILLER_0_96_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14540_ _04536_ _04551_ VGND VGND VPWR VPWR _04552_ sky130_fd_sc_hd__xnor2_1
X_11752_ _00659_ _00757_ VGND VGND VPWR VPWR _01691_ sky130_fd_sc_hd__nand2_1
X_10703_ _00539_ _00637_ _00640_ VGND VGND VPWR VPWR _00642_ sky130_fd_sc_hd__nand3_1
X_14471_ _04470_ _04474_ _04475_ VGND VGND VPWR VPWR _04476_ sky130_fd_sc_hd__o21a_1
XFILLER_0_95_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11683_ net385 _00810_ _00409_ net564 VGND VGND VPWR VPWR _01622_ sky130_fd_sc_hd__a22oi_1
X_16210_ net285 _06307_ _06308_ VGND VGND VPWR VPWR _06389_ sky130_fd_sc_hd__and3_1
XFILLER_0_153_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13422_ _03373_ _03378_ VGND VGND VPWR VPWR _03379_ sky130_fd_sc_hd__or2b_1
XFILLER_0_36_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17190_ net323 _06408_ _06401_ net319 VGND VGND VPWR VPWR _07467_ sky130_fd_sc_hd__a22o_1
X_10634_ net376 _06062_ _00477_ VGND VGND VPWR VPWR _00573_ sky130_fd_sc_hd__and3_1
X_16141_ prev_error\[17\] _04995_ VGND VGND VPWR VPWR _06313_ sky130_fd_sc_hd__nand2_2
X_13353_ _03251_ _03254_ _03253_ VGND VGND VPWR VPWR _03306_ sky130_fd_sc_hd__a21o_1
X_10565_ net352 _09583_ _00398_ VGND VGND VPWR VPWR _00504_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12304_ _02071_ _02208_ _02186_ _02207_ VGND VGND VPWR VPWR _02243_ sky130_fd_sc_hd__o211ai_2
X_16072_ _06181_ _06236_ VGND VGND VPWR VPWR _06237_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13284_ net262 net258 _01851_ _01873_ VGND VGND VPWR VPWR _03237_ sky130_fd_sc_hd__and4_1
XFILLER_0_122_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10496_ _00301_ _00303_ VGND VGND VPWR VPWR _00435_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15023_ _05055_ _05057_ _05082_ VGND VGND VPWR VPWR _05084_ sky130_fd_sc_hd__a21oi_1
X_12235_ _02011_ _02043_ VGND VGND VPWR VPWR _02174_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12166_ _01895_ _02104_ VGND VGND VPWR VPWR _02105_ sky130_fd_sc_hd__xnor2_1
X_11117_ net383 _06634_ VGND VGND VPWR VPWR _01056_ sky130_fd_sc_hd__nand2_1
X_12097_ net234 _01787_ VGND VGND VPWR VPWR _02036_ sky130_fd_sc_hd__nand2_1
X_16974_ _07223_ _07218_ VGND VGND VPWR VPWR _07230_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18713_ _06104_ _06065_ _06103_ VGND VGND VPWR VPWR _09143_ sky130_fd_sc_hd__and3_1
X_15925_ _05948_ _05546_ VGND VGND VPWR VPWR _06076_ sky130_fd_sc_hd__nor2_1
X_11048_ _00935_ _00960_ _00974_ VGND VGND VPWR VPWR _00987_ sky130_fd_sc_hd__a21o_1
Xinput8 measurement[15] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15856_ _04384_ _04476_ VGND VGND VPWR VPWR _06000_ sky130_fd_sc_hd__and2b_1
X_18644_ _09062_ _09066_ VGND VGND VPWR VPWR _09067_ sky130_fd_sc_hd__and2b_1
XFILLER_0_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14807_ _04816_ _04842_ _04844_ VGND VGND VPWR VPWR _04846_ sky130_fd_sc_hd__nand3_1
X_15787_ _05887_ _05907_ _05923_ VGND VGND VPWR VPWR _05924_ sky130_fd_sc_hd__and3_1
X_18575_ _08896_ _08990_ _08964_ VGND VGND VPWR VPWR _08991_ sky130_fd_sc_hd__mux2_1
X_12999_ _02923_ _02925_ VGND VGND VPWR VPWR _02938_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14738_ _04768_ _04759_ _04766_ VGND VGND VPWR VPWR _04770_ sky130_fd_sc_hd__and3_1
X_17526_ _07664_ _07672_ VGND VGND VPWR VPWR _07837_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17457_ _07673_ _07689_ VGND VGND VPWR VPWR _07761_ sky130_fd_sc_hd__nor2_1
X_14669_ _04617_ _04682_ _04686_ VGND VGND VPWR VPWR _04694_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_156_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16408_ _06455_ _06457_ VGND VGND VPWR VPWR _06607_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17388_ _07667_ _07670_ VGND VGND VPWR VPWR _07685_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19127_ _09155_ _09156_ _09550_ VGND VGND VPWR VPWR _09555_ sky130_fd_sc_hd__a21o_1
X_16339_ _06399_ _06404_ _06449_ _06446_ VGND VGND VPWR VPWR _06531_ sky130_fd_sc_hd__o31a_1
XFILLER_0_70_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19058_ _09447_ _09484_ _09451_ VGND VGND VPWR VPWR _09511_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_112_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18009_ _08365_ _08367_ VGND VGND VPWR VPWR _08368_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09713_ net14 net72 VGND VGND VPWR VPWR _04192_ sky130_fd_sc_hd__or2b_2
X_09644_ net57 _03358_ _03391_ net235 VGND VGND VPWR VPWR _00017_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10350_ _00210_ _00208_ VGND VGND VPWR VPWR _00289_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10281_ _00218_ _00219_ VGND VGND VPWR VPWR _00220_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12020_ _01883_ _01958_ VGND VGND VPWR VPWR _01959_ sky130_fd_sc_hd__xor2_1
X_13971_ _03938_ _03942_ VGND VGND VPWR VPWR _03943_ sky130_fd_sc_hd__xnor2_1
X_15710_ net478 net185 VGND VGND VPWR VPWR _05839_ sky130_fd_sc_hd__nand2_1
X_12922_ _02859_ _02860_ VGND VGND VPWR VPWR _02861_ sky130_fd_sc_hd__nand2_1
X_16690_ _06915_ _06916_ VGND VGND VPWR VPWR _06917_ sky130_fd_sc_hd__or2_1
X_15641_ net455 net457 net195 net191 VGND VGND VPWR VPWR _05763_ sky130_fd_sc_hd__and4_1
X_12853_ _02782_ _02791_ _02789_ VGND VGND VPWR VPWR _02792_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_69_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18360_ _08752_ _08753_ _08601_ VGND VGND VPWR VPWR _08754_ sky130_fd_sc_hd__a21o_1
X_11804_ _01742_ VGND VGND VPWR VPWR _01743_ sky130_fd_sc_hd__inv_2
X_15572_ net466 net180 net164 net483 VGND VGND VPWR VPWR _05687_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_29_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12784_ net223 _02091_ _02721_ _02722_ VGND VGND VPWR VPWR _02723_ sky130_fd_sc_hd__a31oi_1
X_17311_ _07577_ _07599_ VGND VGND VPWR VPWR _07600_ sky130_fd_sc_hd__xnor2_1
X_14523_ _04494_ _04502_ _04515_ VGND VGND VPWR VPWR _04534_ sky130_fd_sc_hd__nand3_1
XFILLER_0_68_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11735_ _01411_ _01668_ _01408_ VGND VGND VPWR VPWR _01674_ sky130_fd_sc_hd__or3_1
XFILLER_0_113_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18291_ _08677_ _06668_ VGND VGND VPWR VPWR _08678_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_154_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_1_Left_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17242_ _07521_ _07522_ _07518_ VGND VGND VPWR VPWR _07524_ sky130_fd_sc_hd__a21o_1
X_14454_ _04356_ _04457_ VGND VGND VPWR VPWR _04458_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11666_ _01593_ _01602_ VGND VGND VPWR VPWR _01605_ sky130_fd_sc_hd__xnor2_1
X_13405_ net249 _02223_ _03359_ VGND VGND VPWR VPWR _03361_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17173_ _07434_ _07440_ VGND VGND VPWR VPWR _07449_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10617_ _00497_ _00499_ _00555_ VGND VGND VPWR VPWR _00556_ sky130_fd_sc_hd__a21o_1
X_14385_ _04375_ _04380_ _04381_ VGND VGND VPWR VPWR _04382_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11597_ _01510_ _01511_ VGND VGND VPWR VPWR _01536_ sky130_fd_sc_hd__xor2_1
XFILLER_0_52_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16124_ _01704_ _05930_ VGND VGND VPWR VPWR _06295_ sky130_fd_sc_hd__nor2_1
X_13336_ net225 _02746_ VGND VGND VPWR VPWR _03289_ sky130_fd_sc_hd__nand2_1
X_10548_ net368 _05996_ _06183_ net364 VGND VGND VPWR VPWR _00487_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_11_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16055_ _06217_ _06218_ VGND VGND VPWR VPWR _06219_ sky130_fd_sc_hd__nand2_1
X_13267_ _02935_ VGND VGND VPWR VPWR _03220_ sky130_fd_sc_hd__buf_4
X_10479_ _00405_ _00416_ _00417_ VGND VGND VPWR VPWR _00418_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15006_ _04939_ _04942_ _04943_ VGND VGND VPWR VPWR _05065_ sky130_fd_sc_hd__or3_1
X_12218_ _01984_ _02156_ VGND VGND VPWR VPWR _02157_ sky130_fd_sc_hd__nor2_1
X_13198_ _03149_ _03150_ VGND VGND VPWR VPWR _03151_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12149_ _02085_ _02087_ VGND VGND VPWR VPWR _02088_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_138_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16957_ net302 _06437_ VGND VGND VPWR VPWR _07211_ sky130_fd_sc_hd__nand2_1
X_15908_ _05200_ _05955_ VGND VGND VPWR VPWR _06057_ sky130_fd_sc_hd__xor2_2
X_16888_ _07064_ _07134_ VGND VGND VPWR VPWR _07135_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18627_ _06112_ _09047_ VGND VGND VPWR VPWR _09048_ sky130_fd_sc_hd__nand2_2
X_15839_ _04894_ _05967_ _05980_ VGND VGND VPWR VPWR _05981_ sky130_fd_sc_hd__a21oi_1
X_18558_ _08971_ _06012_ VGND VGND VPWR VPWR _08972_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_63_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17509_ _07574_ _07575_ VGND VGND VPWR VPWR _07818_ sky130_fd_sc_hd__and2_1
XFILLER_0_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18489_ _06173_ _06266_ _08895_ VGND VGND VPWR VPWR _08896_ sky130_fd_sc_hd__nor3_1
XFILLER_0_28_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_13 kp\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_24 net406 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_35 net404 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09627_ net47 _03091_ _03124_ net127 VGND VGND VPWR VPWR _00026_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11520_ _01431_ _01458_ VGND VGND VPWR VPWR _01459_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11451_ _01306_ _01389_ VGND VGND VPWR VPWR _01390_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10402_ _00319_ _00339_ VGND VGND VPWR VPWR _00341_ sky130_fd_sc_hd__xnor2_1
X_14170_ _04127_ _04143_ VGND VGND VPWR VPWR _04145_ sky130_fd_sc_hd__and2_1
X_11382_ net395 _08185_ _01319_ VGND VGND VPWR VPWR _01321_ sky130_fd_sc_hd__and3_1
X_13121_ _03056_ _03061_ _03063_ VGND VGND VPWR VPWR _03067_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10333_ _00218_ _00219_ VGND VGND VPWR VPWR _00272_ sky130_fd_sc_hd__nor2_1
X_13052_ _02989_ _02584_ _02990_ VGND VGND VPWR VPWR _02991_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_131_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10264_ _09395_ _00202_ VGND VGND VPWR VPWR _00203_ sky130_fd_sc_hd__and2_1
X_12003_ net218 _01810_ _01941_ VGND VGND VPWR VPWR _01942_ sky130_fd_sc_hd__and3_1
X_17860_ _08202_ _08203_ VGND VGND VPWR VPWR _08204_ sky130_fd_sc_hd__or2b_1
X_10195_ _08218_ _08251_ VGND VGND VPWR VPWR _09491_ sky130_fd_sc_hd__xnor2_1
X_16811_ net566 _01755_ _06316_ _06309_ net317 VGND VGND VPWR VPWR _07050_ sky130_fd_sc_hd__a32oi_2
X_17791_ _08126_ _08127_ VGND VGND VPWR VPWR _08128_ sky130_fd_sc_hd__or2_1
Xfanout380 kp\[6\] VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_108_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout391 kp\[3\] VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__buf_2
XFILLER_0_89_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16742_ _06957_ _06973_ VGND VGND VPWR VPWR _06974_ sky130_fd_sc_hd__nor2_1
X_13954_ _03922_ _03925_ VGND VGND VPWR VPWR _03926_ sky130_fd_sc_hd__xor2_1
X_12905_ net216 _02409_ _02843_ VGND VGND VPWR VPWR _02844_ sky130_fd_sc_hd__and3_1
X_16673_ _06879_ _06897_ VGND VGND VPWR VPWR _06899_ sky130_fd_sc_hd__and2b_1
X_13885_ _03609_ _03848_ _03850_ VGND VGND VPWR VPWR _03851_ sky130_fd_sc_hd__a21oi_2
X_18412_ _08810_ VGND VGND VPWR VPWR _08811_ sky130_fd_sc_hd__inv_2
X_12836_ _02762_ _02774_ VGND VGND VPWR VPWR _02775_ sky130_fd_sc_hd__nand2_1
X_15624_ net466 net484 net183 net166 VGND VGND VPWR VPWR _05745_ sky130_fd_sc_hd__and4_1
XFILLER_0_57_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15555_ _05616_ _05668_ VGND VGND VPWR VPWR _05669_ sky130_fd_sc_hd__or2_1
X_18343_ _08529_ _08734_ VGND VGND VPWR VPWR _08736_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12767_ _02598_ _02703_ _02705_ VGND VGND VPWR VPWR _02706_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_139_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14506_ _04513_ _04514_ VGND VGND VPWR VPWR _04515_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11718_ _01645_ _01656_ _01612_ _01648_ VGND VGND VPWR VPWR _01657_ sky130_fd_sc_hd__o2bb2a_1
X_18274_ _08656_ _08659_ VGND VGND VPWR VPWR _08660_ sky130_fd_sc_hd__xnor2_1
X_15486_ _05591_ _05592_ VGND VGND VPWR VPWR _05593_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12698_ prev_error\[3\] _00600_ VGND VGND VPWR VPWR _02637_ sky130_fd_sc_hd__xnor2_4
X_14437_ _04425_ _04427_ _04438_ VGND VGND VPWR VPWR _04439_ sky130_fd_sc_hd__a21oi_1
X_17225_ net308 net305 _06619_ _06721_ VGND VGND VPWR VPWR _07506_ sky130_fd_sc_hd__and4_1
Xinput11 measurement[18] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_1
X_11649_ net564 net385 _00815_ _01001_ VGND VGND VPWR VPWR _01588_ sky130_fd_sc_hd__nand4_2
Xinput22 reg_addr[10] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput33 reg_addr[3] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_1
X_17156_ _07405_ _07421_ _07429_ VGND VGND VPWR VPWR _07430_ sky130_fd_sc_hd__a21o_1
Xinput44 reg_data[13] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14368_ _04360_ _04362_ VGND VGND VPWR VPWR _04363_ sky130_fd_sc_hd__nor2_1
Xinput55 reg_data[6] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_4
XFILLER_0_40_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput66 target[15] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput77 target[8] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_1
X_16107_ _02928_ _01717_ _06275_ VGND VGND VPWR VPWR _06276_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13319_ _03259_ _03260_ VGND VGND VPWR VPWR _03272_ sky130_fd_sc_hd__xnor2_1
X_17087_ _07319_ _07328_ VGND VGND VPWR VPWR _07354_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14299_ _04041_ _04042_ _04044_ VGND VGND VPWR VPWR _04287_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16038_ _07382_ _08966_ _08834_ VGND VGND VPWR VPWR _06200_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17989_ _08292_ _08344_ _08338_ _08343_ VGND VGND VPWR VPWR _08346_ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10951_ _00887_ _00781_ _00889_ VGND VGND VPWR VPWR _00890_ sky130_fd_sc_hd__a21oi_1
X_13670_ _03586_ _03632_ VGND VGND VPWR VPWR _03633_ sky130_fd_sc_hd__nor2_1
X_10882_ net337 _00812_ _00817_ _00820_ VGND VGND VPWR VPWR _00821_ sky130_fd_sc_hd__a31o_1
X_12621_ _02473_ _02528_ VGND VGND VPWR VPWR _02560_ sky130_fd_sc_hd__xor2_1
XFILLER_0_156_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_125_Right_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15340_ _05431_ VGND VGND VPWR VPWR _05432_ sky130_fd_sc_hd__inv_2
X_12552_ _02429_ _02432_ VGND VGND VPWR VPWR _02491_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11503_ _01432_ _01441_ VGND VGND VPWR VPWR _01442_ sky130_fd_sc_hd__and2b_1
X_15271_ _05351_ _05352_ _05354_ VGND VGND VPWR VPWR _05356_ sky130_fd_sc_hd__nand3_1
XFILLER_0_151_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12483_ _02418_ _02421_ VGND VGND VPWR VPWR _02422_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_91_Left_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17010_ _07260_ _07268_ VGND VGND VPWR VPWR _07269_ sky130_fd_sc_hd__and2_1
X_14222_ _04200_ _04201_ VGND VGND VPWR VPWR _04202_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11434_ _01357_ _01372_ VGND VGND VPWR VPWR _01373_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14153_ _03921_ VGND VGND VPWR VPWR _04127_ sky130_fd_sc_hd__inv_2
X_11365_ net362 _00814_ _00614_ net366 VGND VGND VPWR VPWR _01304_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_132_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13104_ _03023_ _03048_ VGND VGND VPWR VPWR _03049_ sky130_fd_sc_hd__and2_1
X_10316_ _00225_ _00254_ VGND VGND VPWR VPWR _00255_ sky130_fd_sc_hd__xnor2_1
X_14084_ _04024_ _04026_ _04055_ VGND VGND VPWR VPWR _04056_ sky130_fd_sc_hd__o21ai_2
X_18961_ net408 net130 _09235_ _09234_ VGND VGND VPWR VPWR _09415_ sky130_fd_sc_hd__a31o_1
X_11296_ net358 _00815_ _01234_ VGND VGND VPWR VPWR _01235_ sky130_fd_sc_hd__and3_1
X_13035_ _02945_ _02972_ _02973_ VGND VGND VPWR VPWR _02974_ sky130_fd_sc_hd__a21bo_1
X_17912_ _08201_ _08255_ _08244_ _08254_ VGND VGND VPWR VPWR _08261_ sky130_fd_sc_hd__a211oi_1
X_10247_ _00184_ _00185_ VGND VGND VPWR VPWR _00186_ sky130_fd_sc_hd__and2_2
X_18892_ _09337_ _09338_ VGND VGND VPWR VPWR _09339_ sky130_fd_sc_hd__xnor2_1
X_17843_ _08063_ _08065_ _08068_ _08069_ VGND VGND VPWR VPWR _08186_ sky130_fd_sc_hd__a2bb2o_1
X_10178_ net365 _05424_ _07855_ VGND VGND VPWR VPWR _09307_ sky130_fd_sc_hd__a21oi_1
X_17774_ ki\[8\] _07157_ VGND VGND VPWR VPWR _08110_ sky130_fd_sc_hd__nand2_1
X_14986_ _04915_ _05042_ VGND VGND VPWR VPWR _05043_ sky130_fd_sc_hd__nor2_1
X_16725_ _06870_ _06955_ VGND VGND VPWR VPWR _06956_ sky130_fd_sc_hd__or2_1
X_13937_ _03905_ _03906_ VGND VGND VPWR VPWR _03908_ sky130_fd_sc_hd__and2_1
X_16656_ net286 _06468_ VGND VGND VPWR VPWR _06880_ sky130_fd_sc_hd__nand2_1
X_13868_ _03818_ _03824_ _03833_ VGND VGND VPWR VPWR _03834_ sky130_fd_sc_hd__or3b_1
X_15607_ _05664_ _05724_ _05712_ _05723_ VGND VGND VPWR VPWR _05726_ sky130_fd_sc_hd__o211ai_1
X_12819_ kd_1\[18\] _02748_ _02757_ VGND VGND VPWR VPWR _02758_ sky130_fd_sc_hd__and3_1
X_16587_ net278 _06621_ _06723_ net274 VGND VGND VPWR VPWR _06804_ sky130_fd_sc_hd__a22o_1
X_13799_ _03761_ _03762_ _03764_ VGND VGND VPWR VPWR _03765_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_151_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18326_ _06376_ _08716_ VGND VGND VPWR VPWR _08717_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15538_ _05564_ _05649_ VGND VGND VPWR VPWR _05650_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15469_ _05497_ _05496_ VGND VGND VPWR VPWR _05574_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18257_ _08639_ _08640_ VGND VGND VPWR VPWR _08641_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17208_ _07485_ _07486_ VGND VGND VPWR VPWR _07487_ sky130_fd_sc_hd__xnor2_2
X_18188_ i_error\[2\] _08554_ _08555_ VGND VGND VPWR VPWR _08565_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17139_ _07168_ _07170_ VGND VGND VPWR VPWR _07411_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09961_ _06909_ VGND VGND VPWR VPWR _06920_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09892_ _05897_ _06150_ VGND VGND VPWR VPWR _06161_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_139_Left_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11150_ _01004_ _01088_ VGND VGND VPWR VPWR _01089_ sky130_fd_sc_hd__xor2_1
X_10101_ _08130_ _08394_ VGND VGND VPWR VPWR _08460_ sky130_fd_sc_hd__or2_1
X_11081_ _00899_ _01019_ VGND VGND VPWR VPWR _01020_ sky130_fd_sc_hd__xnor2_1
X_10032_ _07591_ _07690_ VGND VGND VPWR VPWR _07701_ sky130_fd_sc_hd__nor2_1
X_14840_ _04791_ _04853_ VGND VGND VPWR VPWR _04882_ sky130_fd_sc_hd__xnor2_1
X_14771_ _04801_ _04804_ VGND VGND VPWR VPWR _04806_ sky130_fd_sc_hd__nor2_1
X_11983_ _01825_ _01846_ _01893_ VGND VGND VPWR VPWR _01922_ sky130_fd_sc_hd__or3_1
X_13722_ _03645_ _03646_ VGND VGND VPWR VPWR _03688_ sky130_fd_sc_hd__nand2_1
X_16510_ _06273_ _06287_ _02087_ VGND VGND VPWR VPWR _06719_ sky130_fd_sc_hd__a21o_1
X_10934_ _00871_ _00872_ _04841_ _04852_ VGND VGND VPWR VPWR _00873_ sky130_fd_sc_hd__or4bb_4
X_17490_ _07766_ _07796_ VGND VGND VPWR VPWR _07797_ sky130_fd_sc_hd__xor2_2
XFILLER_0_14_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16441_ _06617_ _06640_ _06642_ VGND VGND VPWR VPWR _06643_ sky130_fd_sc_hd__a21oi_2
X_13653_ net269 net251 _02544_ _02089_ VGND VGND VPWR VPWR _03615_ sky130_fd_sc_hd__and4_1
XFILLER_0_129_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10865_ net340 _00614_ VGND VGND VPWR VPWR _00804_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12604_ _02541_ _02542_ VGND VGND VPWR VPWR _02543_ sky130_fd_sc_hd__xor2_4
XFILLER_0_128_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19160_ net501 net477 VGND VGND VPWR VPWR _09575_ sky130_fd_sc_hd__or2_1
X_16372_ _06565_ _06566_ VGND VGND VPWR VPWR _06567_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13584_ _03518_ _03542_ VGND VGND VPWR VPWR _03543_ sky130_fd_sc_hd__xor2_1
XFILLER_0_66_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10796_ _00732_ _00733_ VGND VGND VPWR VPWR _00735_ sky130_fd_sc_hd__xor2_1
XFILLER_0_27_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18111_ _07425_ _07443_ VGND VGND VPWR VPWR _08480_ sky130_fd_sc_hd__xor2_2
X_15323_ _05409_ _05405_ _05407_ VGND VGND VPWR VPWR _05414_ sky130_fd_sc_hd__or3_1
XFILLER_0_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12535_ _02442_ _02444_ VGND VGND VPWR VPWR _02474_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19091_ net499 prev_error\[7\] VGND VGND VPWR VPWR _09532_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15254_ net437 net189 VGND VGND VPWR VPWR _05338_ sky130_fd_sc_hd__nand2_1
X_18042_ _08348_ _08387_ VGND VGND VPWR VPWR _08404_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12466_ _02325_ _02404_ VGND VGND VPWR VPWR _02405_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14205_ _04182_ _04183_ VGND VGND VPWR VPWR _04184_ sky130_fd_sc_hd__and2_1
X_11417_ net385 _00243_ VGND VGND VPWR VPWR _01356_ sky130_fd_sc_hd__and2_1
X_15185_ _05261_ _05240_ VGND VGND VPWR VPWR _05262_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12397_ _02323_ _02335_ VGND VGND VPWR VPWR _02336_ sky130_fd_sc_hd__and2b_1
X_14136_ net415 net134 net130 net419 VGND VGND VPWR VPWR _04108_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11348_ net386 _01286_ _05963_ _05974_ VGND VGND VPWR VPWR _01287_ sky130_fd_sc_hd__and4_1
XFILLER_0_120_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18944_ _09394_ _09396_ VGND VGND VPWR VPWR _09397_ sky130_fd_sc_hd__xnor2_1
X_14067_ _03980_ _04022_ _04038_ VGND VGND VPWR VPWR _04039_ sky130_fd_sc_hd__a21o_1
X_11279_ net370 _00324_ _01146_ VGND VGND VPWR VPWR _01218_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13018_ _02954_ _02950_ _02952_ VGND VGND VPWR VPWR _02957_ sky130_fd_sc_hd__or3_1
X_18875_ _01979_ _02157_ _09320_ VGND VGND VPWR VPWR _09321_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17826_ _08050_ _08051_ _08166_ VGND VGND VPWR VPWR _08167_ sky130_fd_sc_hd__nand3_1
XFILLER_0_89_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17757_ net301 _07182_ VGND VGND VPWR VPWR _08091_ sky130_fd_sc_hd__nand2_1
X_14969_ net472 net474 net144 net138 VGND VGND VPWR VPWR _05024_ sky130_fd_sc_hd__and4_1
X_16708_ _06904_ _06925_ VGND VGND VPWR VPWR _06937_ sky130_fd_sc_hd__xnor2_1
X_17688_ net291 net540 _07929_ VGND VGND VPWR VPWR _08015_ sky130_fd_sc_hd__a21oi_1
X_16639_ net296 _06409_ VGND VGND VPWR VPWR _06861_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18309_ _08694_ _08697_ VGND VGND VPWR VPWR _08698_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19289_ clknet_4_8_0_clock _00038_ VGND VGND VPWR VPWR ki\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_147_Left_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09944_ _06722_ VGND VGND VPWR VPWR _06733_ sky130_fd_sc_hd__inv_2
X_09875_ _05919_ VGND VGND VPWR VPWR _05974_ sky130_fd_sc_hd__buf_2
XFILLER_0_95_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_156_Left_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10650_ _00582_ _00587_ VGND VGND VPWR VPWR _00589_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10581_ _00517_ _00518_ _00519_ VGND VGND VPWR VPWR _00520_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_146_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12320_ _01765_ _02258_ _01762_ VGND VGND VPWR VPWR _02259_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_51_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12251_ _02187_ _02188_ VGND VGND VPWR VPWR _02190_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11202_ _01140_ _00765_ VGND VGND VPWR VPWR _01141_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12182_ _02120_ _02000_ VGND VGND VPWR VPWR _02121_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11133_ _01070_ _01071_ VGND VGND VPWR VPWR _01072_ sky130_fd_sc_hd__xnor2_1
X_16990_ _06398_ _07157_ _07191_ VGND VGND VPWR VPWR _07247_ sky130_fd_sc_hd__o21ba_1
X_15941_ _06077_ _06079_ VGND VGND VPWR VPWR _06093_ sky130_fd_sc_hd__or2_1
X_11064_ net367 _00243_ _00324_ net363 VGND VGND VPWR VPWR _01003_ sky130_fd_sc_hd__a22oi_1
X_10015_ _07426_ _07503_ VGND VGND VPWR VPWR _07514_ sky130_fd_sc_hd__xnor2_1
X_18660_ _06136_ _09082_ _09083_ VGND VGND VPWR VPWR _09084_ sky130_fd_sc_hd__nand3_1
X_15872_ _04382_ _06016_ VGND VGND VPWR VPWR _06017_ sky130_fd_sc_hd__xnor2_1
X_17611_ net291 _07570_ _07929_ VGND VGND VPWR VPWR _07930_ sky130_fd_sc_hd__and3_1
XFILLER_0_99_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14823_ _04860_ _04862_ VGND VGND VPWR VPWR _04864_ sky130_fd_sc_hd__or2_1
X_18591_ _08998_ _09007_ VGND VGND VPWR VPWR _09008_ sky130_fd_sc_hd__xor2_1
X_17542_ _07840_ _07853_ VGND VGND VPWR VPWR _07854_ sky130_fd_sc_hd__or2b_1
X_14754_ _04680_ _04785_ VGND VGND VPWR VPWR _04788_ sky130_fd_sc_hd__nand2_1
X_11966_ _01709_ _01732_ VGND VGND VPWR VPWR _01905_ sky130_fd_sc_hd__nand2_2
XFILLER_0_157_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13705_ _03656_ _03659_ _03657_ VGND VGND VPWR VPWR _03671_ sky130_fd_sc_hd__a21o_1
X_10917_ _00829_ _00855_ VGND VGND VPWR VPWR _00856_ sky130_fd_sc_hd__xnor2_4
X_14685_ _04710_ _04711_ VGND VGND VPWR VPWR _04712_ sky130_fd_sc_hd__and2_1
X_17473_ _07773_ _07777_ VGND VGND VPWR VPWR _07779_ sky130_fd_sc_hd__xor2_2
X_11897_ _01835_ VGND VGND VPWR VPWR _01836_ sky130_fd_sc_hd__clkbuf_4
X_19212_ clknet_4_15_0_clock _00094_ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16424_ net272 _06621_ _06624_ VGND VGND VPWR VPWR _06625_ sky130_fd_sc_hd__and3_1
X_13636_ _03589_ _03594_ _03539_ _03595_ VGND VGND VPWR VPWR _03596_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_39_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10848_ _00702_ _00704_ VGND VGND VPWR VPWR _00787_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19143_ _09559_ _09017_ _09564_ net495 VGND VGND VPWR VPWR _00126_ sky130_fd_sc_hd__o211a_1
X_13567_ _03477_ _03525_ VGND VGND VPWR VPWR _03526_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16355_ _06536_ _06548_ VGND VGND VPWR VPWR _06549_ sky130_fd_sc_hd__or2_2
X_10779_ _00710_ _00716_ _00701_ VGND VGND VPWR VPWR _00718_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12518_ _02455_ _02456_ VGND VGND VPWR VPWR _02457_ sky130_fd_sc_hd__nor2_1
X_15306_ _05327_ _05394_ VGND VGND VPWR VPWR _05395_ sky130_fd_sc_hd__xnor2_1
X_16286_ net278 _06431_ _06434_ VGND VGND VPWR VPWR _06473_ sky130_fd_sc_hd__and3_2
X_19074_ net505 net542 net496 VGND VGND VPWR VPWR _09522_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13498_ _03444_ _03455_ _03456_ VGND VGND VPWR VPWR _03457_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_140_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18025_ _08351_ _08371_ VGND VGND VPWR VPWR _08386_ sky130_fd_sc_hd__xnor2_1
X_12449_ _02319_ _02387_ VGND VGND VPWR VPWR _02388_ sky130_fd_sc_hd__nor2_1
X_15237_ _05219_ _05221_ VGND VGND VPWR VPWR _05319_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15168_ net441 net446 net181 net177 VGND VGND VPWR VPWR _05243_ sky130_fd_sc_hd__and4_1
X_14119_ _03921_ _03953_ _03916_ VGND VGND VPWR VPWR _04091_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout209 net210 VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_2
X_15099_ _05062_ _05166_ VGND VGND VPWR VPWR _05167_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18927_ _09368_ _09377_ VGND VGND VPWR VPWR _09378_ sky130_fd_sc_hd__xnor2_1
X_09660_ _03636_ VGND VGND VPWR VPWR _03647_ sky130_fd_sc_hd__clkbuf_4
X_18858_ _09284_ _09301_ VGND VGND VPWR VPWR _09302_ sky130_fd_sc_hd__xnor2_1
X_17809_ _08139_ _08140_ VGND VGND VPWR VPWR _08148_ sky130_fd_sc_hd__nand2_1
X_18789_ _04161_ _04211_ VGND VGND VPWR VPWR _09226_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09927_ _06535_ VGND VGND VPWR VPWR _06546_ sky130_fd_sc_hd__inv_2
X_09858_ net356 net353 _05182_ _04885_ VGND VGND VPWR VPWR _05787_ sky130_fd_sc_hd__and4_1
X_09789_ net69 net11 VGND VGND VPWR VPWR _05028_ sky130_fd_sc_hd__xnor2_1
X_11820_ _01754_ _01757_ _05600_ _01758_ VGND VGND VPWR VPWR _01759_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_139_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11751_ _00866_ _00959_ net569 _01689_ _00865_ VGND VGND VPWR VPWR _01690_ sky130_fd_sc_hd__a32o_2
XFILLER_0_96_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10702_ _00539_ _00637_ _00640_ VGND VGND VPWR VPWR _00641_ sky130_fd_sc_hd__a21o_1
X_14470_ _04378_ _04377_ VGND VGND VPWR VPWR _04475_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11682_ net399 _00614_ _01620_ _01618_ VGND VGND VPWR VPWR _01621_ sky130_fd_sc_hd__a31o_1
XFILLER_0_83_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13421_ _03376_ _03377_ VGND VGND VPWR VPWR _03378_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10633_ net376 _06062_ _00477_ VGND VGND VPWR VPWR _00572_ sky130_fd_sc_hd__a21o_1
XFILLER_0_107_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16140_ ki\[11\] _06311_ VGND VGND VPWR VPWR _06312_ sky130_fd_sc_hd__nand2_1
X_13352_ _03303_ _03304_ VGND VGND VPWR VPWR _03305_ sky130_fd_sc_hd__nor2_1
X_10564_ net565 _09558_ _09565_ VGND VGND VPWR VPWR _00503_ sky130_fd_sc_hd__and3_2
XFILLER_0_107_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12303_ _02240_ _02241_ VGND VGND VPWR VPWR _02242_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16071_ _06179_ _06189_ _06187_ VGND VGND VPWR VPWR _06236_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13283_ _03234_ _03235_ VGND VGND VPWR VPWR _03236_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_121_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10495_ _00373_ _00372_ VGND VGND VPWR VPWR _00434_ sky130_fd_sc_hd__xnor2_2
X_15022_ _04948_ _04950_ VGND VGND VPWR VPWR _05082_ sky130_fd_sc_hd__xnor2_1
X_12234_ _02171_ _02172_ VGND VGND VPWR VPWR _02173_ sky130_fd_sc_hd__nand2_1
X_12165_ _01920_ _01919_ VGND VGND VPWR VPWR _02104_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11116_ _01053_ _01054_ VGND VGND VPWR VPWR _01055_ sky130_fd_sc_hd__xnor2_1
X_12096_ _02013_ _02034_ VGND VGND VPWR VPWR _02035_ sky130_fd_sc_hd__or2_1
X_16973_ net305 _06438_ _07225_ _07227_ VGND VGND VPWR VPWR _07229_ sky130_fd_sc_hd__a31o_1
X_18712_ _06065_ _06103_ _06104_ VGND VGND VPWR VPWR _09141_ sky130_fd_sc_hd__a21oi_1
X_15924_ _06072_ _06074_ VGND VGND VPWR VPWR _06075_ sky130_fd_sc_hd__nand2_1
X_11047_ _00981_ _00985_ VGND VGND VPWR VPWR _00986_ sky130_fd_sc_hd__xnor2_2
Xinput9 measurement[16] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
X_18643_ _08912_ _09064_ _08963_ VGND VGND VPWR VPWR _09066_ sky130_fd_sc_hd__mux2_1
X_15855_ _04304_ _05998_ VGND VGND VPWR VPWR _05999_ sky130_fd_sc_hd__or2_1
X_14806_ _04816_ _04842_ _04844_ VGND VGND VPWR VPWR _04845_ sky130_fd_sc_hd__a21o_1
X_18574_ _08989_ _08748_ _08882_ VGND VGND VPWR VPWR _08990_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15786_ _05903_ _05918_ _05915_ _05922_ VGND VGND VPWR VPWR _05923_ sky130_fd_sc_hd__and4b_1
X_12998_ net202 _02935_ _02927_ _02936_ VGND VGND VPWR VPWR _02937_ sky130_fd_sc_hd__nand4_1
XFILLER_0_143_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17525_ _07832_ _07835_ VGND VGND VPWR VPWR _07836_ sky130_fd_sc_hd__nand2_1
X_14737_ _04759_ _04766_ _04768_ VGND VGND VPWR VPWR _04769_ sky130_fd_sc_hd__a21oi_1
X_11949_ _01881_ _01887_ VGND VGND VPWR VPWR _01888_ sky130_fd_sc_hd__xor2_1
XFILLER_0_52_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17456_ _07655_ net537 _07758_ _07759_ VGND VGND VPWR VPWR _07760_ sky130_fd_sc_hd__o211ai_4
X_14668_ _04691_ _04692_ VGND VGND VPWR VPWR _04693_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16407_ _06604_ _06605_ VGND VGND VPWR VPWR _06606_ sky130_fd_sc_hd__nor2_1
X_13619_ net265 _02090_ _03530_ _03531_ VGND VGND VPWR VPWR _03578_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17387_ _07682_ _07683_ VGND VGND VPWR VPWR _07684_ sky130_fd_sc_hd__nand2_1
X_14599_ _03917_ _04614_ _04616_ VGND VGND VPWR VPWR _04617_ sky130_fd_sc_hd__nor3_1
XFILLER_0_144_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19126_ net506 net561 net494 _09554_ VGND VGND VPWR VPWR _00118_ sky130_fd_sc_hd__o211a_1
X_16338_ _06506_ _06529_ VGND VGND VPWR VPWR _06530_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19057_ _04126_ net82 VGND VGND VPWR VPWR _09510_ sky130_fd_sc_hd__and2_1
X_16269_ _06354_ _06453_ VGND VGND VPWR VPWR _06454_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18008_ _08335_ _08366_ VGND VGND VPWR VPWR _08367_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09712_ net5 net63 VGND VGND VPWR VPWR _04181_ sky130_fd_sc_hd__or2b_2
X_09643_ net56 _03358_ _03391_ net241 VGND VGND VPWR VPWR _00016_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10280_ _00189_ _00198_ VGND VGND VPWR VPWR _00219_ sky130_fd_sc_hd__xnor2_1
X_13970_ _03939_ _03941_ VGND VGND VPWR VPWR _03942_ sky130_fd_sc_hd__xnor2_1
X_12921_ _02858_ _02849_ _02856_ VGND VGND VPWR VPWR _02860_ sky130_fd_sc_hd__nand3_1
X_15640_ _05760_ _05761_ VGND VGND VPWR VPWR _05762_ sky130_fd_sc_hd__nor2_1
X_12852_ _02789_ _02790_ VGND VGND VPWR VPWR _02791_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11803_ _01740_ _01741_ VGND VGND VPWR VPWR _01742_ sky130_fd_sc_hd__nor2_8
X_15571_ net466 net483 net180 net164 VGND VGND VPWR VPWR _05686_ sky130_fd_sc_hd__and4_1
X_12783_ net227 _01909_ _02615_ VGND VGND VPWR VPWR _02722_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17310_ _07597_ _07598_ VGND VGND VPWR VPWR _07599_ sky130_fd_sc_hd__nor2_1
X_14522_ _04526_ _04531_ VGND VGND VPWR VPWR _04532_ sky130_fd_sc_hd__and2_1
X_11734_ _01408_ _01672_ VGND VGND VPWR VPWR _01673_ sky130_fd_sc_hd__xnor2_4
X_18290_ _08675_ _08676_ VGND VGND VPWR VPWR _08677_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17241_ _07518_ _07521_ _07522_ VGND VGND VPWR VPWR _07523_ sky130_fd_sc_hd__nand3_1
X_14453_ _04351_ _04353_ _04355_ VGND VGND VPWR VPWR _04457_ sky130_fd_sc_hd__or3_1
X_11665_ _01591_ _01603_ VGND VGND VPWR VPWR _01604_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13404_ net249 _02223_ _03359_ VGND VGND VPWR VPWR _03360_ sky130_fd_sc_hd__and3_1
X_10616_ _00500_ _00526_ VGND VGND VPWR VPWR _00555_ sky130_fd_sc_hd__nor2_1
X_17172_ _07432_ _07433_ VGND VGND VPWR VPWR _07447_ sky130_fd_sc_hd__nand2_1
X_14384_ _04293_ _04292_ VGND VGND VPWR VPWR _04381_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11596_ _01529_ _01530_ _01534_ VGND VGND VPWR VPWR _01535_ sky130_fd_sc_hd__nand3_1
XFILLER_0_51_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13335_ _03207_ _03210_ VGND VGND VPWR VPWR _03288_ sky130_fd_sc_hd__xor2_1
X_16123_ net115 _06291_ _06292_ VGND VGND VPWR VPWR _06294_ sky130_fd_sc_hd__a21o_1
X_10547_ net361 _06634_ VGND VGND VPWR VPWR _00486_ sky130_fd_sc_hd__nand2_1
X_16054_ _06215_ _06214_ VGND VGND VPWR VPWR _06218_ sky130_fd_sc_hd__or2b_1
X_13266_ _03216_ _03218_ VGND VGND VPWR VPWR _03219_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10478_ _00328_ _00338_ VGND VGND VPWR VPWR _00417_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12217_ _02147_ _02155_ VGND VGND VPWR VPWR _02156_ sky130_fd_sc_hd__xnor2_1
X_15005_ _04985_ _05003_ _05063_ VGND VGND VPWR VPWR _05064_ sky130_fd_sc_hd__or3_2
X_13197_ _03148_ _03145_ VGND VGND VPWR VPWR _03150_ sky130_fd_sc_hd__and2b_1
X_12148_ _02086_ _01731_ VGND VGND VPWR VPWR _02087_ sky130_fd_sc_hd__or2_4
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12079_ _02015_ _02017_ VGND VGND VPWR VPWR _02018_ sky130_fd_sc_hd__nand2_1
X_16956_ _07200_ _07204_ _07209_ VGND VGND VPWR VPWR _07210_ sky130_fd_sc_hd__o21ai_4
X_15907_ _06053_ _06055_ VGND VGND VPWR VPWR _06056_ sky130_fd_sc_hd__nand2_1
X_16887_ _07061_ _07062_ VGND VGND VPWR VPWR _07134_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_139_Right_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18626_ _06111_ _06050_ _06110_ VGND VGND VPWR VPWR _09047_ sky130_fd_sc_hd__nand3_1
XFILLER_0_2_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15838_ _05978_ _05979_ VGND VGND VPWR VPWR _05980_ sky130_fd_sc_hd__nand2_1
X_18557_ _06009_ _06010_ VGND VGND VPWR VPWR _08971_ sky130_fd_sc_hd__nand2_1
X_15769_ _05896_ _05900_ _05903_ VGND VGND VPWR VPWR _05904_ sky130_fd_sc_hd__a21o_1
X_17508_ _07815_ _07816_ VGND VGND VPWR VPWR _07817_ sky130_fd_sc_hd__nand2_1
X_18488_ _06169_ _06170_ _06133_ VGND VGND VPWR VPWR _08895_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_111_Left_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_14 kp\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17439_ _07263_ _07265_ VGND VGND VPWR VPWR _07741_ sky130_fd_sc_hd__nand2_1
XANTENNA_25 net406 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_36 net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19109_ _09536_ _05193_ _09543_ net488 VGND VGND VPWR VPWR _00110_ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_120_Left_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_106_Right_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09626_ net46 _03091_ _03124_ net132 VGND VGND VPWR VPWR _00025_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11450_ net358 _00811_ _01305_ VGND VGND VPWR VPWR _01389_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_151_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10401_ _00339_ VGND VGND VPWR VPWR _00340_ sky130_fd_sc_hd__inv_2
X_11381_ _01257_ _01319_ VGND VGND VPWR VPWR _01320_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13120_ _02225_ _03065_ _02926_ VGND VGND VPWR VPWR _03066_ sky130_fd_sc_hd__or3_1
XFILLER_0_61_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10332_ _00257_ _00270_ VGND VGND VPWR VPWR _00271_ sky130_fd_sc_hd__or2_1
X_13051_ net251 _01859_ _01797_ net267 VGND VGND VPWR VPWR _02990_ sky130_fd_sc_hd__a22o_1
X_10263_ _09362_ _09384_ VGND VGND VPWR VPWR _00202_ sky130_fd_sc_hd__nand2_1
X_12002_ net215 _01787_ VGND VGND VPWR VPWR _01941_ sky130_fd_sc_hd__and2_1
X_10194_ _08097_ _08207_ VGND VGND VPWR VPWR _09483_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16810_ net312 _06335_ VGND VGND VPWR VPWR _07049_ sky130_fd_sc_hd__nand2_1
X_17790_ _08124_ _08125_ VGND VGND VPWR VPWR _08127_ sky130_fd_sc_hd__nor2_1
Xfanout370 net373 VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__clkbuf_4
Xfanout381 net382 VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__clkbuf_4
X_16741_ _06970_ _06972_ VGND VGND VPWR VPWR _06973_ sky130_fd_sc_hd__and2b_1
Xfanout392 kp\[3\] VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__clkbuf_4
X_13953_ net119 _03923_ _03924_ VGND VGND VPWR VPWR _03925_ sky130_fd_sc_hd__a21bo_1
X_12904_ _02737_ _02842_ VGND VGND VPWR VPWR _02843_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16672_ _06883_ _06886_ _06896_ VGND VGND VPWR VPWR _06897_ sky130_fd_sc_hd__a21bo_1
X_13884_ _03553_ _03849_ VGND VGND VPWR VPWR _03850_ sky130_fd_sc_hd__or2_1
X_18411_ _08809_ _08566_ VGND VGND VPWR VPWR _08810_ sky130_fd_sc_hd__xor2_2
X_15623_ _05738_ _05740_ _05742_ VGND VGND VPWR VPWR _05744_ sky130_fd_sc_hd__o21ai_1
X_12835_ _02760_ _02761_ VGND VGND VPWR VPWR _02774_ sky130_fd_sc_hd__or2_1
X_18342_ i_error\[15\] _08528_ VGND VGND VPWR VPWR _08734_ sky130_fd_sc_hd__or2_1
X_15554_ _05634_ _05665_ _05667_ VGND VGND VPWR VPWR _05668_ sky130_fd_sc_hd__a21boi_1
X_12766_ net235 _01853_ _02704_ VGND VGND VPWR VPWR _02705_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14505_ _04509_ _04512_ VGND VGND VPWR VPWR _04514_ sky130_fd_sc_hd__nor2_1
X_11717_ _01634_ _01646_ _01652_ _01654_ _01655_ VGND VGND VPWR VPWR _01656_ sky130_fd_sc_hd__o221a_1
X_18273_ _06561_ _08657_ _06328_ VGND VGND VPWR VPWR _08659_ sky130_fd_sc_hd__and3b_1
X_15485_ _05587_ _05577_ _05590_ VGND VGND VPWR VPWR _05592_ sky130_fd_sc_hd__nor3_1
X_12697_ _01715_ _01719_ _01720_ VGND VGND VPWR VPWR _02636_ sky130_fd_sc_hd__a21o_1
X_17224_ _07489_ _07494_ _07491_ VGND VGND VPWR VPWR _07505_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_154_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14436_ _04361_ _04363_ VGND VGND VPWR VPWR _04438_ sky130_fd_sc_hd__xnor2_1
X_11648_ _01576_ _01586_ VGND VGND VPWR VPWR _01587_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput12 measurement[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_6
Xinput23 reg_addr[11] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput34 reg_addr[4] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17155_ _07388_ _07403_ VGND VGND VPWR VPWR _07429_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput45 reg_data[14] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14367_ _04359_ _04350_ _04356_ VGND VGND VPWR VPWR _04362_ sky130_fd_sc_hd__and3_1
X_11579_ net377 _00810_ VGND VGND VPWR VPWR _01518_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput56 reg_data[7] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_4
Xinput67 target[16] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16106_ prev_error\[1\] _00813_ VGND VGND VPWR VPWR _06275_ sky130_fd_sc_hd__nand2_1
Xinput78 target[9] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13318_ _03230_ _03265_ VGND VGND VPWR VPWR _03271_ sky130_fd_sc_hd__xnor2_1
X_17086_ _07333_ _07343_ _07332_ VGND VGND VPWR VPWR _07353_ sky130_fd_sc_hd__a21bo_1
X_14298_ _04282_ _04283_ _04285_ VGND VGND VPWR VPWR _04286_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16037_ _06196_ _06197_ VGND VGND VPWR VPWR _06199_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13249_ net212 _02915_ _03132_ VGND VGND VPWR VPWR _03202_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17988_ _08338_ _08343_ _08292_ _08344_ VGND VGND VPWR VPWR _08345_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_74_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16939_ _07172_ _07190_ VGND VGND VPWR VPWR _07191_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18609_ _09026_ _09027_ _08964_ VGND VGND VPWR VPWR _09028_ sky130_fd_sc_hd__mux2_2
XFILLER_0_87_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10950_ net359 _00324_ _00888_ VGND VGND VPWR VPWR _00889_ sky130_fd_sc_hd__and3_1
XFILLER_0_86_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09609_ _03113_ VGND VGND VPWR VPWR _03124_ sky130_fd_sc_hd__clkbuf_4
X_10881_ _00804_ _00819_ VGND VGND VPWR VPWR _00820_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12620_ _02532_ _02558_ VGND VGND VPWR VPWR _02559_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12551_ _02488_ _02489_ VGND VGND VPWR VPWR _02490_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11502_ _01437_ _01440_ VGND VGND VPWR VPWR _01441_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12482_ net199 _02419_ _02420_ VGND VGND VPWR VPWR _02421_ sky130_fd_sc_hd__and3_1
X_15270_ _05351_ _05352_ _05354_ VGND VGND VPWR VPWR _05355_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14221_ _04127_ _04199_ VGND VGND VPWR VPWR _04201_ sky130_fd_sc_hd__and2_1
X_11433_ net381 _00324_ VGND VGND VPWR VPWR _01372_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14152_ _04122_ _04123_ _04059_ _04062_ VGND VGND VPWR VPWR _04125_ sky130_fd_sc_hd__a211oi_1
X_11364_ net366 net362 _00814_ _00613_ VGND VGND VPWR VPWR _01303_ sky130_fd_sc_hd__and4_1
XFILLER_0_10_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13103_ _03023_ _03045_ _03046_ VGND VGND VPWR VPWR _03048_ sky130_fd_sc_hd__nand3_1
XFILLER_0_104_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10315_ _00227_ _00252_ _00253_ VGND VGND VPWR VPWR _00254_ sky130_fd_sc_hd__o21ba_1
X_14083_ _04048_ _04054_ VGND VGND VPWR VPWR _04055_ sky130_fd_sc_hd__xnor2_1
X_18960_ _04138_ _09253_ _04128_ VGND VGND VPWR VPWR _09414_ sky130_fd_sc_hd__o21ba_1
X_11295_ _01232_ _01233_ VGND VGND VPWR VPWR _01234_ sky130_fd_sc_hd__nor2_1
X_13034_ _02967_ _02971_ _02833_ _02946_ VGND VGND VPWR VPWR _02973_ sky130_fd_sc_hd__a211o_1
X_17911_ _08257_ _08259_ VGND VGND VPWR VPWR _08260_ sky130_fd_sc_hd__xor2_1
X_10246_ _00182_ _00183_ VGND VGND VPWR VPWR _00185_ sky130_fd_sc_hd__or2_1
X_18891_ _02173_ _03890_ _02171_ VGND VGND VPWR VPWR _09338_ sky130_fd_sc_hd__o21a_1
X_17842_ _08173_ _08182_ _08183_ VGND VGND VPWR VPWR _08184_ sky130_fd_sc_hd__a21o_1
X_10177_ net365 _05424_ _07855_ VGND VGND VPWR VPWR _09296_ sky130_fd_sc_hd__and3_1
X_17773_ _07493_ _08107_ _08079_ _08077_ VGND VGND VPWR VPWR _08109_ sky130_fd_sc_hd__o22ai_2
X_14985_ net436 net173 _04913_ _04914_ VGND VGND VPWR VPWR _05042_ sky130_fd_sc_hd__o2bb2a_1
X_16724_ _06867_ _06869_ VGND VGND VPWR VPWR _06955_ sky130_fd_sc_hd__and2_1
X_13936_ _03905_ _03906_ VGND VGND VPWR VPWR _03907_ sky130_fd_sc_hd__nor2_2
XFILLER_0_88_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16655_ _06806_ _06816_ VGND VGND VPWR VPWR _06879_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13867_ _03828_ _03832_ _03791_ VGND VGND VPWR VPWR _03833_ sky130_fd_sc_hd__and3b_1
X_15606_ _05712_ _05723_ _05664_ _05724_ VGND VGND VPWR VPWR _05725_ sky130_fd_sc_hd__a211o_1
X_12818_ _02736_ _02755_ VGND VGND VPWR VPWR _02757_ sky130_fd_sc_hd__xnor2_1
X_16586_ _06802_ VGND VGND VPWR VPWR _06803_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13798_ net263 _02639_ _03763_ VGND VGND VPWR VPWR _03764_ sky130_fd_sc_hd__and3_1
X_18325_ _06554_ _08665_ _06549_ VGND VGND VPWR VPWR _08716_ sky130_fd_sc_hd__a21bo_1
X_15537_ _05561_ _05563_ VGND VGND VPWR VPWR _05649_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12749_ _02687_ VGND VGND VPWR VPWR _02688_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18256_ _08632_ _08638_ VGND VGND VPWR VPWR _08640_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15468_ net463 net176 _05559_ _05558_ VGND VGND VPWR VPWR _05573_ sky130_fd_sc_hd__a31oi_2
X_17207_ _07474_ _07472_ VGND VGND VPWR VPWR _07486_ sky130_fd_sc_hd__and2b_1
X_14419_ net420 net156 _04344_ _04345_ VGND VGND VPWR VPWR _04419_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_114_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18187_ _08560_ _08562_ _08563_ VGND VGND VPWR VPWR _08564_ sky130_fd_sc_hd__a21o_1
XFILLER_0_108_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15399_ net453 net458 net181 net177 VGND VGND VPWR VPWR _05497_ sky130_fd_sc_hd__and4_1
XFILLER_0_52_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17138_ _06398_ _07095_ VGND VGND VPWR VPWR _07410_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09960_ _06887_ _06898_ _05600_ VGND VGND VPWR VPWR _06909_ sky130_fd_sc_hd__and3b_1
X_17069_ net302 _06438_ _07215_ _07214_ VGND VGND VPWR VPWR _07334_ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09891_ _04599_ _04665_ _05886_ VGND VGND VPWR VPWR _06150_ sky130_fd_sc_hd__nand3_2
XFILLER_0_110_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclone15 _09447_ VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__buf_6
XFILLER_0_146_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10100_ _07756_ _08438_ VGND VGND VPWR VPWR _08449_ sky130_fd_sc_hd__xnor2_1
X_11080_ _00916_ _00915_ VGND VGND VPWR VPWR _01019_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10031_ _07613_ _07679_ _07657_ VGND VGND VPWR VPWR _07690_ sky130_fd_sc_hd__a21oi_1
X_14770_ _04801_ _04804_ VGND VGND VPWR VPWR _04805_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11982_ _01895_ _01919_ _01920_ VGND VGND VPWR VPWR _01921_ sky130_fd_sc_hd__o21ba_1
X_13721_ _03684_ _03686_ VGND VGND VPWR VPWR _03687_ sky130_fd_sc_hd__and2_1
X_10933_ net387 _06062_ VGND VGND VPWR VPWR _00872_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16440_ _06470_ _06641_ ki\[18\] VGND VGND VPWR VPWR _06642_ sky130_fd_sc_hd__and3b_1
X_13652_ _03611_ _02210_ _03612_ VGND VGND VPWR VPWR _03613_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_85_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10864_ _00799_ _00802_ VGND VGND VPWR VPWR _00803_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12603_ _01713_ _01721_ VGND VGND VPWR VPWR _02542_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16371_ _06490_ _06493_ VGND VGND VPWR VPWR _06566_ sky130_fd_sc_hd__and2_1
XFILLER_0_155_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13583_ _03521_ _03522_ VGND VGND VPWR VPWR _03542_ sky130_fd_sc_hd__and2_1
X_10795_ net401 _04841_ _04852_ VGND VGND VPWR VPWR _00734_ sky130_fd_sc_hd__and3_1
X_18110_ _08464_ _08463_ VGND VGND VPWR VPWR _08479_ sky130_fd_sc_hd__and2b_1
X_15322_ _05411_ _05390_ VGND VGND VPWR VPWR _05412_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12534_ _02452_ _02472_ VGND VGND VPWR VPWR _02473_ sky130_fd_sc_hd__nand2_1
X_19090_ _09523_ _00245_ _09531_ net489 VGND VGND VPWR VPWR _00101_ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18041_ _08348_ _08373_ _08387_ _08402_ VGND VGND VPWR VPWR _08403_ sky130_fd_sc_hd__a31o_1
X_15253_ _05335_ _05334_ VGND VGND VPWR VPWR _05337_ sky130_fd_sc_hd__xnor2_1
X_12465_ net206 _02332_ VGND VGND VPWR VPWR _02404_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14204_ _04017_ net140 _04180_ VGND VGND VPWR VPWR _04183_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11416_ _01333_ _01334_ VGND VGND VPWR VPWR _01355_ sky130_fd_sc_hd__xnor2_1
X_12396_ _02324_ _02325_ _02334_ VGND VGND VPWR VPWR _02335_ sky130_fd_sc_hd__o21ai_1
X_15184_ _05135_ _05207_ VGND VGND VPWR VPWR _05261_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14135_ net415 net418 net134 net130 VGND VGND VPWR VPWR _04107_ sky130_fd_sc_hd__and4_1
X_11347_ net564 _09558_ _09565_ VGND VGND VPWR VPWR _01286_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18943_ net210 _01772_ VGND VGND VPWR VPWR _09396_ sky130_fd_sc_hd__nand2_1
X_14066_ _04023_ _04037_ VGND VGND VPWR VPWR _04038_ sky130_fd_sc_hd__xnor2_1
X_11278_ net381 _09577_ _01215_ _01216_ VGND VGND VPWR VPWR _01217_ sky130_fd_sc_hd__a31o_1
X_10229_ _00165_ _00167_ VGND VGND VPWR VPWR _00168_ sky130_fd_sc_hd__and2_1
X_13017_ _02799_ _02882_ VGND VGND VPWR VPWR _02956_ sky130_fd_sc_hd__xnor2_2
X_18874_ _01984_ _09319_ VGND VGND VPWR VPWR _09320_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17825_ _08158_ _08162_ _08165_ VGND VGND VPWR VPWR _08166_ sky130_fd_sc_hd__o21a_1
XFILLER_0_146_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17756_ _08067_ _08068_ VGND VGND VPWR VPWR _08090_ sky130_fd_sc_hd__nand2_1
X_14968_ net478 net135 VGND VGND VPWR VPWR _05023_ sky130_fd_sc_hd__nand2_1
X_16707_ _06929_ _06927_ VGND VGND VPWR VPWR _06936_ sky130_fd_sc_hd__xor2_2
X_13919_ _02252_ _02254_ VGND VGND VPWR VPWR _03888_ sky130_fd_sc_hd__xnor2_1
X_17687_ _07919_ _08012_ _08011_ _07995_ VGND VGND VPWR VPWR _08014_ sky130_fd_sc_hd__a211oi_2
X_14899_ _04938_ _04944_ _04946_ VGND VGND VPWR VPWR _04947_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_76_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16638_ _06858_ _06859_ VGND VGND VPWR VPWR _06860_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_147_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16569_ _06649_ _06698_ VGND VGND VPWR VPWR _06784_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18308_ _08695_ _08696_ VGND VGND VPWR VPWR _08697_ sky130_fd_sc_hd__xnor2_1
X_19288_ clknet_4_6_0_clock _00066_ VGND VGND VPWR VPWR kp\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18239_ _01698_ _08617_ VGND VGND VPWR VPWR _08621_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09943_ _06513_ _06546_ _06711_ VGND VGND VPWR VPWR _06722_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09874_ _05908_ VGND VGND VPWR VPWR _05963_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10580_ kp\[15\] net340 _00410_ _00325_ VGND VGND VPWR VPWR _00519_ sky130_fd_sc_hd__nand4_1
XFILLER_0_51_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_7_0_clock clknet_0_clock VGND VGND VPWR VPWR clknet_4_7_0_clock sky130_fd_sc_hd__clkbuf_8
XFILLER_0_133_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12250_ _02187_ _02188_ VGND VGND VPWR VPWR _02189_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11201_ net388 _06623_ VGND VGND VPWR VPWR _01140_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12181_ _01929_ _01998_ VGND VGND VPWR VPWR _02120_ sky130_fd_sc_hd__or2b_1
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11132_ net373 _09583_ VGND VGND VPWR VPWR _01071_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15940_ _06089_ _06091_ VGND VGND VPWR VPWR _06092_ sky130_fd_sc_hd__nand2_1
X_11063_ net367 _01001_ _00887_ VGND VGND VPWR VPWR _01002_ sky130_fd_sc_hd__and3_1
X_10014_ _05666_ _07492_ VGND VGND VPWR VPWR _07503_ sky130_fd_sc_hd__xor2_1
X_15871_ _04304_ _06001_ VGND VGND VPWR VPWR _06016_ sky130_fd_sc_hd__xnor2_1
X_17610_ _07927_ _07928_ VGND VGND VPWR VPWR _07929_ sky130_fd_sc_hd__nor2_1
X_14822_ _04860_ _04861_ net426 kd_2\[5\] VGND VGND VPWR VPWR _04862_ sky130_fd_sc_hd__and4b_1
X_18590_ _06121_ _09000_ _09003_ _09006_ VGND VGND VPWR VPWR _09007_ sky130_fd_sc_hd__o31a_1
X_17541_ _07845_ _07847_ _07852_ VGND VGND VPWR VPWR _07853_ sky130_fd_sc_hd__a21bo_1
X_14753_ _04680_ _04785_ VGND VGND VPWR VPWR _04787_ sky130_fd_sc_hd__or2_1
X_11965_ net205 _01875_ VGND VGND VPWR VPWR _01904_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13704_ _03631_ _03664_ VGND VGND VPWR VPWR _03670_ sky130_fd_sc_hd__xnor2_1
X_10916_ _00830_ _00853_ _00854_ VGND VGND VPWR VPWR _00855_ sky130_fd_sc_hd__a21bo_2
X_17472_ _07775_ _07776_ VGND VGND VPWR VPWR _07777_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_157_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14684_ _04690_ _04706_ _04708_ VGND VGND VPWR VPWR _04711_ sky130_fd_sc_hd__or3_1
X_11896_ _01834_ VGND VGND VPWR VPWR _01835_ sky130_fd_sc_hd__buf_2
XFILLER_0_74_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19211_ clknet_4_15_0_clock _00093_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dfxtp_1
X_16423_ _06473_ _06622_ VGND VGND VPWR VPWR _06624_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13635_ _03536_ _03538_ _03537_ VGND VGND VPWR VPWR _03595_ sky130_fd_sc_hd__o21a_1
X_10847_ _00784_ _00785_ VGND VGND VPWR VPWR _00786_ sky130_fd_sc_hd__nand2_1
X_19142_ net504 i_error\[12\] VGND VGND VPWR VPWR _09564_ sky130_fd_sc_hd__or2_1
X_16354_ _06542_ _06547_ VGND VGND VPWR VPWR _06548_ sky130_fd_sc_hd__nand2_1
X_13566_ _03474_ _03475_ VGND VGND VPWR VPWR _03525_ sky130_fd_sc_hd__nor2_1
X_10778_ _00701_ _00710_ _00716_ VGND VGND VPWR VPWR _00717_ sky130_fd_sc_hd__nand3_1
XFILLER_0_125_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15305_ _05329_ _05328_ VGND VGND VPWR VPWR _05394_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12517_ _02454_ _02447_ _02452_ VGND VGND VPWR VPWR _02456_ sky130_fd_sc_hd__and3_1
X_19073_ _09515_ _09520_ VGND VGND VPWR VPWR _00093_ sky130_fd_sc_hd__nor2_1
X_16285_ net279 _06404_ _06438_ net276 VGND VGND VPWR VPWR _06472_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_14_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13497_ _03403_ _03221_ VGND VGND VPWR VPWR _03456_ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18024_ _08381_ _08384_ VGND VGND VPWR VPWR _08385_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15236_ _05315_ _05317_ VGND VGND VPWR VPWR _05318_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12448_ net209 _01910_ _02318_ VGND VGND VPWR VPWR _02387_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15167_ net441 net181 net178 net447 VGND VGND VPWR VPWR _05242_ sky130_fd_sc_hd__a22oi_2
X_12379_ _02316_ _02317_ VGND VGND VPWR VPWR _02318_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14118_ _04088_ _04089_ VGND VGND VPWR VPWR _04090_ sky130_fd_sc_hd__or2_1
X_15098_ _05057_ _05058_ _05060_ VGND VGND VPWR VPWR _05166_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18926_ _09369_ _09376_ VGND VGND VPWR VPWR _09377_ sky130_fd_sc_hd__xnor2_1
X_14049_ _04018_ _04020_ VGND VGND VPWR VPWR _04021_ sky130_fd_sc_hd__and2_1
XFILLER_0_157_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18857_ _09299_ _09300_ VGND VGND VPWR VPWR _09301_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17808_ _08129_ _08146_ VGND VGND VPWR VPWR _08147_ sky130_fd_sc_hd__and2_1
X_18788_ _06127_ _06129_ _08965_ VGND VGND VPWR VPWR _09225_ sky130_fd_sc_hd__or3_1
XFILLER_0_89_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17739_ _08063_ _08070_ VGND VGND VPWR VPWR _08071_ sky130_fd_sc_hd__or2b_1
XFILLER_0_49_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09926_ _06227_ _06524_ VGND VGND VPWR VPWR _06535_ sky130_fd_sc_hd__or2_1
X_09857_ net353 _05182_ _04896_ net356 VGND VGND VPWR VPWR _05776_ sky130_fd_sc_hd__a22oi_1
X_09788_ _04159_ _04797_ _04786_ _04808_ _04940_ VGND VGND VPWR VPWR _05017_ sky130_fd_sc_hd__a311o_4
XFILLER_0_96_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11750_ _00864_ _00957_ VGND VGND VPWR VPWR _01689_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10701_ net397 _04885_ _00638_ _00639_ VGND VGND VPWR VPWR _00640_ sky130_fd_sc_hd__a31o_1
XFILLER_0_49_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11681_ _01618_ _01619_ VGND VGND VPWR VPWR _01620_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13420_ _03356_ _03360_ _03375_ VGND VGND VPWR VPWR _03377_ sky130_fd_sc_hd__or3_1
X_10632_ _00475_ _00570_ VGND VGND VPWR VPWR _00571_ sky130_fd_sc_hd__xor2_1
XFILLER_0_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13351_ _03287_ _03300_ _03302_ VGND VGND VPWR VPWR _03304_ sky130_fd_sc_hd__and3_1
X_10563_ _00416_ _00501_ VGND VGND VPWR VPWR _00502_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12302_ _02239_ _02234_ VGND VGND VPWR VPWR _02241_ sky130_fd_sc_hd__and2b_1
X_16070_ net349 _08889_ _07448_ VGND VGND VPWR VPWR _06235_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13282_ _03147_ _03146_ VGND VGND VPWR VPWR _03235_ sky130_fd_sc_hd__and2b_1
X_10494_ _00309_ _00310_ VGND VGND VPWR VPWR _00433_ sky130_fd_sc_hd__xor2_1
XFILLER_0_134_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15021_ net409 net194 _05080_ VGND VGND VPWR VPWR _05081_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12233_ _02118_ _02170_ VGND VGND VPWR VPWR _02172_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_15_Left_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12164_ _02050_ _02067_ VGND VGND VPWR VPWR _02103_ sky130_fd_sc_hd__and2_1
X_11115_ net405 net509 _05369_ VGND VGND VPWR VPWR _01054_ sky130_fd_sc_hd__and3_1
X_12095_ _02011_ _02012_ VGND VGND VPWR VPWR _02034_ sky130_fd_sc_hd__nor2_1
X_16972_ _07212_ _07226_ VGND VGND VPWR VPWR _07227_ sky130_fd_sc_hd__nor2_1
X_15923_ _03425_ _03854_ VGND VGND VPWR VPWR _06074_ sky130_fd_sc_hd__xnor2_2
X_18711_ _08918_ _09075_ _09077_ VGND VGND VPWR VPWR _09140_ sky130_fd_sc_hd__nand3b_1
X_11046_ net370 _09583_ _00983_ _00984_ VGND VGND VPWR VPWR _00985_ sky130_fd_sc_hd__a31oi_2
X_18642_ _09063_ _08841_ _08882_ VGND VGND VPWR VPWR _09064_ sky130_fd_sc_hd__mux2_1
X_15854_ _04477_ _05994_ _05997_ VGND VGND VPWR VPWR _05998_ sky130_fd_sc_hd__and3_1
XFILLER_0_36_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14805_ _04733_ _04843_ VGND VGND VPWR VPWR _04844_ sky130_fd_sc_hd__or2_1
X_18573_ _08750_ VGND VGND VPWR VPWR _08989_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_24_Left_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15785_ _05901_ _05902_ VGND VGND VPWR VPWR _05922_ sky130_fd_sc_hd__nand2_1
X_12997_ kd_1\[16\] _02915_ _02747_ net207 VGND VGND VPWR VPWR _02936_ sky130_fd_sc_hd__a22o_1
X_17524_ _07820_ _07834_ VGND VGND VPWR VPWR _07835_ sky130_fd_sc_hd__and2_1
X_14736_ _04573_ _04767_ VGND VGND VPWR VPWR _04768_ sky130_fd_sc_hd__nand2_1
X_11948_ _01882_ _01886_ VGND VGND VPWR VPWR _01887_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17455_ _07732_ _07733_ _07757_ VGND VGND VPWR VPWR _07759_ sky130_fd_sc_hd__a21o_1
X_14667_ net461 net133 VGND VGND VPWR VPWR _04692_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11879_ net213 _01817_ _01810_ net217 VGND VGND VPWR VPWR _01818_ sky130_fd_sc_hd__a22oi_1
X_16406_ _06603_ _06597_ VGND VGND VPWR VPWR _06605_ sky130_fd_sc_hd__and2b_1
X_13618_ net266 _02222_ _03576_ VGND VGND VPWR VPWR _03577_ sky130_fd_sc_hd__and3_1
X_17386_ _07675_ _07593_ _07681_ VGND VGND VPWR VPWR _07683_ sky130_fd_sc_hd__o21ai_1
X_14598_ _04615_ VGND VGND VPWR VPWR _04616_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19125_ _09171_ _09172_ _09550_ VGND VGND VPWR VPWR _09554_ sky130_fd_sc_hd__a21o_1
X_16337_ _06507_ _06528_ VGND VGND VPWR VPWR _06529_ sky130_fd_sc_hd__xor2_1
X_13549_ _03439_ _03507_ VGND VGND VPWR VPWR _03508_ sky130_fd_sc_hd__nor2_1
X_19056_ _09508_ _09509_ net493 VGND VGND VPWR VPWR _00086_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16268_ net289 _06345_ VGND VGND VPWR VPWR _06453_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_33_Left_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18007_ _08332_ _08322_ _08334_ VGND VGND VPWR VPWR _08366_ sky130_fd_sc_hd__a21oi_1
X_15219_ _05289_ _05298_ VGND VGND VPWR VPWR _05299_ sky130_fd_sc_hd__or2_1
X_16199_ ki\[9\] ki\[10\] VGND VGND VPWR VPWR _06377_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09711_ net7 net65 VGND VGND VPWR VPWR _04170_ sky130_fd_sc_hd__or2b_2
X_18909_ net101 _09349_ VGND VGND VPWR VPWR _09358_ sky130_fd_sc_hd__or2b_1
X_09642_ net55 _03358_ _03391_ net245 VGND VGND VPWR VPWR _00015_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09909_ net348 _05754_ _05798_ _05787_ VGND VGND VPWR VPWR _06348_ sky130_fd_sc_hd__a31o_1
X_12920_ _02849_ _02856_ _02858_ VGND VGND VPWR VPWR _02859_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12851_ _02788_ _02783_ _02786_ VGND VGND VPWR VPWR _02790_ sky130_fd_sc_hd__nor3_1
X_11802_ prev_error\[13\] _05292_ _05303_ VGND VGND VPWR VPWR _01741_ sky130_fd_sc_hd__and3_2
X_15570_ _05680_ _05682_ _05684_ VGND VGND VPWR VPWR _05685_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_68_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12782_ net227 _01909_ _02615_ VGND VGND VPWR VPWR _02721_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14521_ _04529_ _04530_ VGND VGND VPWR VPWR _04531_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11733_ _01411_ _01668_ _01407_ VGND VGND VPWR VPWR _01672_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_84_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17240_ net328 _06351_ _07519_ _07520_ VGND VGND VPWR VPWR _07522_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14452_ _04450_ _04452_ _04454_ VGND VGND VPWR VPWR _04455_ sky130_fd_sc_hd__o21ai_1
X_11664_ _01518_ _01588_ _01590_ VGND VGND VPWR VPWR _01603_ sky130_fd_sc_hd__and3_1
XFILLER_0_36_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13403_ _03356_ _03357_ VGND VGND VPWR VPWR _03359_ sky130_fd_sc_hd__nor2_1
X_17171_ _07436_ _07438_ _07445_ VGND VGND VPWR VPWR _07446_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_142_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10615_ _00466_ _00553_ VGND VGND VPWR VPWR _00554_ sky130_fd_sc_hd__xnor2_1
X_14383_ _04377_ _04378_ VGND VGND VPWR VPWR _04380_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11595_ net399 _01001_ _01532_ _01533_ VGND VGND VPWR VPWR _01534_ sky130_fd_sc_hd__a31o_1
X_16122_ prev_error\[9\] _01178_ _01179_ VGND VGND VPWR VPWR _06292_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13334_ _03278_ _03285_ _03286_ VGND VGND VPWR VPWR _03287_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10546_ _00484_ _00385_ VGND VGND VPWR VPWR _00485_ sky130_fd_sc_hd__xor2_1
XFILLER_0_52_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16053_ _06214_ _06215_ VGND VGND VPWR VPWR _06217_ sky130_fd_sc_hd__or2b_1
X_13265_ _03128_ _03217_ VGND VGND VPWR VPWR _03218_ sky130_fd_sc_hd__xor2_1
X_10477_ _00413_ _00415_ VGND VGND VPWR VPWR _00416_ sky130_fd_sc_hd__nand2_1
X_15004_ _05036_ _05062_ VGND VGND VPWR VPWR _05063_ sky130_fd_sc_hd__nor2_1
X_12216_ _01929_ _02154_ VGND VGND VPWR VPWR _02155_ sky130_fd_sc_hd__xnor2_1
X_13196_ _03145_ _03148_ VGND VGND VPWR VPWR _03149_ sky130_fd_sc_hd__and2b_1
X_12147_ _01709_ VGND VGND VPWR VPWR _02086_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16955_ _07205_ _07208_ VGND VGND VPWR VPWR _07209_ sky130_fd_sc_hd__or2b_1
X_12078_ _01978_ _02013_ _02014_ VGND VGND VPWR VPWR _02017_ sky130_fd_sc_hd__or3_1
X_15906_ _03866_ _06054_ VGND VGND VPWR VPWR _06055_ sky130_fd_sc_hd__and2_1
X_11029_ _00962_ _00967_ VGND VGND VPWR VPWR _00968_ sky130_fd_sc_hd__xnor2_4
X_16886_ _07130_ _07132_ VGND VGND VPWR VPWR _07133_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_2_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15837_ _05976_ _05977_ VGND VGND VPWR VPWR _05979_ sky130_fd_sc_hd__nand2_1
X_18625_ _09042_ _09045_ VGND VGND VPWR VPWR _09046_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15768_ _05901_ _05902_ VGND VGND VPWR VPWR _05903_ sky130_fd_sc_hd__nor2_1
X_18556_ _08968_ _08969_ VGND VGND VPWR VPWR _08970_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14719_ _04736_ _04738_ _04748_ VGND VGND VPWR VPWR _04749_ sky130_fd_sc_hd__a21o_1
X_17507_ _07804_ _07806_ VGND VGND VPWR VPWR _07816_ sky130_fd_sc_hd__xor2_1
XFILLER_0_157_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18487_ _08893_ VGND VGND VPWR VPWR _08894_ sky130_fd_sc_hd__inv_2
X_15699_ _05825_ _05826_ VGND VGND VPWR VPWR _05827_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17438_ net282 _07157_ _07648_ _07739_ VGND VGND VPWR VPWR _07740_ sky130_fd_sc_hd__a31o_1
XFILLER_0_157_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_15 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 net431 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_37 net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17369_ _07658_ _07663_ VGND VGND VPWR VPWR _07664_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19108_ net500 prev_error\[15\] VGND VGND VPWR VPWR _09543_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19039_ net563 net94 VGND VGND VPWR VPWR _09496_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09625_ net45 _03091_ _03124_ net136 VGND VGND VPWR VPWR _00024_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10400_ _00328_ _00338_ _00336_ VGND VGND VPWR VPWR _00339_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_22_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11380_ net391 _09558_ _09565_ VGND VGND VPWR VPWR _01319_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10331_ _00255_ _00256_ VGND VGND VPWR VPWR _00270_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10262_ _00193_ _00196_ _00200_ VGND VGND VPWR VPWR _00201_ sky130_fd_sc_hd__a21o_1
X_13050_ net269 _01859_ VGND VGND VPWR VPWR _02989_ sky130_fd_sc_hd__nand2_2
X_12001_ net218 _01787_ _01810_ net215 VGND VGND VPWR VPWR _01940_ sky130_fd_sc_hd__a22oi_1
X_10193_ _09450_ _09461_ VGND VGND VPWR VPWR _09472_ sky130_fd_sc_hd__nand2_2
XFILLER_0_100_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout360 net361 VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout371 net373 VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__clkbuf_4
X_16740_ _06957_ _06971_ VGND VGND VPWR VPWR _06972_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout382 kp\[5\] VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__buf_2
X_13952_ net440 net119 net116 net444 VGND VGND VPWR VPWR _03924_ sky130_fd_sc_hd__a22o_1
Xfanout393 kp\[3\] VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_89_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12903_ net224 _02223_ VGND VGND VPWR VPWR _02842_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16671_ _06888_ _06894_ _06895_ VGND VGND VPWR VPWR _06896_ sky130_fd_sc_hd__o21ai_2
X_13883_ _03551_ _03552_ VGND VGND VPWR VPWR _03849_ sky130_fd_sc_hd__nor2_1
X_15622_ _05682_ _05741_ VGND VGND VPWR VPWR _05742_ sky130_fd_sc_hd__nor2_1
X_18410_ _08567_ _08552_ VGND VGND VPWR VPWR _08809_ sky130_fd_sc_hd__or2b_1
X_12834_ _02766_ _02764_ VGND VGND VPWR VPWR _02773_ sky130_fd_sc_hd__xor2_1
X_18341_ _08620_ _08732_ VGND VGND VPWR VPWR _08733_ sky130_fd_sc_hd__nand2_1
X_15553_ _05660_ _05664_ _05603_ _05635_ VGND VGND VPWR VPWR _05667_ sky130_fd_sc_hd__o211ai_2
X_12765_ _02598_ _02703_ VGND VGND VPWR VPWR _02704_ sky130_fd_sc_hd__xor2_2
XFILLER_0_57_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14504_ _04509_ _04512_ VGND VGND VPWR VPWR _04513_ sky130_fd_sc_hd__and2_1
X_11716_ _01644_ _01643_ VGND VGND VPWR VPWR _01655_ sky130_fd_sc_hd__xnor2_1
X_18272_ net290 net287 VGND VGND VPWR VPWR _08657_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15484_ _05587_ _05577_ _05590_ VGND VGND VPWR VPWR _05591_ sky130_fd_sc_hd__o21a_1
X_12696_ net207 _02545_ VGND VGND VPWR VPWR _02635_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17223_ net302 _06891_ _07502_ _07500_ VGND VGND VPWR VPWR _07504_ sky130_fd_sc_hd__a31o_1
X_14435_ _04409_ _04433_ _04436_ VGND VGND VPWR VPWR _04437_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11647_ _01573_ _01575_ _01574_ VGND VGND VPWR VPWR _01586_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput13 measurement[2] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_1
X_17154_ _07409_ _07419_ _07427_ VGND VGND VPWR VPWR _07428_ sky130_fd_sc_hd__a21bo_1
Xinput24 reg_addr[12] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14366_ _04017_ net165 VGND VGND VPWR VPWR _04361_ sky130_fd_sc_hd__nor2_1
Xinput35 reg_addr[5] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput46 reg_data[15] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_4
X_11578_ _01513_ _01515_ VGND VGND VPWR VPWR _01517_ sky130_fd_sc_hd__xnor2_1
Xinput57 reg_data[8] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__buf_4
XFILLER_0_107_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput68 target[17] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16105_ prev_error\[4\] _00408_ VGND VGND VPWR VPWR _06274_ sky130_fd_sc_hd__or2_1
X_13317_ _03267_ _03269_ VGND VGND VPWR VPWR _03270_ sky130_fd_sc_hd__or2_1
X_10529_ net387 _00363_ _04885_ VGND VGND VPWR VPWR _00468_ sky130_fd_sc_hd__and3_1
X_17085_ _07346_ _07351_ VGND VGND VPWR VPWR _07352_ sky130_fd_sc_hd__nand2_1
Xinput79 write_enable VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_4
X_14297_ _04256_ _04284_ VGND VGND VPWR VPWR _04285_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16036_ _06196_ _06197_ VGND VGND VPWR VPWR _06198_ sky130_fd_sc_hd__nor2_1
X_13248_ _03198_ _03200_ VGND VGND VPWR VPWR _03201_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13179_ net220 _02640_ _02746_ net216 VGND VGND VPWR VPWR _03131_ sky130_fd_sc_hd__a22o_1
X_17987_ _08283_ _08291_ _08290_ VGND VGND VPWR VPWR _08344_ sky130_fd_sc_hd__o21a_1
X_16938_ _07178_ _07179_ _07189_ VGND VGND VPWR VPWR _07190_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_79_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16869_ _07084_ _07113_ VGND VGND VPWR VPWR _07114_ sky130_fd_sc_hd__and2_1
X_18608_ _08858_ _08861_ _08882_ VGND VGND VPWR VPWR _09027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18539_ _08898_ net528 _08755_ _08764_ _08899_ VGND VGND VPWR VPWR _08951_ sky130_fd_sc_hd__a32oi_1
XFILLER_0_90_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09608_ _03069_ _03080_ net487 VGND VGND VPWR VPWR _03113_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10880_ net343 _00818_ VGND VGND VPWR VPWR _00819_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12550_ _02483_ _02487_ VGND VGND VPWR VPWR _02489_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11501_ _01437_ _01415_ _01438_ _01439_ VGND VGND VPWR VPWR _01440_ sky130_fd_sc_hd__nand4_1
X_12481_ _02398_ _02417_ VGND VGND VPWR VPWR _02420_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14220_ _04127_ _04199_ VGND VGND VPWR VPWR _04200_ sky130_fd_sc_hd__nor2_1
X_11432_ _01329_ _01370_ VGND VGND VPWR VPWR _01371_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14151_ _04059_ _04062_ _04122_ _04123_ VGND VGND VPWR VPWR _04124_ sky130_fd_sc_hd__o211a_1
X_11363_ _01235_ _01301_ VGND VGND VPWR VPWR _01302_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13102_ _02965_ _03022_ _03005_ _03021_ VGND VGND VPWR VPWR _03046_ sky130_fd_sc_hd__a211o_1
X_10314_ _00237_ _00251_ _00228_ VGND VGND VPWR VPWR _00253_ sky130_fd_sc_hd__o21a_1
X_14082_ _04051_ _04053_ VGND VGND VPWR VPWR _04054_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11294_ net366 _00515_ _00613_ net362 VGND VGND VPWR VPWR _01233_ sky130_fd_sc_hd__a22oi_1
X_13033_ _02833_ _02946_ _02967_ _02971_ VGND VGND VPWR VPWR _02972_ sky130_fd_sc_hd__o211ai_2
X_17910_ _08245_ _08247_ _08258_ VGND VGND VPWR VPWR _08259_ sky130_fd_sc_hd__a21bo_1
X_10245_ _00182_ _00183_ VGND VGND VPWR VPWR _00184_ sky130_fd_sc_hd__nand2_1
X_18890_ _09335_ _09336_ VGND VGND VPWR VPWR _09337_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10176_ net360 _05424_ _07888_ VGND VGND VPWR VPWR _09285_ sky130_fd_sc_hd__a21oi_1
X_17841_ _08181_ _08176_ VGND VGND VPWR VPWR _08183_ sky130_fd_sc_hd__and2b_1
X_14984_ _05037_ _05040_ VGND VGND VPWR VPWR _05041_ sky130_fd_sc_hd__nor2_1
X_17772_ net334 _06890_ VGND VGND VPWR VPWR _08107_ sky130_fd_sc_hd__nand2_1
Xfanout190 kd_2\[2\] VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16723_ _06951_ _06952_ VGND VGND VPWR VPWR _06954_ sky130_fd_sc_hd__nand2_1
X_13935_ _03898_ _03900_ _03897_ VGND VGND VPWR VPWR _03906_ sky130_fd_sc_hd__o21ba_1
X_16654_ _06875_ _06877_ VGND VGND VPWR VPWR _06878_ sky130_fd_sc_hd__and2_1
X_13866_ _02747_ _03792_ _03811_ _03220_ net267 VGND VGND VPWR VPWR _03832_ sky130_fd_sc_hd__o2111a_1
X_15605_ _05659_ _05663_ _05662_ VGND VGND VPWR VPWR _05724_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_147_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12817_ _02736_ _02755_ VGND VGND VPWR VPWR _02756_ sky130_fd_sc_hd__and2b_1
XFILLER_0_85_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16585_ _06801_ VGND VGND VPWR VPWR _06802_ sky130_fd_sc_hd__clkbuf_4
X_13797_ _03761_ _03762_ VGND VGND VPWR VPWR _03763_ sky130_fd_sc_hd__xor2_1
X_15536_ _05645_ _05647_ VGND VGND VPWR VPWR _05648_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18324_ _08675_ _08714_ VGND VGND VPWR VPWR _08715_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12748_ net255 net199 _01813_ _02686_ VGND VGND VPWR VPWR _02687_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18255_ _08632_ _08638_ VGND VGND VPWR VPWR _08639_ sky130_fd_sc_hd__and2_1
X_15467_ _05569_ _05570_ _05571_ VGND VGND VPWR VPWR _05572_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_72_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12679_ net222 _01909_ _02616_ _02617_ VGND VGND VPWR VPWR _02618_ sky130_fd_sc_hd__and4_1
XFILLER_0_44_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17206_ net328 net514 VGND VGND VPWR VPWR _07485_ sky130_fd_sc_hd__nand2_1
X_14418_ _04416_ _04414_ VGND VGND VPWR VPWR _04418_ sky130_fd_sc_hd__xnor2_1
X_18186_ i_error\[1\] _08434_ _08561_ VGND VGND VPWR VPWR _08563_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_7_Left_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15398_ net452 net181 net177 net457 VGND VGND VPWR VPWR _05496_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_53_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17137_ _07368_ _07378_ _07408_ VGND VGND VPWR VPWR _07409_ sky130_fd_sc_hd__a21bo_1
X_14349_ _04251_ _04253_ VGND VGND VPWR VPWR _04342_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17068_ _07328_ _07331_ _07330_ VGND VGND VPWR VPWR _07333_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_100_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16019_ net339 _05754_ _08603_ _08592_ VGND VGND VPWR VPWR _06179_ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09890_ net344 net341 _05996_ _06073_ VGND VGND VPWR VPWR _06139_ sky130_fd_sc_hd__and4_1
XFILLER_0_85_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10030_ _07657_ _07668_ VGND VGND VPWR VPWR _07679_ sky130_fd_sc_hd__nor2_1
Xclkbuf_4_3_0_clock clknet_0_clock VGND VGND VPWR VPWR clknet_4_3_0_clock sky130_fd_sc_hd__clkbuf_8
X_11981_ _01903_ _01918_ _01896_ VGND VGND VPWR VPWR _01920_ sky130_fd_sc_hd__a21oi_1
X_13720_ _03679_ _03685_ VGND VGND VPWR VPWR _03686_ sky130_fd_sc_hd__nor2_1
X_10932_ net405 VGND VGND VPWR VPWR _00871_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13651_ net251 _02544_ VGND VGND VPWR VPWR _03612_ sky130_fd_sc_hd__nand2_1
X_10863_ net346 _00516_ _00801_ VGND VGND VPWR VPWR _00802_ sky130_fd_sc_hd__and3_1
XFILLER_0_155_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12602_ _01722_ _01712_ VGND VGND VPWR VPWR _02541_ sky130_fd_sc_hd__nor2b_4
XFILLER_0_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16370_ _06563_ _06564_ VGND VGND VPWR VPWR _06565_ sky130_fd_sc_hd__xor2_1
X_13582_ _03536_ net107 _03484_ _03540_ VGND VGND VPWR VPWR _03541_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_93_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10794_ net397 _05138_ _05149_ VGND VGND VPWR VPWR _00733_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15321_ _05392_ _05389_ VGND VGND VPWR VPWR _05411_ sky130_fd_sc_hd__nor2_1
X_12533_ _02449_ _02451_ VGND VGND VPWR VPWR _02472_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18040_ _08388_ _08390_ _08393_ _08401_ VGND VGND VPWR VPWR _08402_ sky130_fd_sc_hd__or4b_1
X_15252_ _05239_ _05302_ VGND VGND VPWR VPWR _05335_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12464_ _02334_ _02402_ VGND VGND VPWR VPWR _02403_ sky130_fd_sc_hd__and2_1
X_14203_ _04017_ net140 _04180_ VGND VGND VPWR VPWR _04182_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11415_ _01352_ _01353_ VGND VGND VPWR VPWR _01354_ sky130_fd_sc_hd__nor2_1
X_15183_ _05256_ _05257_ _05247_ _05252_ VGND VGND VPWR VPWR _05260_ sky130_fd_sc_hd__a211o_1
XFILLER_0_105_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12395_ net201 _02332_ _02333_ VGND VGND VPWR VPWR _02334_ sky130_fd_sc_hd__nand3_1
X_14134_ _04071_ _04072_ _04073_ VGND VGND VPWR VPWR _04106_ sky130_fd_sc_hd__o21ba_1
X_11346_ net564 _05963_ _05974_ net385 _09577_ VGND VGND VPWR VPWR _01285_ sky130_fd_sc_hd__a32o_1
X_18942_ net201 _01810_ VGND VGND VPWR VPWR _09394_ sky130_fd_sc_hd__nand2_1
X_14065_ _04035_ _04036_ VGND VGND VPWR VPWR _04037_ sky130_fd_sc_hd__nor2_1
X_11277_ net406 net386 _08185_ _06051_ VGND VGND VPWR VPWR _01216_ sky130_fd_sc_hd__and4_1
X_13016_ _02950_ _02952_ _02954_ VGND VGND VPWR VPWR _02955_ sky130_fd_sc_hd__o21ai_1
X_10228_ _00162_ _00164_ VGND VGND VPWR VPWR _00167_ sky130_fd_sc_hd__nand2_1
X_18873_ _09316_ _09317_ VGND VGND VPWR VPWR _09319_ sky130_fd_sc_hd__and2_1
X_17824_ _08159_ _08161_ VGND VGND VPWR VPWR _08165_ sky130_fd_sc_hd__nand2_2
X_10159_ _09076_ _09087_ VGND VGND VPWR VPWR _09098_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14967_ net472 net144 net138 net474 VGND VGND VPWR VPWR _05022_ sky130_fd_sc_hd__a22oi_2
X_17755_ net301 net540 _08084_ _08088_ VGND VGND VPWR VPWR _08089_ sky130_fd_sc_hd__a31o_1
X_16706_ _06838_ _06932_ VGND VGND VPWR VPWR _06935_ sky130_fd_sc_hd__xor2_1
X_13918_ _02464_ _03884_ _03886_ VGND VGND VPWR VPWR _03887_ sky130_fd_sc_hd__o21ai_1
X_14898_ _04873_ _04945_ VGND VGND VPWR VPWR _04946_ sky130_fd_sc_hd__nand2_1
X_17686_ _07995_ _08011_ _08012_ _07919_ VGND VGND VPWR VPWR _08013_ sky130_fd_sc_hd__o211a_1
X_16637_ _06687_ _06774_ _06773_ VGND VGND VPWR VPWR _06859_ sky130_fd_sc_hd__o21a_1
X_13849_ _03680_ _03814_ VGND VGND VPWR VPWR _03815_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16568_ _06770_ _06782_ VGND VGND VPWR VPWR _06783_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18307_ _08634_ _08659_ VGND VGND VPWR VPWR _08696_ sky130_fd_sc_hd__xor2_1
XFILLER_0_127_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15519_ _05623_ _05628_ VGND VGND VPWR VPWR _05629_ sky130_fd_sc_hd__and2_1
XFILLER_0_143_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19287_ clknet_4_7_0_clock _00065_ VGND VGND VPWR VPWR kp\[17\] sky130_fd_sc_hd__dfxtp_1
X_16499_ _06682_ _06704_ _06706_ VGND VGND VPWR VPWR _06707_ sky130_fd_sc_hd__a21o_1
X_18238_ _08619_ VGND VGND VPWR VPWR _08620_ sky130_fd_sc_hd__buf_4
XFILLER_0_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18169_ i_error\[5\] _08543_ VGND VGND VPWR VPWR _08544_ sky130_fd_sc_hd__nor2_1
Xmax_cap110 _08299_ VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__buf_1
XFILLER_0_13_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09942_ _06568_ _06689_ _06700_ VGND VGND VPWR VPWR _06711_ sky130_fd_sc_hd__o21a_1
XFILLER_0_110_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09873_ _05347_ _05446_ VGND VGND VPWR VPWR _05952_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11200_ _01063_ _01138_ VGND VGND VPWR VPWR _01139_ sky130_fd_sc_hd__xnor2_1
X_12180_ _01952_ _01966_ _01969_ VGND VGND VPWR VPWR _02119_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_102_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11131_ _00984_ _00983_ VGND VGND VPWR VPWR _01070_ sky130_fd_sc_hd__and2b_1
XFILLER_0_102_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_79_Left_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11062_ _00323_ VGND VGND VPWR VPWR _01001_ sky130_fd_sc_hd__buf_4
X_10013_ _06920_ _07481_ VGND VGND VPWR VPWR _07492_ sky130_fd_sc_hd__xor2_1
X_15870_ _03886_ _06014_ VGND VGND VPWR VPWR _06015_ sky130_fd_sc_hd__xnor2_1
X_14821_ net567 net174 net169 net436 VGND VGND VPWR VPWR _04861_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14752_ _04780_ _04784_ VGND VGND VPWR VPWR _04785_ sky130_fd_sc_hd__and2_1
X_17540_ _07848_ _07849_ _07851_ VGND VGND VPWR VPWR _07852_ sky130_fd_sc_hd__or3_1
X_11964_ _01897_ _01900_ _01902_ VGND VGND VPWR VPWR _01903_ sky130_fd_sc_hd__o21ai_1
X_13703_ _03550_ _03668_ VGND VGND VPWR VPWR _03669_ sky130_fd_sc_hd__xnor2_1
X_17471_ _07205_ _07208_ VGND VGND VPWR VPWR _07776_ sky130_fd_sc_hd__xnor2_2
X_10915_ _00848_ _00852_ _00831_ _00832_ VGND VGND VPWR VPWR _00854_ sky130_fd_sc_hd__a211o_1
X_14683_ _04690_ _04706_ _04708_ VGND VGND VPWR VPWR _04710_ sky130_fd_sc_hd__o21ai_1
X_11895_ _01739_ _01742_ VGND VGND VPWR VPWR _01834_ sky130_fd_sc_hd__xnor2_4
XPHY_EDGE_ROW_88_Left_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19210_ clknet_4_15_0_clock _00092_ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dfxtp_1
X_16422_ net275 _06470_ VGND VGND VPWR VPWR _06622_ sky130_fd_sc_hd__nand2_1
X_13634_ _03589_ _03591_ _03593_ VGND VGND VPWR VPWR _03594_ sky130_fd_sc_hd__nand3_2
X_10846_ _00783_ _00778_ VGND VGND VPWR VPWR _00785_ sky130_fd_sc_hd__or2b_1
XFILLER_0_55_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19141_ _09559_ _09028_ _09563_ net496 VGND VGND VPWR VPWR _00125_ sky130_fd_sc_hd__o211a_1
X_16353_ _06543_ _06544_ _06545_ VGND VGND VPWR VPWR _06547_ sky130_fd_sc_hd__mux2_2
X_13565_ _03486_ _03489_ _03488_ VGND VGND VPWR VPWR _03524_ sky130_fd_sc_hd__o21a_1
X_10777_ _00713_ _00715_ VGND VGND VPWR VPWR _00716_ sky130_fd_sc_hd__nand2_2
X_15304_ _05389_ _05390_ _05392_ VGND VGND VPWR VPWR _05393_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_82_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12516_ _02447_ _02452_ _02454_ VGND VGND VPWR VPWR _02455_ sky130_fd_sc_hd__a21oi_1
X_19072_ net506 net546 net496 VGND VGND VPWR VPWR _09520_ sky130_fd_sc_hd__o21ai_1
X_16284_ net272 _06470_ VGND VGND VPWR VPWR _06471_ sky130_fd_sc_hd__nand2_1
X_13496_ _03445_ _03454_ VGND VGND VPWR VPWR _03455_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15235_ _05309_ _05316_ VGND VGND VPWR VPWR _05317_ sky130_fd_sc_hd__and2_1
X_18023_ _08370_ _08382_ VGND VGND VPWR VPWR _08384_ sky130_fd_sc_hd__or2_1
X_12447_ _02379_ _02385_ VGND VGND VPWR VPWR _02386_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15166_ net437 net184 VGND VGND VPWR VPWR _05241_ sky130_fd_sc_hd__nand2_1
X_12378_ net219 _01853_ _01874_ net214 VGND VGND VPWR VPWR _02317_ sky130_fd_sc_hd__a22oi_1
XPHY_EDGE_ROW_97_Left_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14117_ _03921_ _04087_ VGND VGND VPWR VPWR _04089_ sky130_fd_sc_hd__nor2_1
X_11329_ _01265_ _01266_ _01267_ VGND VGND VPWR VPWR _01268_ sky130_fd_sc_hd__nand3_4
X_15097_ _05140_ _05162_ _05163_ _05164_ VGND VGND VPWR VPWR _05165_ sky130_fd_sc_hd__nor4_1
X_14048_ _04015_ _04019_ VGND VGND VPWR VPWR _04020_ sky130_fd_sc_hd__nor2_1
X_18925_ _09370_ _09375_ VGND VGND VPWR VPWR _09376_ sky130_fd_sc_hd__xnor2_1
X_18856_ _02134_ _09286_ _09298_ VGND VGND VPWR VPWR _09300_ sky130_fd_sc_hd__and3_1
X_17807_ _08134_ _08144_ VGND VGND VPWR VPWR _08146_ sky130_fd_sc_hd__xnor2_1
X_18787_ _08982_ _08996_ _09206_ _08981_ VGND VGND VPWR VPWR _09224_ sky130_fd_sc_hd__a31o_1
X_15999_ _06155_ _06156_ VGND VGND VPWR VPWR _06157_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_82_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17738_ _08063_ _08065_ _08068_ _08069_ VGND VGND VPWR VPWR _08070_ sky130_fd_sc_hd__or4bb_1
X_17669_ _07993_ _07901_ VGND VGND VPWR VPWR _07994_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_92_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19339_ clknet_4_2_0_clock _00022_ VGND VGND VPWR VPWR kd_2\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09925_ net338 _06194_ _06216_ VGND VGND VPWR VPWR _06524_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_111_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09856_ net348 _05754_ VGND VGND VPWR VPWR _05765_ sky130_fd_sc_hd__nand2_1
X_09787_ net539 VGND VGND VPWR VPWR _05006_ sky130_fd_sc_hd__buf_2
XFILLER_0_96_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10700_ net393 net568 _05171_ VGND VGND VPWR VPWR _00639_ sky130_fd_sc_hd__and3_1
X_11680_ net390 _00810_ _00814_ net394 VGND VGND VPWR VPWR _01619_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_36_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10631_ _00478_ _00476_ VGND VGND VPWR VPWR _00570_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13350_ _03287_ _03300_ _03302_ VGND VGND VPWR VPWR _03303_ sky130_fd_sc_hd__a21oi_1
X_10562_ _00413_ _00415_ VGND VGND VPWR VPWR _00501_ sky130_fd_sc_hd__or2_1
X_12301_ _02234_ _02239_ VGND VGND VPWR VPWR _02240_ sky130_fd_sc_hd__and2b_1
XFILLER_0_51_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13281_ net265 _01834_ VGND VGND VPWR VPWR _03234_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10493_ _00379_ _00392_ VGND VGND VPWR VPWR _00432_ sky130_fd_sc_hd__xor2_1
XFILLER_0_51_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15020_ _05078_ _05079_ VGND VGND VPWR VPWR _05080_ sky130_fd_sc_hd__nor2_1
X_12232_ _02118_ _02170_ VGND VGND VPWR VPWR _02171_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12163_ _02075_ _02098_ _02101_ VGND VGND VPWR VPWR _02102_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11114_ net388 _06172_ VGND VGND VPWR VPWR _01053_ sky130_fd_sc_hd__nand2_1
X_12094_ _02032_ VGND VGND VPWR VPWR _02033_ sky130_fd_sc_hd__inv_2
X_16971_ net311 _06401_ VGND VGND VPWR VPWR _07226_ sky130_fd_sc_hd__nand2_2
X_18710_ _08961_ _08962_ _08781_ _08881_ _09138_ VGND VGND VPWR VPWR _09139_ sky130_fd_sc_hd__a221o_1
X_15922_ _05950_ _06071_ VGND VGND VPWR VPWR _06072_ sky130_fd_sc_hd__and2_1
X_11045_ net378 _06612_ _00982_ VGND VGND VPWR VPWR _00984_ sky130_fd_sc_hd__and3_1
XFILLER_0_36_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18641_ _08843_ VGND VGND VPWR VPWR _09063_ sky130_fd_sc_hd__inv_2
X_15853_ _05987_ _05995_ VGND VGND VPWR VPWR _05997_ sky130_fd_sc_hd__or2_1
X_14804_ _04729_ _04732_ VGND VGND VPWR VPWR _04843_ sky130_fd_sc_hd__nor2_1
X_18572_ _06122_ _08986_ VGND VGND VPWR VPWR _08987_ sky130_fd_sc_hd__xnor2_4
X_15784_ _05907_ _05909_ _05920_ VGND VGND VPWR VPWR _05921_ sky130_fd_sc_hd__and3_1
X_12996_ _02934_ VGND VGND VPWR VPWR _02935_ sky130_fd_sc_hd__buf_4
XFILLER_0_86_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17523_ _07807_ _07817_ _07819_ VGND VGND VPWR VPWR _07834_ sky130_fd_sc_hd__nand3_1
XFILLER_0_157_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11947_ _01884_ _01885_ VGND VGND VPWR VPWR _01886_ sky130_fd_sc_hd__and2_1
X_14735_ _04570_ _04572_ VGND VGND VPWR VPWR _04767_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14666_ _04689_ _04690_ VGND VGND VPWR VPWR _04691_ sky130_fd_sc_hd__nor2_1
X_17454_ _07732_ _07733_ _07757_ VGND VGND VPWR VPWR _07758_ sky130_fd_sc_hd__nand3_2
X_11878_ _01814_ VGND VGND VPWR VPWR _01817_ sky130_fd_sc_hd__clkbuf_4
X_13617_ _03574_ _03575_ VGND VGND VPWR VPWR _03576_ sky130_fd_sc_hd__nor2_1
X_16405_ _06597_ _06603_ VGND VGND VPWR VPWR _06604_ sky130_fd_sc_hd__and2b_1
XFILLER_0_156_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10829_ _00763_ _00767_ VGND VGND VPWR VPWR _00768_ sky130_fd_sc_hd__and2b_1
X_14597_ net470 net124 net121 net475 VGND VGND VPWR VPWR _04615_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17385_ _07675_ _07593_ _07681_ VGND VGND VPWR VPWR _07682_ sky130_fd_sc_hd__or3_1
X_19124_ _09536_ _09091_ _09553_ net494 VGND VGND VPWR VPWR _00117_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13548_ net236 _02641_ _03438_ VGND VGND VPWR VPWR _03507_ sky130_fd_sc_hd__a21oi_1
X_16336_ _06526_ _06527_ VGND VGND VPWR VPWR _06528_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19055_ _09447_ _09484_ _09452_ VGND VGND VPWR VPWR _09509_ sky130_fd_sc_hd__a21oi_1
X_16267_ _06437_ VGND VGND VPWR VPWR _06452_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13479_ _03371_ _03437_ VGND VGND VPWR VPWR _03438_ sky130_fd_sc_hd__xor2_1
XFILLER_0_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15218_ _05268_ _05280_ _05288_ VGND VGND VPWR VPWR _05298_ sky130_fd_sc_hd__nor3_1
X_18006_ _08358_ _08364_ VGND VGND VPWR VPWR _08365_ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16198_ _06372_ _06375_ VGND VGND VPWR VPWR _06376_ sky130_fd_sc_hd__nor2_4
XFILLER_0_22_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15149_ _05219_ _05221_ VGND VGND VPWR VPWR _05222_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09710_ net8 net66 VGND VGND VPWR VPWR _04159_ sky130_fd_sc_hd__or2b_2
X_18908_ _09353_ _09224_ _09352_ VGND VGND VPWR VPWR _09357_ sky130_fd_sc_hd__a21o_1
X_09641_ net54 _03358_ _03391_ net249 VGND VGND VPWR VPWR _00014_ sky130_fd_sc_hd__a22o_1
X_18839_ _02122_ _02140_ _02138_ VGND VGND VPWR VPWR _09281_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09908_ _06293_ _06326_ VGND VGND VPWR VPWR _06337_ sky130_fd_sc_hd__xnor2_1
X_09839_ _05556_ _05567_ _05072_ VGND VGND VPWR VPWR _05578_ sky130_fd_sc_hd__and3b_1
X_12850_ _02783_ _02786_ _02788_ VGND VGND VPWR VPWR _02789_ sky130_fd_sc_hd__o21a_1
X_11801_ prev_error\[13\] _05314_ VGND VGND VPWR VPWR _01740_ sky130_fd_sc_hd__nor2_2
X_12781_ _02618_ _02719_ VGND VGND VPWR VPWR _02720_ sky130_fd_sc_hd__or2b_1
X_14520_ net421 net165 _04527_ _04528_ VGND VGND VPWR VPWR _04530_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_68_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11732_ _01411_ _01666_ _01670_ VGND VGND VPWR VPWR _01671_ sky130_fd_sc_hd__and3b_2
XFILLER_0_56_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14451_ _04449_ _04453_ VGND VGND VPWR VPWR _04454_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11663_ _01595_ _01600_ _01601_ VGND VGND VPWR VPWR _01602_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_153_Right_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13402_ _02989_ _03355_ VGND VGND VPWR VPWR _03357_ sky130_fd_sc_hd__and2_1
X_17170_ _07435_ _07439_ VGND VGND VPWR VPWR _07445_ sky130_fd_sc_hd__or2b_1
X_10614_ _00527_ _00552_ _00550_ VGND VGND VPWR VPWR _00553_ sky130_fd_sc_hd__a21oi_1
X_14382_ _04367_ _04370_ VGND VGND VPWR VPWR _04378_ sky130_fd_sc_hd__nand2_1
X_11594_ net390 _00514_ _01488_ VGND VGND VPWR VPWR _01533_ sky130_fd_sc_hd__and3_1
XFILLER_0_52_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16121_ prev_error\[8\] _08185_ VGND VGND VPWR VPWR _06291_ sky130_fd_sc_hd__and2_1
X_13333_ _03203_ _03212_ VGND VGND VPWR VPWR _03286_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10545_ net361 _06183_ VGND VGND VPWR VPWR _00484_ sky130_fd_sc_hd__nand2_1
X_16052_ _08537_ _08757_ _08801_ VGND VGND VPWR VPWR _06215_ sky130_fd_sc_hd__a21bo_1
X_13264_ _03066_ _03137_ VGND VGND VPWR VPWR _03217_ sky130_fd_sc_hd__nand2_1
X_10476_ _00405_ _00414_ VGND VGND VPWR VPWR _00415_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15003_ _05057_ _05058_ _05060_ VGND VGND VPWR VPWR _05062_ sky130_fd_sc_hd__and3_1
X_12215_ _02152_ _02153_ VGND VGND VPWR VPWR _02154_ sky130_fd_sc_hd__xor2_1
XFILLER_0_110_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13195_ net265 _01834_ _03146_ _03147_ VGND VGND VPWR VPWR _03148_ sky130_fd_sc_hd__a31o_1
XFILLER_0_103_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12146_ _01710_ _01728_ _01729_ _01730_ VGND VGND VPWR VPWR _02085_ sky130_fd_sc_hd__a31o_2
X_16954_ _07177_ _07207_ VGND VGND VPWR VPWR _07208_ sky130_fd_sc_hd__and2_1
X_12077_ _01845_ _01832_ _01843_ VGND VGND VPWR VPWR _02016_ sky130_fd_sc_hd__nor3_1
X_15905_ _03865_ _03178_ _03863_ VGND VGND VPWR VPWR _06054_ sky130_fd_sc_hd__nand3_1
X_11028_ _00963_ _00966_ VGND VGND VPWR VPWR _00967_ sky130_fd_sc_hd__and2b_2
X_16885_ _07131_ _07022_ VGND VGND VPWR VPWR _07132_ sky130_fd_sc_hd__xor2_2
X_18624_ _06165_ _09041_ VGND VGND VPWR VPWR _09045_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15836_ _05976_ _05977_ VGND VGND VPWR VPWR _05978_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18555_ _08967_ _01698_ VGND VGND VPWR VPWR _08969_ sky130_fd_sc_hd__or2b_1
X_15767_ _05896_ _05900_ VGND VGND VPWR VPWR _05902_ sky130_fd_sc_hd__xnor2_1
X_12979_ _02856_ _02917_ VGND VGND VPWR VPWR _02918_ sky130_fd_sc_hd__nand2_1
X_17506_ _07809_ _07814_ VGND VGND VPWR VPWR _07815_ sky130_fd_sc_hd__nand2_1
X_14718_ _04557_ _04579_ VGND VGND VPWR VPWR _04748_ sky130_fd_sc_hd__xnor2_1
X_18486_ _06174_ _06265_ _08892_ VGND VGND VPWR VPWR _08893_ sky130_fd_sc_hd__or3_2
X_15698_ _05736_ _05783_ VGND VGND VPWR VPWR _05826_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17437_ _07254_ _07590_ VGND VGND VPWR VPWR _07739_ sky130_fd_sc_hd__nor2_1
X_14649_ _04670_ _04671_ VGND VGND VPWR VPWR _04672_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_16 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_120_Right_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_27 net440 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17368_ _07563_ _07659_ _07662_ VGND VGND VPWR VPWR _07663_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_12_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19107_ _09536_ _05754_ _09542_ net488 VGND VGND VPWR VPWR _00109_ sky130_fd_sc_hd__o211a_1
X_16319_ _06416_ _06424_ VGND VGND VPWR VPWR _06509_ sky130_fd_sc_hd__and2_1
XFILLER_0_141_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17299_ _07550_ _07551_ _07553_ VGND VGND VPWR VPWR _07587_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_113_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19038_ _09494_ _09495_ net492 VGND VGND VPWR VPWR _00080_ sky130_fd_sc_hd__o21a_1
XFILLER_0_112_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09624_ net44 _03091_ _03124_ net137 VGND VGND VPWR VPWR _00023_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10330_ _00261_ _00259_ VGND VGND VPWR VPWR _00269_ sky130_fd_sc_hd__xor2_4
XFILLER_0_104_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10261_ _00195_ _05545_ VGND VGND VPWR VPWR _00200_ sky130_fd_sc_hd__and2b_1
XFILLER_0_103_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12000_ net210 _01817_ VGND VGND VPWR VPWR _01939_ sky130_fd_sc_hd__nand2_1
X_10192_ _09252_ _09417_ _09439_ VGND VGND VPWR VPWR _09461_ sky130_fd_sc_hd__nand3_1
Xfanout350 kp\[14\] VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout361 kp\[11\] VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__buf_2
Xfanout372 net373 VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__buf_2
X_13951_ net440 net444 net117 VGND VGND VPWR VPWR _03923_ sky130_fd_sc_hd__and3_1
Xfanout383 net384 VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__clkbuf_4
Xfanout394 net398 VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__clkbuf_4
X_12902_ _01847_ _02747_ VGND VGND VPWR VPWR _02841_ sky130_fd_sc_hd__or2_1
X_16670_ _06883_ _06886_ VGND VGND VPWR VPWR _06895_ sky130_fd_sc_hd__xor2_1
X_13882_ _03554_ _03667_ _03669_ _03847_ VGND VGND VPWR VPWR _03848_ sky130_fd_sc_hd__or4bb_1
X_12833_ _02769_ _02771_ VGND VGND VPWR VPWR _02772_ sky130_fd_sc_hd__nor2_1
X_15621_ net478 net171 _05680_ _05681_ VGND VGND VPWR VPWR _05741_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_96_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18340_ _06261_ _08731_ VGND VGND VPWR VPWR _08732_ sky130_fd_sc_hd__nand2_1
X_12764_ net238 _01860_ VGND VGND VPWR VPWR _02703_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15552_ _05603_ _05635_ _05660_ _05664_ VGND VGND VPWR VPWR _05665_ sky130_fd_sc_hd__a211o_1
XFILLER_0_127_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14503_ _04446_ _04510_ VGND VGND VPWR VPWR _04512_ sky130_fd_sc_hd__nor2_1
X_11715_ _01651_ _01653_ _01617_ VGND VGND VPWR VPWR _01654_ sky130_fd_sc_hd__and3b_1
XFILLER_0_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15483_ _05515_ _05588_ VGND VGND VPWR VPWR _05590_ sky130_fd_sc_hd__and2_1
X_18271_ net281 _06379_ VGND VGND VPWR VPWR _08656_ sky130_fd_sc_hd__nand2_1
X_12695_ _02553_ _02633_ VGND VGND VPWR VPWR _02634_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17222_ _07500_ _07501_ VGND VGND VPWR VPWR _07502_ sky130_fd_sc_hd__nor2_1
X_14434_ _04341_ _04435_ VGND VGND VPWR VPWR _04436_ sky130_fd_sc_hd__nand2_1
X_11646_ _01521_ _01584_ VGND VGND VPWR VPWR _01585_ sky130_fd_sc_hd__xor2_1
Xinput14 measurement[3] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_1
XFILLER_0_126_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17153_ _07407_ _07420_ VGND VGND VPWR VPWR _07427_ sky130_fd_sc_hd__or2b_1
XFILLER_0_142_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14365_ _04350_ _04356_ _04359_ VGND VGND VPWR VPWR _04360_ sky130_fd_sc_hd__a21oi_2
Xinput25 reg_addr[13] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
Xinput36 reg_addr[6] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
X_11577_ _01513_ _01515_ VGND VGND VPWR VPWR _01516_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput47 reg_data[16] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput58 reg_data[9] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_4
X_13316_ _03180_ _03266_ VGND VGND VPWR VPWR _03269_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16104_ prev_error\[7\] _09577_ VGND VGND VPWR VPWR _06273_ sky130_fd_sc_hd__or2_2
Xinput69 target[18] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dlymetal6s2s_1
X_10528_ net388 _04885_ _00363_ VGND VGND VPWR VPWR _00467_ sky130_fd_sc_hd__a21oi_1
X_17084_ _07346_ _07347_ _07350_ VGND VGND VPWR VPWR _07351_ sky130_fd_sc_hd__nand3_2
X_14296_ _03986_ _04255_ _04230_ _04254_ VGND VGND VPWR VPWR _04284_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16035_ _08669_ _08680_ _08702_ _08724_ VGND VGND VPWR VPWR _06197_ sky130_fd_sc_hd__o31a_1
XFILLER_0_0_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13247_ _03118_ _03199_ VGND VGND VPWR VPWR _03200_ sky130_fd_sc_hd__or2_1
X_10459_ net565 _08185_ VGND VGND VPWR VPWR _00398_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13178_ _03129_ _03057_ VGND VGND VPWR VPWR _03130_ sky130_fd_sc_hd__or2_1
X_12129_ _02052_ _02066_ VGND VGND VPWR VPWR _02068_ sky130_fd_sc_hd__or2_1
X_17986_ _08337_ _08341_ _08342_ VGND VGND VPWR VPWR _08343_ sky130_fd_sc_hd__or3_2
X_16937_ _07187_ _07188_ VGND VGND VPWR VPWR _07189_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16868_ _07110_ _07112_ VGND VGND VPWR VPWR _07113_ sky130_fd_sc_hd__or2b_1
X_18607_ _08905_ VGND VGND VPWR VPWR _09026_ sky130_fd_sc_hd__inv_2
X_15819_ _04893_ _05958_ VGND VGND VPWR VPWR _05959_ sky130_fd_sc_hd__or2_1
X_16799_ _06937_ _07036_ VGND VGND VPWR VPWR _07037_ sky130_fd_sc_hd__xnor2_1
X_18538_ _08893_ _08739_ net525 net521 VGND VGND VPWR VPWR _08950_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18469_ net530 _08870_ _08872_ VGND VGND VPWR VPWR _08874_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09607_ _03091_ VGND VGND VPWR VPWR _03102_ sky130_fd_sc_hd__buf_2
XFILLER_0_78_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Left_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11500_ _01379_ _01433_ _01436_ VGND VGND VPWR VPWR _01439_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12480_ _02332_ VGND VGND VPWR VPWR _02419_ sky130_fd_sc_hd__inv_2
X_11431_ _01325_ _01327_ _01328_ _01323_ VGND VGND VPWR VPWR _01370_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_105_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14150_ _04084_ _04103_ _04121_ VGND VGND VPWR VPWR _04123_ sky130_fd_sc_hd__nand3_1
X_11362_ net358 _00815_ _01234_ VGND VGND VPWR VPWR _01301_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13101_ _03043_ _03044_ VGND VGND VPWR VPWR _03045_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10313_ _00228_ _00237_ _00251_ VGND VGND VPWR VPWR _00252_ sky130_fd_sc_hd__nor3_1
X_14081_ net408 net144 _04049_ _04052_ VGND VGND VPWR VPWR _04053_ sky130_fd_sc_hd__o2bb2a_1
X_11293_ net366 net362 _00514_ _00613_ VGND VGND VPWR VPWR _01232_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_60_Left_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13032_ _02969_ _02970_ VGND VGND VPWR VPWR _02971_ sky130_fd_sc_hd__nand2_1
X_10244_ _07734_ _08493_ VGND VGND VPWR VPWR _00183_ sky130_fd_sc_hd__xor2_1
X_17840_ _08176_ _08181_ VGND VGND VPWR VPWR _08182_ sky130_fd_sc_hd__xnor2_1
X_10175_ _09252_ _09263_ VGND VGND VPWR VPWR _09274_ sky130_fd_sc_hd__nand2_1
X_17771_ net301 _07183_ _08094_ _08092_ VGND VGND VPWR VPWR _08106_ sky130_fd_sc_hd__a31o_1
Xfanout180 kd_2\[4\] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_2
X_14983_ _05037_ _05038_ net437 net177 VGND VGND VPWR VPWR _05040_ sky130_fd_sc_hd__and4bb_1
Xfanout191 net192 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__buf_2
X_16722_ _06944_ _06946_ VGND VGND VPWR VPWR _06952_ sky130_fd_sc_hd__xor2_1
X_13934_ _03902_ _03904_ VGND VGND VPWR VPWR _03905_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16653_ _06855_ _06872_ _06874_ VGND VGND VPWR VPWR _06877_ sky130_fd_sc_hd__or3_1
X_13865_ _03820_ _03830_ VGND VGND VPWR VPWR _03831_ sky130_fd_sc_hd__nand2_1
X_15604_ _05719_ _05722_ VGND VGND VPWR VPWR _05723_ sky130_fd_sc_hd__nand2_1
X_12816_ _02741_ _02743_ _02754_ VGND VGND VPWR VPWR _02755_ sky130_fd_sc_hd__a21bo_1
X_16584_ _06800_ VGND VGND VPWR VPWR _06801_ sky130_fd_sc_hd__clkbuf_4
X_13796_ net256 _02913_ VGND VGND VPWR VPWR _03762_ sky130_fd_sc_hd__nand2_2
XFILLER_0_56_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18323_ _08708_ _08712_ VGND VGND VPWR VPWR _08714_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15535_ _05641_ _05646_ VGND VGND VPWR VPWR _05647_ sky130_fd_sc_hd__and2_1
X_12747_ net259 _01798_ _02684_ _02685_ VGND VGND VPWR VPWR _02686_ sky130_fd_sc_hd__and4_1
XFILLER_0_57_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18254_ _08633_ _08637_ VGND VGND VPWR VPWR _08638_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12678_ net231 _01853_ _01874_ net227 VGND VGND VPWR VPWR _02617_ sky130_fd_sc_hd__a22o_1
X_15466_ net452 net457 net185 net180 VGND VGND VPWR VPWR _05571_ sky130_fd_sc_hd__and4_1
XFILLER_0_5_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17205_ net328 _06401_ _07482_ _07483_ VGND VGND VPWR VPWR _07484_ sky130_fd_sc_hd__a31oi_2
X_14417_ _04414_ _04416_ VGND VGND VPWR VPWR _04417_ sky130_fd_sc_hd__and2b_1
X_11629_ _01565_ _01567_ VGND VGND VPWR VPWR _01568_ sky130_fd_sc_hd__xnor2_1
X_18185_ _08434_ _08561_ i_error\[1\] VGND VGND VPWR VPWR _08562_ sky130_fd_sc_hd__a21o_1
X_15397_ net449 net184 VGND VGND VPWR VPWR _05495_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17136_ _07379_ _07366_ VGND VGND VPWR VPWR _07408_ sky130_fd_sc_hd__or2b_1
XFILLER_0_80_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14348_ _04337_ _04338_ _04340_ VGND VGND VPWR VPWR _04341_ sky130_fd_sc_hd__or3_1
X_14279_ net411 net160 net156 net416 VGND VGND VPWR VPWR _04265_ sky130_fd_sc_hd__a22oi_1
X_17067_ _07328_ _07330_ _07331_ VGND VGND VPWR VPWR _07332_ sky130_fd_sc_hd__or3_1
X_16018_ _08097_ _05754_ VGND VGND VPWR VPWR _06178_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17969_ net322 net318 _07181_ _07567_ VGND VGND VPWR VPWR _08324_ sky130_fd_sc_hd__and4_1
XFILLER_0_109_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_108_Left_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_117_Left_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_126_Left_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11980_ _01896_ _01903_ _01918_ VGND VGND VPWR VPWR _01919_ sky130_fd_sc_hd__and3_1
X_10931_ _00674_ _05930_ VGND VGND VPWR VPWR _00870_ sky130_fd_sc_hd__nor2_1
X_13650_ net269 VGND VGND VPWR VPWR _03611_ sky130_fd_sc_hd__inv_2
X_10862_ _00799_ _00800_ VGND VGND VPWR VPWR _00801_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12601_ _02534_ _02537_ _02539_ VGND VGND VPWR VPWR _02540_ sky130_fd_sc_hd__o21ai_1
X_13581_ _03480_ _03483_ _03482_ VGND VGND VPWR VPWR _03540_ sky130_fd_sc_hd__a21o_1
X_10793_ net393 net509 _05369_ VGND VGND VPWR VPWR _00732_ sky130_fd_sc_hd__and3_1
XFILLER_0_137_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12532_ _02423_ _02457_ VGND VGND VPWR VPWR _02471_ sky130_fd_sc_hd__xnor2_2
X_15320_ _05405_ _05407_ _05409_ VGND VGND VPWR VPWR _05410_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_135_Left_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12463_ net201 _02332_ _02333_ VGND VGND VPWR VPWR _02402_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15251_ _05321_ _05333_ VGND VGND VPWR VPWR _05334_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14202_ _04178_ _04179_ VGND VGND VPWR VPWR _04180_ sky130_fd_sc_hd__nand2_1
X_11414_ _01343_ _01342_ _01314_ VGND VGND VPWR VPWR _01353_ sky130_fd_sc_hd__a21oi_1
X_15182_ _05247_ _05252_ _05256_ _05257_ VGND VGND VPWR VPWR _05258_ sky130_fd_sc_hd__o211ai_2
X_12394_ _02324_ _02325_ VGND VGND VPWR VPWR _02333_ sky130_fd_sc_hd__xor2_1
X_14133_ _04051_ _04048_ _04053_ VGND VGND VPWR VPWR _04105_ sky130_fd_sc_hd__or3_1
X_11345_ _01221_ _01283_ VGND VGND VPWR VPWR _01284_ sky130_fd_sc_hd__xnor2_1
X_18941_ net201 _01817_ _09290_ _09392_ VGND VGND VPWR VPWR _09393_ sky130_fd_sc_hd__a31o_1
X_14064_ _04034_ _04009_ _04012_ VGND VGND VPWR VPWR _04036_ sky130_fd_sc_hd__and3_1
X_11276_ net386 _08185_ _06051_ net406 VGND VGND VPWR VPWR _01215_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13015_ _02953_ _02785_ VGND VGND VPWR VPWR _02954_ sky130_fd_sc_hd__xnor2_1
X_10227_ _09274_ _09406_ VGND VGND VPWR VPWR _00166_ sky130_fd_sc_hd__xnor2_2
X_18872_ _09308_ _09315_ VGND VGND VPWR VPWR _09317_ sky130_fd_sc_hd__nand2_1
X_17823_ _08052_ _08158_ _08162_ VGND VGND VPWR VPWR _08164_ sky130_fd_sc_hd__nor3_1
X_10158_ _06788_ _07712_ _07701_ VGND VGND VPWR VPWR _09087_ sky130_fd_sc_hd__a21oi_1
X_17754_ _08085_ _08087_ VGND VGND VPWR VPWR _08088_ sky130_fd_sc_hd__nor2_1
X_10089_ _06656_ _06678_ VGND VGND VPWR VPWR _08328_ sky130_fd_sc_hd__xor2_1
X_14966_ net478 net131 _04960_ _04964_ VGND VGND VPWR VPWR _05021_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_89_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16705_ _06837_ _06933_ VGND VGND VPWR VPWR _06934_ sky130_fd_sc_hd__nand2_1
X_13917_ _02354_ _03885_ VGND VGND VPWR VPWR _03886_ sky130_fd_sc_hd__and2_1
X_17685_ _07905_ _07906_ _07918_ VGND VGND VPWR VPWR _08012_ sky130_fd_sc_hd__o21ai_1
X_14897_ _04871_ _04872_ VGND VGND VPWR VPWR _04945_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16636_ net293 _06410_ VGND VGND VPWR VPWR _06858_ sky130_fd_sc_hd__nand2_1
X_13848_ _03810_ _03812_ VGND VGND VPWR VPWR _03814_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16567_ _06772_ _06776_ _06781_ VGND VGND VPWR VPWR _06782_ sky130_fd_sc_hd__a21oi_2
X_13779_ _03690_ _03702_ _03701_ VGND VGND VPWR VPWR _03745_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18306_ net281 _06379_ _08659_ _06561_ VGND VGND VPWR VPWR _08695_ sky130_fd_sc_hd__a31o_1
X_15518_ _05617_ _05619_ _05621_ VGND VGND VPWR VPWR _05628_ sky130_fd_sc_hd__or3_1
XFILLER_0_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19286_ clknet_4_7_0_clock _00064_ VGND VGND VPWR VPWR kp\[16\] sky130_fd_sc_hd__dfxtp_2
X_16498_ _06642_ _06705_ VGND VGND VPWR VPWR _06706_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18237_ _06261_ _08618_ VGND VGND VPWR VPWR _08619_ sky130_fd_sc_hd__or2b_1
XFILLER_0_26_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15449_ _05550_ _05551_ net479 net164 VGND VGND VPWR VPWR _05552_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_127_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18168_ _08441_ _08491_ VGND VGND VPWR VPWR _08543_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_5_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap100 _08896_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__buf_1
XFILLER_0_20_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17119_ _07354_ _07356_ VGND VGND VPWR VPWR _07389_ sky130_fd_sc_hd__and2b_1
XFILLER_0_40_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18099_ _07769_ _07780_ VGND VGND VPWR VPWR _08467_ sky130_fd_sc_hd__and2b_1
XFILLER_0_123_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09941_ _06513_ _06535_ VGND VGND VPWR VPWR _06700_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09872_ net568 _05930_ VGND VGND VPWR VPWR _05941_ sky130_fd_sc_hd__nand2_2
XFILLER_0_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11130_ net383 _06634_ _01055_ VGND VGND VPWR VPWR _01069_ sky130_fd_sc_hd__and3_1
X_11061_ _00889_ _00999_ VGND VGND VPWR VPWR _01000_ sky130_fd_sc_hd__nor2_1
X_10012_ _07437_ _07470_ VGND VGND VPWR VPWR _07481_ sky130_fd_sc_hd__xnor2_1
X_14820_ net436 net174 _04558_ VGND VGND VPWR VPWR _04860_ sky130_fd_sc_hd__and3_1
X_14751_ _04782_ _04783_ VGND VGND VPWR VPWR _04784_ sky130_fd_sc_hd__or2b_1
X_11963_ _01877_ _01901_ VGND VGND VPWR VPWR _01902_ sky130_fd_sc_hd__and2_1
X_13702_ _03554_ _03608_ _03549_ VGND VGND VPWR VPWR _03668_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_157_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10914_ _00831_ _00832_ _00848_ _00852_ VGND VGND VPWR VPWR _00853_ sky130_fd_sc_hd__o211ai_4
X_17470_ _07699_ _07707_ _07774_ VGND VGND VPWR VPWR _07775_ sky130_fd_sc_hd__a21boi_2
X_11894_ _01827_ _01831_ VGND VGND VPWR VPWR _01833_ sky130_fd_sc_hd__xor2_1
X_14682_ _04496_ _04707_ VGND VGND VPWR VPWR _04708_ sky130_fd_sc_hd__xor2_1
X_16421_ _06620_ VGND VGND VPWR VPWR _06621_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13633_ _03588_ _03580_ _03586_ VGND VGND VPWR VPWR _03593_ sky130_fd_sc_hd__or3_1
X_10845_ _00778_ _00783_ VGND VGND VPWR VPWR _00784_ sky130_fd_sc_hd__or2b_1
XPHY_EDGE_ROW_143_Left_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19140_ net504 i_error\[11\] VGND VGND VPWR VPWR _09563_ sky130_fd_sc_hd__or2_1
X_16352_ _06364_ _06362_ _06324_ VGND VGND VPWR VPWR _06545_ sky130_fd_sc_hd__and3b_1
XFILLER_0_26_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13564_ _03518_ _03521_ _03522_ _03517_ _03515_ VGND VGND VPWR VPWR _03523_ sky130_fd_sc_hd__a32o_1
XFILLER_0_82_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10776_ _00710_ _00714_ VGND VGND VPWR VPWR _00715_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15303_ net468 net486 net162 net144 VGND VGND VPWR VPWR _05392_ sky130_fd_sc_hd__and4_1
X_12515_ _02304_ _02453_ VGND VGND VPWR VPWR _02454_ sky130_fd_sc_hd__nand2_1
X_19071_ _09515_ _09519_ VGND VGND VPWR VPWR _00092_ sky130_fd_sc_hd__nor2_1
X_16283_ _06468_ VGND VGND VPWR VPWR _06470_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_136_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13495_ _03447_ _03451_ _03453_ VGND VGND VPWR VPWR _03454_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18022_ _08360_ _08369_ VGND VGND VPWR VPWR _08382_ sky130_fd_sc_hd__nor2_1
X_12446_ _02381_ _02384_ VGND VGND VPWR VPWR _02385_ sky130_fd_sc_hd__nor2_1
X_15234_ _05308_ _05304_ _05306_ VGND VGND VPWR VPWR _05316_ sky130_fd_sc_hd__or3_1
XFILLER_0_124_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12377_ net219 net214 _01853_ _01874_ VGND VGND VPWR VPWR _02316_ sky130_fd_sc_hd__and4_1
XFILLER_0_23_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15165_ _05225_ _05239_ VGND VGND VPWR VPWR _05240_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14116_ _03921_ _04087_ VGND VGND VPWR VPWR _04088_ sky130_fd_sc_hd__and2_1
X_11328_ _01250_ _01251_ _01264_ VGND VGND VPWR VPWR _01267_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_152_Left_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15096_ _05139_ _05123_ _05135_ VGND VGND VPWR VPWR _05164_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18924_ _09371_ _09374_ VGND VGND VPWR VPWR _09375_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_157_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14047_ _04014_ _03997_ _04003_ VGND VGND VPWR VPWR _04019_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11259_ _01192_ _01195_ _01196_ _01197_ VGND VGND VPWR VPWR _01198_ sky130_fd_sc_hd__a211o_2
X_18855_ _02134_ _09286_ _09298_ VGND VGND VPWR VPWR _09299_ sky130_fd_sc_hd__a21oi_1
X_17806_ _08134_ _08144_ VGND VGND VPWR VPWR _08145_ sky130_fd_sc_hd__and2b_1
X_18786_ _04115_ _09215_ _09218_ _09222_ VGND VGND VPWR VPWR _09223_ sky130_fd_sc_hd__or4b_4
X_15998_ _01209_ _01210_ VGND VGND VPWR VPWR _06156_ sky130_fd_sc_hd__and2b_2
X_17737_ net313 _07094_ _08066_ _08067_ VGND VGND VPWR VPWR _08069_ sky130_fd_sc_hd__a22o_1
X_14949_ _04990_ _05001_ VGND VGND VPWR VPWR _05002_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17668_ _07890_ _07892_ VGND VGND VPWR VPWR _07993_ sky130_fd_sc_hd__xor2_1
XFILLER_0_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16619_ _06823_ _06824_ VGND VGND VPWR VPWR _06839_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17599_ _07912_ _07915_ VGND VGND VPWR VPWR _07917_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19338_ clknet_4_2_0_clock _00021_ VGND VGND VPWR VPWR kd_2\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19269_ clknet_4_11_0_clock _00151_ VGND VGND VPWR VPWR prev_d_error\[18\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_155_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09924_ net353 _05336_ _05380_ _06502_ VGND VGND VPWR VPWR _06513_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09855_ _05424_ VGND VGND VPWR VPWR _05754_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09786_ _04984_ VGND VGND VPWR VPWR _04995_ sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_134_Right_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10630_ net384 _05413_ _00566_ _00568_ VGND VGND VPWR VPWR _00569_ sky130_fd_sc_hd__a31o_1
XFILLER_0_48_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10561_ _00497_ _00499_ VGND VGND VPWR VPWR _00500_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_11_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12300_ _02237_ _02238_ VGND VGND VPWR VPWR _02239_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13280_ _03154_ _03232_ VGND VGND VPWR VPWR _03233_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10492_ _00299_ _00430_ VGND VGND VPWR VPWR _00431_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12231_ _02168_ _02169_ VGND VGND VPWR VPWR _02170_ sky130_fd_sc_hd__xor2_1
XFILLER_0_106_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12162_ _02099_ _02100_ VGND VGND VPWR VPWR _02101_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11113_ _00966_ _01046_ _01051_ VGND VGND VPWR VPWR _01052_ sky130_fd_sc_hd__nand3_1
XFILLER_0_130_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12093_ _02025_ _02031_ VGND VGND VPWR VPWR _02032_ sky130_fd_sc_hd__and2_1
X_16970_ net311 _06409_ _06401_ net308 VGND VGND VPWR VPWR _07225_ sky130_fd_sc_hd__a22o_1
X_15921_ _05467_ _05949_ VGND VGND VPWR VPWR _06071_ sky130_fd_sc_hd__nand2_1
X_11044_ net378 _06612_ _00982_ VGND VGND VPWR VPWR _00983_ sky130_fd_sc_hd__a21o_1
X_18640_ _06110_ _09061_ VGND VGND VPWR VPWR _09062_ sky130_fd_sc_hd__nand2_2
X_15852_ _05990_ _05993_ _04480_ VGND VGND VPWR VPWR _05995_ sky130_fd_sc_hd__o21a_1
X_14803_ _04823_ _04818_ VGND VGND VPWR VPWR _04842_ sky130_fd_sc_hd__or2b_1
X_18571_ _06019_ _06123_ VGND VGND VPWR VPWR _08986_ sky130_fd_sc_hd__or2_2
X_15783_ _05915_ _05916_ _05870_ _05918_ VGND VGND VPWR VPWR _05920_ sky130_fd_sc_hd__and4b_1
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12995_ _02933_ VGND VGND VPWR VPWR _02934_ sky130_fd_sc_hd__clkbuf_4
X_17522_ _07827_ _07831_ VGND VGND VPWR VPWR _07832_ sky130_fd_sc_hd__or2_1
X_14734_ _04760_ _04762_ _04765_ VGND VGND VPWR VPWR _04766_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_87_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11946_ net203 _01836_ _01808_ net205 VGND VGND VPWR VPWR _01885_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17453_ _07754_ _07755_ VGND VGND VPWR VPWR _07757_ sky130_fd_sc_hd__xnor2_1
X_14665_ net465 net129 _04482_ VGND VGND VPWR VPWR _04690_ sky130_fd_sc_hd__and3_1
X_11877_ net213 _01810_ _01815_ VGND VGND VPWR VPWR _01816_ sky130_fd_sc_hd__and3_1
XFILLER_0_157_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16404_ net293 _06386_ _06602_ _06599_ VGND VGND VPWR VPWR _06603_ sky130_fd_sc_hd__a31o_1
X_13616_ net260 _02330_ _02408_ net256 VGND VGND VPWR VPWR _03575_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_27_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17384_ _07676_ _07680_ VGND VGND VPWR VPWR _07681_ sky130_fd_sc_hd__xnor2_1
X_10828_ _00676_ _00764_ _00766_ VGND VGND VPWR VPWR _00767_ sky130_fd_sc_hd__a21bo_1
X_14596_ net470 net475 net125 net121 VGND VGND VPWR VPWR _04614_ sky130_fd_sc_hd__and4_1
X_19123_ net503 i_error\[3\] VGND VGND VPWR VPWR _09553_ sky130_fd_sc_hd__or2_1
X_16335_ _06525_ _06508_ _06509_ VGND VGND VPWR VPWR _06527_ sky130_fd_sc_hd__nor3_1
X_13547_ _03502_ _03503_ _03505_ VGND VGND VPWR VPWR _03506_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10759_ _00601_ _00697_ VGND VGND VPWR VPWR _00698_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19054_ _04126_ net81 VGND VGND VPWR VPWR _09508_ sky130_fd_sc_hd__and2_1
X_16266_ _06397_ _06450_ VGND VGND VPWR VPWR _06451_ sky130_fd_sc_hd__xnor2_1
X_13478_ net239 _02544_ VGND VGND VPWR VPWR _03437_ sky130_fd_sc_hd__nand2_1
X_18005_ _08362_ _08363_ VGND VGND VPWR VPWR _08364_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15217_ _05291_ _05296_ VGND VGND VPWR VPWR _05297_ sky130_fd_sc_hd__or2_1
X_12429_ _02267_ _02266_ VGND VGND VPWR VPWR _02368_ sky130_fd_sc_hd__and2b_1
XFILLER_0_113_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16197_ _06373_ _06374_ VGND VGND VPWR VPWR _06375_ sky130_fd_sc_hd__and2_1
X_15148_ _05213_ _05220_ VGND VGND VPWR VPWR _05221_ sky130_fd_sc_hd__and2_1
X_15079_ net437 net177 _05037_ _05038_ VGND VGND VPWR VPWR _05145_ sky130_fd_sc_hd__o2bb2a_1
X_18907_ _09209_ _09213_ _09223_ _09355_ VGND VGND VPWR VPWR _09356_ sky130_fd_sc_hd__or4b_4
X_09640_ net53 _03358_ _03391_ net253 VGND VGND VPWR VPWR _00013_ sky130_fd_sc_hd__a22o_1
X_18838_ _02121_ _02141_ _09279_ VGND VGND VPWR VPWR _09280_ sky130_fd_sc_hd__a21bo_1
X_18769_ _08985_ _08995_ VGND VGND VPWR VPWR _09204_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09907_ _06304_ _06315_ VGND VGND VPWR VPWR _06326_ sky130_fd_sc_hd__or2b_1
X_09838_ net380 net376 VGND VGND VPWR VPWR _05567_ sky130_fd_sc_hd__or2_1
X_09769_ net67 net9 VGND VGND VPWR VPWR _04808_ sky130_fd_sc_hd__and2b_1
X_11800_ _01705_ _01706_ _01737_ _06073_ _01738_ VGND VGND VPWR VPWR _01739_ sky130_fd_sc_hd__a32o_2
X_12780_ net222 _01909_ _02616_ _02617_ VGND VGND VPWR VPWR _02719_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11731_ _01461_ _01507_ _01668_ _01669_ VGND VGND VPWR VPWR _01670_ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14450_ _04443_ _04446_ _04448_ VGND VGND VPWR VPWR _04453_ sky130_fd_sc_hd__or3_1
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11662_ _01558_ _01596_ _01599_ VGND VGND VPWR VPWR _01601_ sky130_fd_sc_hd__and3_1
XFILLER_0_83_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13401_ _02989_ _03355_ VGND VGND VPWR VPWR _03356_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10613_ _00550_ _00551_ VGND VGND VPWR VPWR _00552_ sky130_fd_sc_hd__nor2_2
X_14381_ _04375_ _04376_ VGND VGND VPWR VPWR _04377_ sky130_fd_sc_hd__or2_1
X_11593_ _01488_ _01531_ VGND VGND VPWR VPWR _01532_ sky130_fd_sc_hd__xnor2_1
X_16120_ prev_error\[10\] _05897_ _06150_ VGND VGND VPWR VPWR _06290_ sky130_fd_sc_hd__and3_1
X_13332_ _03282_ _03284_ VGND VGND VPWR VPWR _03285_ sky130_fd_sc_hd__or2b_1
X_10544_ _00481_ _00482_ VGND VGND VPWR VPWR _00483_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_122_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16051_ _06212_ _06213_ VGND VGND VPWR VPWR _06214_ sky130_fd_sc_hd__xnor2_1
X_13263_ _03198_ _03200_ _03215_ VGND VGND VPWR VPWR _03216_ sky130_fd_sc_hd__o21a_1
X_10475_ _00399_ _00402_ _00404_ VGND VGND VPWR VPWR _00414_ sky130_fd_sc_hd__or3_1
X_15002_ _05036_ _05059_ VGND VGND VPWR VPWR _05060_ sky130_fd_sc_hd__nor2_1
X_12214_ net223 _01932_ _01990_ VGND VGND VPWR VPWR _02153_ sky130_fd_sc_hd__a21o_2
X_13194_ net260 net257 _01851_ _01859_ VGND VGND VPWR VPWR _03147_ sky130_fd_sc_hd__and4_1
X_12145_ _01912_ _02083_ VGND VGND VPWR VPWR _02084_ sky130_fd_sc_hd__or2_1
X_16953_ net282 _06993_ _07176_ VGND VGND VPWR VPWR _07207_ sky130_fd_sc_hd__a21o_1
X_12076_ _01978_ _02013_ _02014_ VGND VGND VPWR VPWR _02015_ sky130_fd_sc_hd__o21ai_1
X_15904_ _05957_ _06052_ VGND VGND VPWR VPWR _06053_ sky130_fd_sc_hd__and2_1
X_11027_ _00964_ _08735_ _00963_ _00965_ VGND VGND VPWR VPWR _00966_ sky130_fd_sc_hd__or4_1
X_16884_ _07016_ _07021_ _06542_ VGND VGND VPWR VPWR _07131_ sky130_fd_sc_hd__a21o_1
X_18623_ _09034_ _09040_ _09042_ VGND VGND VPWR VPWR _09044_ sky130_fd_sc_hd__or3_1
X_15835_ _04581_ _04678_ _04677_ VGND VGND VPWR VPWR _05977_ sky130_fd_sc_hd__a21oi_1
X_18554_ _01698_ _08967_ VGND VGND VPWR VPWR _08968_ sky130_fd_sc_hd__or2b_1
X_15766_ net483 net183 VGND VGND VPWR VPWR _05901_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12978_ _02853_ _02855_ VGND VGND VPWR VPWR _02917_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17505_ _07810_ _07813_ VGND VGND VPWR VPWR _07814_ sky130_fd_sc_hd__or2b_1
X_14717_ _04721_ _04744_ _04746_ VGND VGND VPWR VPWR _04747_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_157_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11929_ _01856_ _01866_ VGND VGND VPWR VPWR _01868_ sky130_fd_sc_hd__xnor2_1
X_18485_ _06173_ _06131_ VGND VGND VPWR VPWR _08892_ sky130_fd_sc_hd__and2b_1
X_15697_ _05822_ _05824_ VGND VGND VPWR VPWR _05825_ sky130_fd_sc_hd__nand2_1
X_17436_ _07676_ _07680_ VGND VGND VPWR VPWR _07738_ sky130_fd_sc_hd__or2b_1
X_14648_ _04650_ _04651_ _04653_ VGND VGND VPWR VPWR _04671_ sky130_fd_sc_hd__o21ba_1
XANTENNA_17 net330 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_28 net539 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17367_ net281 _02932_ _07661_ VGND VGND VPWR VPWR _07662_ sky130_fd_sc_hd__and3_1
X_14579_ _04584_ _04585_ VGND VGND VPWR VPWR _04595_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19106_ net499 prev_error\[14\] VGND VGND VPWR VPWR _09542_ sky130_fd_sc_hd__or2_1
X_16318_ _06417_ _06423_ VGND VGND VPWR VPWR _06508_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17298_ _07584_ _07585_ VGND VGND VPWR VPWR _07586_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19037_ _09448_ _09485_ _09465_ VGND VGND VPWR VPWR _09495_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16249_ _06273_ _02087_ _06287_ _06292_ _06291_ VGND VGND VPWR VPWR _06432_ sky130_fd_sc_hd__a311o_1
XFILLER_0_125_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09623_ net43 _03091_ _03124_ net142 VGND VGND VPWR VPWR _00022_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10260_ _00189_ _00198_ VGND VGND VPWR VPWR _00199_ sky130_fd_sc_hd__and2b_1
X_10191_ _09252_ _09417_ _09439_ VGND VGND VPWR VPWR _09450_ sky130_fd_sc_hd__a21o_1
XFILLER_0_100_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout340 kp\[16\] VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__clkbuf_4
Xfanout351 kp\[13\] VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__clkbuf_4
Xfanout362 kp\[10\] VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__clkbuf_4
X_13950_ net434 net123 VGND VGND VPWR VPWR _03922_ sky130_fd_sc_hd__nand2_1
Xfanout373 kp\[8\] VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__clkbuf_4
Xfanout384 kp\[5\] VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__clkbuf_4
Xfanout395 net398 VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__dlymetal6s2s_1
X_12901_ _02837_ _02839_ VGND VGND VPWR VPWR _02840_ sky130_fd_sc_hd__xnor2_1
X_13881_ _03610_ _03665_ _03845_ _03846_ VGND VGND VPWR VPWR _03847_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15620_ _05738_ _05739_ net478 net176 VGND VGND VPWR VPWR _05740_ sky130_fd_sc_hd__and4bb_2
X_12832_ _02676_ _02768_ VGND VGND VPWR VPWR _02771_ sky130_fd_sc_hd__and2_1
X_15551_ _05659_ _05662_ _05663_ VGND VGND VPWR VPWR _05664_ sky130_fd_sc_hd__and3_1
X_12763_ _02700_ _02701_ VGND VGND VPWR VPWR _02702_ sky130_fd_sc_hd__xor2_1
XFILLER_0_139_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14502_ net420 net161 _04443_ _04444_ VGND VGND VPWR VPWR _04510_ sky130_fd_sc_hd__o2bb2a_1
X_11714_ _00439_ _00615_ _01638_ _00812_ net564 VGND VGND VPWR VPWR _01653_ sky130_fd_sc_hd__o2111a_1
X_18270_ net292 _06325_ VGND VGND VPWR VPWR _08655_ sky130_fd_sc_hd__and2_1
X_15482_ net432 net197 _05514_ VGND VGND VPWR VPWR _05588_ sky130_fd_sc_hd__a21o_1
XFILLER_0_83_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12694_ _02550_ _02552_ VGND VGND VPWR VPWR _02633_ sky130_fd_sc_hd__or2_1
X_17221_ net308 _06721_ _06802_ net305 VGND VGND VPWR VPWR _07501_ sky130_fd_sc_hd__a22oi_1
X_14433_ _04337_ _04338_ _04340_ VGND VGND VPWR VPWR _04435_ sky130_fd_sc_hd__o21ai_1
X_11645_ _01580_ _01583_ VGND VGND VPWR VPWR _01584_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17152_ _07278_ _07423_ _07424_ VGND VGND VPWR VPWR _07425_ sky130_fd_sc_hd__a21oi_2
X_14364_ _04270_ _04358_ VGND VGND VPWR VPWR _04359_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput15 measurement[4] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_1
XFILLER_0_24_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput26 reg_addr[14] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
X_11576_ _01471_ _01514_ VGND VGND VPWR VPWR _01515_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput37 reg_addr[7] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput48 reg_data[17] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_4
X_16103_ prev_error\[15\] _05171_ _06270_ VGND VGND VPWR VPWR _06272_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_3_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13315_ _03177_ _03179_ _03267_ VGND VGND VPWR VPWR _03268_ sky130_fd_sc_hd__nand3_2
Xinput59 reset VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_1
X_17083_ _07210_ _07348_ VGND VGND VPWR VPWR _07350_ sky130_fd_sc_hd__xor2_2
XFILLER_0_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10527_ _00429_ _00457_ VGND VGND VPWR VPWR _00466_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14295_ _04279_ _04281_ _04273_ _04277_ VGND VGND VPWR VPWR _04283_ sky130_fd_sc_hd__a211o_1
X_16034_ _06177_ _06195_ VGND VGND VPWR VPWR _06196_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13246_ _03115_ _03117_ VGND VGND VPWR VPWR _03199_ sky130_fd_sc_hd__nor2_1
X_10458_ _00322_ VGND VGND VPWR VPWR _00397_ sky130_fd_sc_hd__inv_2
XFILLER_0_149_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13177_ kd_1\[12\] _02746_ VGND VGND VPWR VPWR _03129_ sky130_fd_sc_hd__nand2_1
X_10389_ _00247_ _00320_ _00327_ VGND VGND VPWR VPWR _00328_ sky130_fd_sc_hd__a21o_1
X_12128_ _02052_ _02066_ VGND VGND VPWR VPWR _02067_ sky130_fd_sc_hd__nand2_1
X_17985_ _08336_ _08331_ _08335_ VGND VGND VPWR VPWR _08342_ sky130_fd_sc_hd__nor3_1
X_16936_ _07178_ _07179_ VGND VGND VPWR VPWR _07188_ sky130_fd_sc_hd__xor2_1
X_12059_ _01996_ _01997_ VGND VGND VPWR VPWR _01998_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16867_ _07084_ _07111_ VGND VGND VPWR VPWR _07112_ sky130_fd_sc_hd__and2_1
X_15818_ _04892_ _04887_ _04891_ VGND VGND VPWR VPWR _05958_ sky130_fd_sc_hd__and3_1
X_18606_ _06115_ _06041_ _06114_ VGND VGND VPWR VPWR _09025_ sky130_fd_sc_hd__nand3_2
X_16798_ _07006_ _07034_ _07035_ VGND VGND VPWR VPWR _07036_ sky130_fd_sc_hd__a21oi_1
X_18537_ _08915_ _08948_ _08906_ VGND VGND VPWR VPWR _08949_ sky130_fd_sc_hd__a21oi_1
X_15749_ _05880_ _05881_ VGND VGND VPWR VPWR _05882_ sky130_fd_sc_hd__and2b_1
XFILLER_0_59_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18468_ _08686_ _08870_ _08872_ _08622_ _08615_ VGND VGND VPWR VPWR _08873_ sky130_fd_sc_hd__a32o_1
XFILLER_0_8_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17419_ _07201_ _07718_ VGND VGND VPWR VPWR _07719_ sky130_fd_sc_hd__xor2_1
XFILLER_0_7_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18399_ _08792_ _08794_ _08796_ _08620_ _06146_ VGND VGND VPWR VPWR _08797_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_90_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09606_ _03069_ _03080_ VGND VGND VPWR VPWR _03091_ sky130_fd_sc_hd__nor2_4
XFILLER_0_94_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11430_ _01364_ _01368_ VGND VGND VPWR VPWR _01369_ sky130_fd_sc_hd__xor2_2
XFILLER_0_151_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11361_ _01296_ _01298_ VGND VGND VPWR VPWR _01300_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13100_ _03042_ _03035_ VGND VGND VPWR VPWR _03044_ sky130_fd_sc_hd__and2b_1
X_10312_ _00249_ _00250_ VGND VGND VPWR VPWR _00251_ sky130_fd_sc_hd__and2_1
X_14080_ _04050_ VGND VGND VPWR VPWR _04052_ sky130_fd_sc_hd__inv_2
X_11292_ _01156_ _01230_ VGND VGND VPWR VPWR _01231_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10243_ _00177_ _00180_ _00181_ VGND VGND VPWR VPWR _00182_ sky130_fd_sc_hd__o21a_1
X_13031_ _02947_ _02966_ VGND VGND VPWR VPWR _02970_ sky130_fd_sc_hd__xor2_2
XFILLER_0_119_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10174_ _09164_ _09219_ _09241_ VGND VGND VPWR VPWR _09263_ sky130_fd_sc_hd__or3_1
X_17770_ _07991_ _08103_ _08102_ VGND VGND VPWR VPWR _08105_ sky130_fd_sc_hd__a21oi_1
X_14982_ net441 net173 net168 net446 VGND VGND VPWR VPWR _05038_ sky130_fd_sc_hd__a22oi_1
Xfanout170 net174 VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__buf_2
Xfanout181 net182 VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_4
Xfanout192 net194 VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_2
X_16721_ net306 _06386_ _06847_ _06950_ VGND VGND VPWR VPWR _06951_ sky130_fd_sc_hd__a31o_1
X_13933_ _03896_ _03901_ VGND VGND VPWR VPWR _03904_ sky130_fd_sc_hd__and2_1
X_16652_ _06855_ _06872_ _06874_ VGND VGND VPWR VPWR _06875_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13864_ _03818_ _03819_ VGND VGND VPWR VPWR _03830_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15603_ _05720_ VGND VGND VPWR VPWR _05722_ sky130_fd_sc_hd__inv_2
X_12815_ _02752_ _02753_ VGND VGND VPWR VPWR _02754_ sky130_fd_sc_hd__nand2_1
X_16583_ _02220_ _06798_ VGND VGND VPWR VPWR _06800_ sky130_fd_sc_hd__xnor2_4
X_13795_ net260 _02745_ VGND VGND VPWR VPWR _03761_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18322_ _08710_ _08711_ VGND VGND VPWR VPWR _08712_ sky130_fd_sc_hd__xnor2_1
X_15534_ _05640_ _05636_ _05638_ VGND VGND VPWR VPWR _05646_ sky130_fd_sc_hd__or3_1
X_12746_ net254 _01813_ net199 VGND VGND VPWR VPWR _02685_ sky130_fd_sc_hd__a21o_1
XFILLER_0_155_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18253_ _06514_ _08634_ _08635_ VGND VGND VPWR VPWR _08637_ sky130_fd_sc_hd__o21a_1
X_15465_ net452 net185 net179 net457 VGND VGND VPWR VPWR _05570_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_127_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12677_ _02613_ _02614_ _02507_ VGND VGND VPWR VPWR _02616_ sky130_fd_sc_hd__or3_1
XFILLER_0_154_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17204_ _07473_ _07480_ VGND VGND VPWR VPWR _07483_ sky130_fd_sc_hd__and2_1
X_14416_ _04321_ _04415_ VGND VGND VPWR VPWR _04416_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11628_ _01470_ _01566_ _01541_ VGND VGND VPWR VPWR _01567_ sky130_fd_sc_hd__a21oi_1
X_18184_ net513 _08433_ _08164_ _08430_ VGND VGND VPWR VPWR _08561_ sky130_fd_sc_hd__a211o_1
X_15396_ _05492_ _05493_ VGND VGND VPWR VPWR _05494_ sky130_fd_sc_hd__and2_1
XFILLER_0_114_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17135_ _07406_ _07192_ VGND VGND VPWR VPWR _07407_ sky130_fd_sc_hd__nor2_2
XFILLER_0_52_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14347_ _04318_ _04339_ VGND VGND VPWR VPWR _04340_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11559_ _01494_ _01497_ VGND VGND VPWR VPWR _01498_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17066_ _07319_ _07320_ _07326_ VGND VGND VPWR VPWR _07331_ sky130_fd_sc_hd__o21ba_1
X_14278_ net411 net416 net160 net156 VGND VGND VPWR VPWR _04264_ sky130_fd_sc_hd__and4_1
XFILLER_0_123_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16017_ _05666_ _08922_ _08944_ VGND VGND VPWR VPWR _06177_ sky130_fd_sc_hd__o21bai_2
X_13229_ net244 _02221_ VGND VGND VPWR VPWR _03182_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17968_ _08319_ _08322_ _08249_ VGND VGND VPWR VPWR _08323_ sky130_fd_sc_hd__a21oi_2
X_16919_ net271 _07095_ VGND VGND VPWR VPWR _07169_ sky130_fd_sc_hd__nand2_1
X_17899_ _08246_ _08195_ VGND VGND VPWR VPWR _08247_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10930_ net405 _04841_ _04852_ net387 _06062_ VGND VGND VPWR VPWR _00869_ sky130_fd_sc_hd__a32o_1
XFILLER_0_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10861_ net351 _00409_ _00324_ net357 VGND VGND VPWR VPWR _00800_ sky130_fd_sc_hd__a22oi_1
X_12600_ _02414_ _02538_ VGND VGND VPWR VPWR _02539_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13580_ _03536_ _03537_ _03538_ VGND VGND VPWR VPWR _03539_ sky130_fd_sc_hd__nor3_2
X_10792_ _00729_ _00730_ VGND VGND VPWR VPWR _00731_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_155_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12531_ _02461_ _02469_ VGND VGND VPWR VPWR _02470_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15250_ _05321_ _05331_ _05332_ VGND VGND VPWR VPWR _05333_ sky130_fd_sc_hd__nand3_2
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12462_ net209 _02091_ _02399_ _02400_ VGND VGND VPWR VPWR _02401_ sky130_fd_sc_hd__a31o_1
X_14201_ _04164_ _04114_ _04177_ VGND VGND VPWR VPWR _04179_ sky130_fd_sc_hd__nand3_1
X_11413_ _01314_ _01343_ _01342_ VGND VGND VPWR VPWR _01352_ sky130_fd_sc_hd__and3_1
XFILLER_0_152_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15181_ _05253_ _05235_ _05255_ VGND VGND VPWR VPWR _05257_ sky130_fd_sc_hd__nand3_1
XFILLER_0_2_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12393_ _02331_ VGND VGND VPWR VPWR _02332_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14132_ _04017_ net144 VGND VGND VPWR VPWR _04104_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11344_ _01223_ _01222_ VGND VGND VPWR VPWR _01283_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18940_ _02129_ _09289_ VGND VGND VPWR VPWR _09392_ sky130_fd_sc_hd__nor2_1
X_14063_ _04009_ _04012_ _04034_ VGND VGND VPWR VPWR _04035_ sky130_fd_sc_hd__a21oi_2
X_11275_ _01111_ _01213_ VGND VGND VPWR VPWR _01214_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_148_Right_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13014_ net264 _01797_ VGND VGND VPWR VPWR _02953_ sky130_fd_sc_hd__nand2_1
X_10226_ _00162_ _00164_ VGND VGND VPWR VPWR _00165_ sky130_fd_sc_hd__or2_1
X_18871_ _09308_ _09315_ VGND VGND VPWR VPWR _09316_ sky130_fd_sc_hd__or2_1
X_10157_ _08515_ _09065_ VGND VGND VPWR VPWR _09076_ sky130_fd_sc_hd__xor2_1
X_17822_ _08159_ _08161_ VGND VGND VPWR VPWR _08162_ sky130_fd_sc_hd__xnor2_2
X_10088_ net348 _06007_ _08306_ VGND VGND VPWR VPWR _08317_ sky130_fd_sc_hd__and3_1
X_14965_ _04972_ _05019_ VGND VGND VPWR VPWR _05020_ sky130_fd_sc_hd__nand2_1
X_17753_ net310 _07181_ VGND VGND VPWR VPWR _08087_ sky130_fd_sc_hd__nand2_2
X_13916_ _02256_ _02353_ VGND VGND VPWR VPWR _03885_ sky130_fd_sc_hd__or2_1
X_16704_ _06838_ _06932_ VGND VGND VPWR VPWR _06933_ sky130_fd_sc_hd__or2_1
X_17684_ _07996_ _08010_ VGND VGND VPWR VPWR _08011_ sky130_fd_sc_hd__nor2_1
X_14896_ _04939_ _04942_ _04943_ VGND VGND VPWR VPWR _04944_ sky130_fd_sc_hd__o21ai_2
X_16635_ _06855_ _06856_ VGND VGND VPWR VPWR _06857_ sky130_fd_sc_hd__or2_1
X_13847_ _03810_ _03812_ VGND VGND VPWR VPWR _03813_ sky130_fd_sc_hd__and2_1
X_16566_ _06778_ _06780_ VGND VGND VPWR VPWR _06781_ sky130_fd_sc_hd__nor2_1
X_13778_ _03738_ _03742_ _03743_ VGND VGND VPWR VPWR _03744_ sky130_fd_sc_hd__nand3_2
XFILLER_0_84_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15517_ _05624_ _05625_ _05626_ VGND VGND VPWR VPWR _05627_ sky130_fd_sc_hd__o21ba_1
X_18305_ _08692_ _08693_ VGND VGND VPWR VPWR _08694_ sky130_fd_sc_hd__nor2_1
X_12729_ _02573_ _02667_ VGND VGND VPWR VPWR _02668_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19285_ clknet_4_6_0_clock _00063_ VGND VGND VPWR VPWR kp\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16497_ _06399_ _06470_ _06641_ VGND VGND VPWR VPWR _06705_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_128_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18236_ net101 _01698_ _08617_ VGND VGND VPWR VPWR _08618_ sky130_fd_sc_hd__or3_1
XFILLER_0_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15448_ net471 net171 net166 net476 VGND VGND VPWR VPWR _05551_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_5_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18167_ _08540_ _08541_ i_error\[7\] VGND VGND VPWR VPWR _08542_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_4_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15379_ _05407_ _05474_ VGND VGND VPWR VPWR _05475_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17118_ _07365_ _07380_ _07387_ VGND VGND VPWR VPWR _07388_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_142_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap112 _05188_ VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__buf_1
XFILLER_0_80_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18098_ _08450_ _08461_ VGND VGND VPWR VPWR _08466_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_96_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09940_ _06656_ _06678_ VGND VGND VPWR VPWR _06689_ sky130_fd_sc_hd__nor2_1
X_17049_ _07229_ _07230_ VGND VGND VPWR VPWR _07312_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_115_Right_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09871_ _05908_ _05919_ VGND VGND VPWR VPWR _05930_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11060_ net359 _00325_ _00888_ VGND VGND VPWR VPWR _00999_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10011_ _05677_ _07448_ _07459_ VGND VGND VPWR VPWR _07470_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14750_ _04751_ _04772_ _04749_ VGND VGND VPWR VPWR _04783_ sky130_fd_sc_hd__o21ai_1
X_11962_ net200 _01875_ _01876_ VGND VGND VPWR VPWR _01901_ sky130_fd_sc_hd__a21o_1
X_13701_ _03610_ _03665_ _03608_ _03666_ VGND VGND VPWR VPWR _03667_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_99_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10913_ _00850_ _00851_ VGND VGND VPWR VPWR _00852_ sky130_fd_sc_hd__nand2_1
X_14681_ net452 net133 _04702_ _04497_ VGND VGND VPWR VPWR _04707_ sky130_fd_sc_hd__a31o_1
X_11893_ _01827_ _01831_ VGND VGND VPWR VPWR _01832_ sky130_fd_sc_hd__and2_1
X_16420_ _06619_ VGND VGND VPWR VPWR _06620_ sky130_fd_sc_hd__clkbuf_4
X_13632_ _03570_ _03590_ VGND VGND VPWR VPWR _03591_ sky130_fd_sc_hd__and2_1
X_10844_ _00779_ _00780_ _00782_ VGND VGND VPWR VPWR _00783_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_132_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16351_ net312 VGND VGND VPWR VPWR _06544_ sky130_fd_sc_hd__inv_2
X_13563_ net232 net229 _02935_ _02915_ VGND VGND VPWR VPWR _03522_ sky130_fd_sc_hd__and4_1
XFILLER_0_82_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10775_ _00706_ _00709_ VGND VGND VPWR VPWR _00714_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15302_ net464 net167 VGND VGND VPWR VPWR _05390_ sky130_fd_sc_hd__nand2_1
X_12514_ _02301_ _02303_ VGND VGND VPWR VPWR _02453_ sky130_fd_sc_hd__nand2_1
X_19070_ net505 net543 net496 VGND VGND VPWR VPWR _09519_ sky130_fd_sc_hd__o21ai_1
X_16282_ _06467_ VGND VGND VPWR VPWR _06468_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13494_ net220 _03220_ _03452_ VGND VGND VPWR VPWR _03453_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18021_ _08364_ _08374_ _08380_ VGND VGND VPWR VPWR _08381_ sky130_fd_sc_hd__or3b_1
X_15233_ _05312_ _05313_ VGND VGND VPWR VPWR _05315_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12445_ net222 _01853_ _02383_ VGND VGND VPWR VPWR _02384_ sky130_fd_sc_hd__and3_1
XFILLER_0_152_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15164_ _05225_ _05227_ _05238_ VGND VGND VPWR VPWR _05239_ sky130_fd_sc_hd__nand3_1
XFILLER_0_151_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12376_ _02228_ _02314_ VGND VGND VPWR VPWR _02315_ sky130_fd_sc_hd__or2_1
X_14115_ _04070_ _04086_ VGND VGND VPWR VPWR _04087_ sky130_fd_sc_hd__xnor2_1
X_11327_ _01226_ _01224_ VGND VGND VPWR VPWR _01266_ sky130_fd_sc_hd__xnor2_2
X_15095_ _05161_ _05147_ _05153_ VGND VGND VPWR VPWR _05163_ sky130_fd_sc_hd__nor3_1
X_18923_ _09289_ _09372_ VGND VGND VPWR VPWR _09374_ sky130_fd_sc_hd__xor2_1
X_14046_ _04017_ net156 VGND VGND VPWR VPWR _04018_ sky130_fd_sc_hd__nor2_1
X_11258_ _01081_ _01101_ _01100_ VGND VGND VPWR VPWR _01197_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10209_ _09577_ VGND VGND VPWR VPWR _09583_ sky130_fd_sc_hd__clkbuf_4
X_18854_ _09287_ _09297_ VGND VGND VPWR VPWR _09298_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11189_ _01126_ _01127_ VGND VGND VPWR VPWR _01128_ sky130_fd_sc_hd__and2b_1
X_17805_ _08137_ _08143_ VGND VGND VPWR VPWR _08144_ sky130_fd_sc_hd__xor2_1
X_18785_ _09220_ _09221_ VGND VGND VPWR VPWR _09222_ sky130_fd_sc_hd__xnor2_1
X_15997_ _01281_ _01680_ VGND VGND VPWR VPWR _06155_ sky130_fd_sc_hd__nand2_4
XFILLER_0_89_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14948_ _04954_ _04988_ _04989_ _04987_ VGND VGND VPWR VPWR _05001_ sky130_fd_sc_hd__a22o_1
X_17736_ net313 _07094_ _08066_ _08067_ VGND VGND VPWR VPWR _08068_ sky130_fd_sc_hd__nand4_1
XFILLER_0_89_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14879_ _04921_ _04924_ VGND VGND VPWR VPWR _04925_ sky130_fd_sc_hd__and2_1
X_17667_ _07984_ _07991_ VGND VGND VPWR VPWR _07992_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16618_ _06831_ _06829_ VGND VGND VPWR VPWR _06838_ sky130_fd_sc_hd__xor2_1
XFILLER_0_15_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17598_ _07912_ _07915_ VGND VGND VPWR VPWR _07916_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19337_ clknet_4_2_0_clock _00020_ VGND VGND VPWR VPWR kd_2\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16549_ net303 _06336_ _06761_ VGND VGND VPWR VPWR _06762_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19268_ clknet_4_3_0_clock _00150_ VGND VGND VPWR VPWR prev_d_error\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18219_ i_error\[11\] _08586_ VGND VGND VPWR VPWR _08599_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19199_ clknet_4_12_0_clock _00081_ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09923_ _06469_ _06491_ VGND VGND VPWR VPWR _06502_ sky130_fd_sc_hd__nor2_1
X_09854_ _05688_ _05732_ VGND VGND VPWR VPWR _05743_ sky130_fd_sc_hd__xor2_1
X_09785_ _04973_ VGND VGND VPWR VPWR _04984_ sky130_fd_sc_hd__buf_8
XFILLER_0_56_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10560_ _00498_ _00420_ VGND VGND VPWR VPWR _00499_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10491_ _00313_ _00312_ VGND VGND VPWR VPWR _00430_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12230_ _01925_ _02028_ _02027_ VGND VGND VPWR VPWR _02169_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12161_ _02075_ _02098_ VGND VGND VPWR VPWR _02100_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11112_ _01047_ _01048_ _01050_ VGND VGND VPWR VPWR _01051_ sky130_fd_sc_hd__o21bai_1
X_12092_ _02022_ _02024_ VGND VGND VPWR VPWR _02031_ sky130_fd_sc_hd__or2_1
X_15920_ _06067_ _06069_ VGND VGND VPWR VPWR _06070_ sky130_fd_sc_hd__nand2_1
X_11043_ kp\[7\] _08185_ VGND VGND VPWR VPWR _00982_ sky130_fd_sc_hd__and2_1
X_15851_ _04480_ _05993_ VGND VGND VPWR VPWR _05994_ sky130_fd_sc_hd__or2_1
X_14802_ _04837_ _04839_ VGND VGND VPWR VPWR _04840_ sky130_fd_sc_hd__and2_1
X_15782_ _05917_ _05904_ VGND VGND VPWR VPWR _05918_ sky130_fd_sc_hd__xnor2_1
X_18570_ _08979_ _08984_ VGND VGND VPWR VPWR _08985_ sky130_fd_sc_hd__nand2_1
X_12994_ _02932_ VGND VGND VPWR VPWR _02933_ sky130_fd_sc_hd__buf_4
X_14733_ _04759_ _04763_ VGND VGND VPWR VPWR _04765_ sky130_fd_sc_hd__and2_1
X_17521_ _07828_ _07830_ VGND VGND VPWR VPWR _07831_ sky130_fd_sc_hd__and2_1
X_11945_ _01883_ _01857_ VGND VGND VPWR VPWR _01884_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17452_ _07670_ _07684_ VGND VGND VPWR VPWR _07755_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14664_ net465 net129 _04482_ VGND VGND VPWR VPWR _04689_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11876_ net217 _01814_ VGND VGND VPWR VPWR _01815_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16403_ _06599_ _06600_ VGND VGND VPWR VPWR _06602_ sky130_fd_sc_hd__nor2_1
X_13615_ net261 net257 _02330_ _02407_ VGND VGND VPWR VPWR _03574_ sky130_fd_sc_hd__and4_1
XFILLER_0_95_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17383_ _07677_ _07678_ VGND VGND VPWR VPWR _07680_ sky130_fd_sc_hd__and2_1
X_10827_ net387 _00765_ _04984_ VGND VGND VPWR VPWR _00766_ sky130_fd_sc_hd__nand3_1
X_14595_ _04501_ _04498_ VGND VGND VPWR VPWR _04613_ sky130_fd_sc_hd__xnor2_1
X_19122_ net503 net556 net494 _09551_ VGND VGND VPWR VPWR _00116_ sky130_fd_sc_hd__o211a_1
X_16334_ _06508_ _06509_ _06525_ VGND VGND VPWR VPWR _06526_ sky130_fd_sc_hd__o21a_1
X_13546_ net248 _02410_ _03504_ VGND VGND VPWR VPWR _03505_ sky130_fd_sc_hd__nand3_1
X_10758_ _00624_ _00623_ VGND VGND VPWR VPWR _00697_ sky130_fd_sc_hd__nor2_1
X_19053_ _09505_ _09506_ net492 VGND VGND VPWR VPWR _00085_ sky130_fd_sc_hd__o21a_1
X_16265_ _06405_ _06449_ VGND VGND VPWR VPWR _06450_ sky130_fd_sc_hd__xnor2_1
X_13477_ _03434_ _03430_ VGND VGND VPWR VPWR _03436_ sky130_fd_sc_hd__xor2_1
XFILLER_0_113_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10689_ _00580_ _00593_ VGND VGND VPWR VPWR _00628_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15216_ _05205_ _05290_ VGND VGND VPWR VPWR _05296_ sky130_fd_sc_hd__and2_1
X_18004_ _08357_ _08355_ VGND VGND VPWR VPWR _08363_ sky130_fd_sc_hd__xnor2_1
X_12428_ net234 _01814_ VGND VGND VPWR VPWR _02367_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16196_ _06365_ _06371_ VGND VGND VPWR VPWR _06374_ sky130_fd_sc_hd__xor2_2
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15147_ _05212_ _05208_ _05210_ VGND VGND VPWR VPWR _05220_ sky130_fd_sc_hd__or3_1
X_12359_ _02294_ _02297_ _02292_ VGND VGND VPWR VPWR _02298_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15078_ _05141_ _05142_ _05143_ VGND VGND VPWR VPWR _05144_ sky130_fd_sc_hd__o21ba_1
X_14029_ _03989_ _03991_ _03996_ VGND VGND VPWR VPWR _04001_ sky130_fd_sc_hd__or3_1
X_18906_ _09224_ _09354_ VGND VGND VPWR VPWR _09355_ sky130_fd_sc_hd__xnor2_1
X_18837_ _02144_ _02142_ VGND VGND VPWR VPWR _09279_ sky130_fd_sc_hd__or2b_1
XFILLER_0_93_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18768_ _09033_ _09200_ _09202_ VGND VGND VPWR VPWR _09203_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17719_ _07969_ _07977_ _08048_ VGND VGND VPWR VPWR _08049_ sky130_fd_sc_hd__a21oi_2
X_18699_ _09075_ _09077_ _09125_ _09126_ VGND VGND VPWR VPWR _09127_ sky130_fd_sc_hd__a211o_1
XFILLER_0_93_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire2 _08904_ VGND VGND VPWR VPWR net536 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout500 net1 VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09906_ net342 _05336_ _05424_ net344 VGND VGND VPWR VPWR _06315_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09837_ net380 net376 _05061_ VGND VGND VPWR VPWR _05556_ sky130_fd_sc_hd__and3_1
X_09768_ net9 net67 VGND VGND VPWR VPWR _04797_ sky130_fd_sc_hd__or2b_1
XFILLER_0_68_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09699_ net43 _03870_ _03903_ net565 VGND VGND VPWR VPWR _00060_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11730_ _01405_ _01667_ _01456_ _01459_ VGND VGND VPWR VPWR _01669_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_139_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11661_ _01558_ _01596_ _01599_ VGND VGND VPWR VPWR _01600_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13400_ net252 _02089_ VGND VGND VPWR VPWR _03355_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10612_ _00528_ _00549_ VGND VGND VPWR VPWR _00551_ sky130_fd_sc_hd__and2_1
X_14380_ _04286_ _04374_ _04343_ _04373_ VGND VGND VPWR VPWR _04376_ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11592_ net390 _00514_ VGND VGND VPWR VPWR _01531_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13331_ _03278_ _03283_ VGND VGND VPWR VPWR _03284_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10543_ _00389_ _00391_ VGND VGND VPWR VPWR _00482_ sky130_fd_sc_hd__xor2_2
XFILLER_0_150_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16050_ _08823_ _09010_ _08988_ VGND VGND VPWR VPWR _06213_ sky130_fd_sc_hd__a21oi_1
X_13262_ _03201_ _03214_ VGND VGND VPWR VPWR _03215_ sky130_fd_sc_hd__or2_1
X_10474_ net337 _00410_ _00411_ _00412_ VGND VGND VPWR VPWR _00413_ sky130_fd_sc_hd__a31o_1
XFILLER_0_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15001_ _04979_ _05004_ _05035_ VGND VGND VPWR VPWR _05059_ sky130_fd_sc_hd__a21oi_1
X_12213_ _02150_ _02151_ VGND VGND VPWR VPWR _02152_ sky130_fd_sc_hd__xnor2_1
X_13193_ net257 _01851_ _01859_ net260 VGND VGND VPWR VPWR _03146_ sky130_fd_sc_hd__a22o_1
X_12144_ net205 _01910_ VGND VGND VPWR VPWR _02083_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16952_ _07200_ _07204_ VGND VGND VPWR VPWR _07205_ sky130_fd_sc_hd__xnor2_2
X_12075_ _01972_ _02011_ VGND VGND VPWR VPWR _02014_ sky130_fd_sc_hd__xnor2_1
X_15903_ _05102_ _05956_ VGND VGND VPWR VPWR _06052_ sky130_fd_sc_hd__nand2_1
X_11026_ net392 _05963_ _05974_ _06051_ net396 VGND VGND VPWR VPWR _00965_ sky130_fd_sc_hd__a32oi_1
X_16883_ _07125_ _07127_ _07128_ VGND VGND VPWR VPWR _07130_ sky130_fd_sc_hd__a21o_1
X_18622_ _06165_ _09041_ VGND VGND VPWR VPWR _09042_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15834_ _05968_ _05975_ VGND VGND VPWR VPWR _05976_ sky130_fd_sc_hd__xor2_1
XFILLER_0_99_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18553_ _06130_ _08965_ VGND VGND VPWR VPWR _08967_ sky130_fd_sc_hd__xnor2_1
X_15765_ _05898_ _05899_ VGND VGND VPWR VPWR _05900_ sky130_fd_sc_hd__xnor2_1
X_12977_ _01847_ _02915_ VGND VGND VPWR VPWR _02916_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17504_ _07809_ _07812_ VGND VGND VPWR VPWR _07813_ sky130_fd_sc_hd__and2_1
X_11928_ _01856_ _01866_ VGND VGND VPWR VPWR _01867_ sky130_fd_sc_hd__nor2_1
X_14716_ _04639_ _04745_ VGND VGND VPWR VPWR _04746_ sky130_fd_sc_hd__nand2_1
X_15696_ _05782_ _05823_ VGND VGND VPWR VPWR _05824_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18484_ _08886_ _08890_ VGND VGND VPWR VPWR _08891_ sky130_fd_sc_hd__or2_1
XFILLER_0_157_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14647_ _04430_ _04432_ VGND VGND VPWR VPWR _04670_ sky130_fd_sc_hd__xnor2_1
X_17435_ net273 net540 VGND VGND VPWR VPWR _07737_ sky130_fd_sc_hd__nand2_1
X_11859_ _01797_ VGND VGND VPWR VPWR _01798_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_86_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_18 net566 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14578_ _04592_ _04593_ VGND VGND VPWR VPWR _04594_ sky130_fd_sc_hd__xnor2_1
X_17366_ _07563_ _07659_ _07660_ VGND VGND VPWR VPWR _07661_ sky130_fd_sc_hd__o21a_1
XANTENNA_29 ki\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19105_ _09536_ _05336_ _09541_ net488 VGND VGND VPWR VPWR _00108_ sky130_fd_sc_hd__o211a_1
X_13529_ _03455_ _03487_ VGND VGND VPWR VPWR _03488_ sky130_fd_sc_hd__or2_1
X_16317_ _06399_ _06410_ VGND VGND VPWR VPWR _06507_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17297_ net291 _06993_ _07583_ VGND VGND VPWR VPWR _07585_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_153_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19036_ net563 net93 VGND VGND VPWR VPWR _09494_ sky130_fd_sc_hd__and2_1
X_16248_ net115 _06289_ _06430_ VGND VGND VPWR VPWR _06431_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_113_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16179_ _06347_ _06354_ VGND VGND VPWR VPWR _06355_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09622_ net42 _03091_ _03124_ net147 VGND VGND VPWR VPWR _00021_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10190_ _08383_ _09428_ VGND VGND VPWR VPWR _09439_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout330 ki\[1\] VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__clkbuf_4
Xfanout341 net342 VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__buf_2
Xfanout352 kp\[13\] VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__buf_1
XFILLER_0_17_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout363 kp\[10\] VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__clkbuf_2
Xfanout374 kp\[7\] VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__clkbuf_4
Xfanout385 net389 VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__clkbuf_4
X_12900_ _02758_ _02838_ VGND VGND VPWR VPWR _02839_ sky130_fd_sc_hd__nor2_1
Xfanout396 net398 VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__clkbuf_4
X_13880_ _03670_ _03715_ VGND VGND VPWR VPWR _03846_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12831_ _02675_ _02769_ VGND VGND VPWR VPWR _02770_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15550_ _05582_ _05658_ _05651_ _05657_ VGND VGND VPWR VPWR _05663_ sky130_fd_sc_hd__o211ai_1
X_12762_ _02599_ _02601_ VGND VGND VPWR VPWR _02701_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14501_ _04504_ _04508_ VGND VGND VPWR VPWR _04509_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11713_ _01642_ _01649_ _01651_ VGND VGND VPWR VPWR _01652_ sky130_fd_sc_hd__and3b_1
X_15481_ _05573_ _05575_ VGND VGND VPWR VPWR _05587_ sky130_fd_sc_hd__and2b_1
XFILLER_0_96_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12693_ _02630_ _02631_ VGND VGND VPWR VPWR _02632_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14432_ _04430_ _04432_ VGND VGND VPWR VPWR _04433_ sky130_fd_sc_hd__or2_1
X_17220_ net308 net305 _06721_ _06802_ VGND VGND VPWR VPWR _07500_ sky130_fd_sc_hd__and4_1
XFILLER_0_154_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11644_ _01523_ _01581_ _01582_ VGND VGND VPWR VPWR _01583_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17151_ _07386_ _07422_ VGND VGND VPWR VPWR _07424_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14363_ _04264_ _04266_ _04268_ VGND VGND VPWR VPWR _04358_ sky130_fd_sc_hd__or3_1
X_11575_ _01424_ _01470_ _01473_ VGND VGND VPWR VPWR _01514_ sky130_fd_sc_hd__o21ba_1
Xinput16 measurement[5] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
Xinput27 reg_addr[15] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16102_ prev_error\[14\] _05413_ _01811_ VGND VGND VPWR VPWR _06270_ sky130_fd_sc_hd__and3_1
Xinput38 reg_addr[8] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_1
X_13314_ _03180_ _03266_ VGND VGND VPWR VPWR _03267_ sky130_fd_sc_hd__nor2_1
X_17082_ _07245_ _07244_ VGND VGND VPWR VPWR _07348_ sky130_fd_sc_hd__and2b_1
Xinput49 reg_data[18] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10526_ _00425_ _00459_ VGND VGND VPWR VPWR _00465_ sky130_fd_sc_hd__xnor2_4
X_14294_ _04273_ _04277_ _04279_ _04281_ VGND VGND VPWR VPWR _04282_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16033_ _06178_ _06193_ VGND VGND VPWR VPWR _06195_ sky130_fd_sc_hd__xor2_1
X_13245_ _03186_ _03197_ _03195_ VGND VGND VPWR VPWR _03198_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_21_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10457_ _00378_ _00393_ _00395_ VGND VGND VPWR VPWR _00396_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_150_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13176_ _03064_ _03067_ VGND VGND VPWR VPWR _03128_ sky130_fd_sc_hd__or2b_1
X_10388_ net337 _00325_ _00326_ VGND VGND VPWR VPWR _00327_ sky130_fd_sc_hd__and3_1
X_12127_ _02060_ _02065_ VGND VGND VPWR VPWR _02066_ sky130_fd_sc_hd__nand2_1
X_17984_ _08323_ _08340_ VGND VGND VPWR VPWR _08341_ sky130_fd_sc_hd__or2_1
X_16935_ _07158_ _07180_ _07186_ VGND VGND VPWR VPWR _07187_ sky130_fd_sc_hd__o21bai_1
X_12058_ _01934_ _01995_ _01990_ VGND VGND VPWR VPWR _01997_ sky130_fd_sc_hd__or3_1
X_11009_ _00941_ _00945_ _00946_ _00947_ VGND VGND VPWR VPWR _00948_ sky130_fd_sc_hd__a211o_1
X_16866_ _07066_ _07081_ _07083_ VGND VGND VPWR VPWR _07111_ sky130_fd_sc_hd__or3_1
X_18605_ _09019_ _09023_ VGND VGND VPWR VPWR _09024_ sky130_fd_sc_hd__or2_1
X_15817_ _05102_ _05956_ VGND VGND VPWR VPWR _05957_ sky130_fd_sc_hd__or2_1
X_16797_ _07009_ _07033_ VGND VGND VPWR VPWR _07035_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18536_ _08910_ _08913_ VGND VGND VPWR VPWR _08948_ sky130_fd_sc_hd__or2b_1
X_15748_ _05848_ _05850_ VGND VGND VPWR VPWR _05881_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18467_ _08731_ _08871_ VGND VGND VPWR VPWR _08872_ sky130_fd_sc_hd__nor2_1
X_15679_ net462 net191 _05792_ _05793_ VGND VGND VPWR VPWR _05805_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_118_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17418_ _07203_ _07202_ VGND VGND VPWR VPWR _07718_ sky130_fd_sc_hd__nor2_1
X_18398_ _08560_ _08795_ VGND VGND VPWR VPWR _08796_ sky130_fd_sc_hd__or2_2
XFILLER_0_99_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17349_ _07201_ _07640_ _07641_ VGND VGND VPWR VPWR _07642_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19019_ _09451_ _09452_ _09478_ _09218_ VGND VGND VPWR VPWR _09479_ sky130_fd_sc_hd__a31o_1
XFILLER_0_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09605_ net33 net32 net79 net21 VGND VGND VPWR VPWR _03080_ sky130_fd_sc_hd__or4b_4
XFILLER_0_97_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_129_Right_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11360_ _01296_ _01298_ VGND VGND VPWR VPWR _01299_ sky130_fd_sc_hd__nor2_1
X_10311_ _00236_ _00230_ VGND VGND VPWR VPWR _00250_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_131_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11291_ net358 _00614_ _01155_ VGND VGND VPWR VPWR _01230_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_132_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13030_ _02908_ _02968_ VGND VGND VPWR VPWR _02969_ sky130_fd_sc_hd__nor2_1
X_10242_ _08471_ _08449_ VGND VGND VPWR VPWR _00181_ sky130_fd_sc_hd__xnor2_1
X_10173_ _09164_ _09219_ _09241_ VGND VGND VPWR VPWR _09252_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout160 kd_2\[8\] VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_4
X_14981_ net440 net446 net173 net168 VGND VGND VPWR VPWR _05037_ sky130_fd_sc_hd__and4_1
Xfanout171 net173 VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__buf_2
Xfanout182 kd_2\[4\] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_4
X_16720_ net303 _06346_ _06949_ VGND VGND VPWR VPWR _06950_ sky130_fd_sc_hd__and3_1
X_13932_ _03896_ _03901_ VGND VGND VPWR VPWR _03902_ sky130_fd_sc_hd__nor2_4
Xfanout193 net194 VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__buf_2
XFILLER_0_89_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16651_ _06820_ _06873_ VGND VGND VPWR VPWR _06874_ sky130_fd_sc_hd__and2_1
X_13863_ _03815_ _03825_ _03826_ _03828_ VGND VGND VPWR VPWR _03829_ sky130_fd_sc_hd__or4b_1
X_15602_ _05679_ _05711_ VGND VGND VPWR VPWR _05720_ sky130_fd_sc_hd__xor2_1
X_12814_ _02741_ _02743_ VGND VGND VPWR VPWR _02753_ sky130_fd_sc_hd__xor2_1
X_13794_ _03726_ _03759_ VGND VGND VPWR VPWR _03760_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16582_ _02328_ _06285_ _06286_ VGND VGND VPWR VPWR _06798_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_69_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18321_ _08650_ _08652_ _08648_ VGND VGND VPWR VPWR _08711_ sky130_fd_sc_hd__a21oi_1
X_15533_ _05619_ _05643_ VGND VGND VPWR VPWR _05645_ sky130_fd_sc_hd__nor2_1
X_12745_ net254 net199 _01813_ VGND VGND VPWR VPWR _02684_ sky130_fd_sc_hd__nand3_1
XFILLER_0_155_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15464_ net450 net188 VGND VGND VPWR VPWR _05569_ sky130_fd_sc_hd__nand2_1
X_18252_ net275 _06336_ _06311_ net280 VGND VGND VPWR VPWR _08635_ sky130_fd_sc_hd__a22o_1
X_12676_ _02613_ _02614_ VGND VGND VPWR VPWR _02615_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14415_ net434 net141 _04319_ _04320_ VGND VGND VPWR VPWR _04415_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_37_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17203_ _07473_ _07480_ VGND VGND VPWR VPWR _07482_ sky130_fd_sc_hd__xor2_2
X_11627_ net374 _00811_ VGND VGND VPWR VPWR _01566_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15395_ _05477_ _05480_ _05491_ VGND VGND VPWR VPWR _05493_ sky130_fd_sc_hd__or3_1
X_18183_ i_error\[0\] _08558_ VGND VGND VPWR VPWR _08560_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17134_ _07172_ _07190_ VGND VGND VPWR VPWR _07406_ sky130_fd_sc_hd__and2b_1
X_14346_ _04306_ _04317_ VGND VGND VPWR VPWR _04339_ sky130_fd_sc_hd__or2_1
X_11558_ _01494_ _01495_ _01496_ VGND VGND VPWR VPWR _01497_ sky130_fd_sc_hd__nor3_1
XFILLER_0_52_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10509_ _00437_ _00447_ _07338_ VGND VGND VPWR VPWR _00448_ sky130_fd_sc_hd__o21bai_4
X_17065_ _07289_ _07296_ _07329_ VGND VGND VPWR VPWR _07330_ sky130_fd_sc_hd__a21boi_1
X_14277_ _04257_ _04260_ _04262_ VGND VGND VPWR VPWR _04263_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_0_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11489_ _01421_ _01427_ VGND VGND VPWR VPWR _01428_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16016_ _09065_ _08515_ VGND VGND VPWR VPWR _06176_ sky130_fd_sc_hd__or2b_1
X_13228_ net237 _02331_ VGND VGND VPWR VPWR _03181_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13159_ net224 _02409_ _03028_ VGND VGND VPWR VPWR _03109_ sky130_fd_sc_hd__a21oi_1
X_17967_ _06544_ _03065_ _08321_ VGND VGND VPWR VPWR _08322_ sky130_fd_sc_hd__or3b_2
XFILLER_0_109_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16918_ net282 _06891_ _07166_ _07167_ VGND VGND VPWR VPWR _07168_ sky130_fd_sc_hd__a31o_1
X_17898_ net301 _02931_ VGND VGND VPWR VPWR _08246_ sky130_fd_sc_hd__nand2_1
X_16849_ _07090_ _07091_ VGND VGND VPWR VPWR _07092_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18519_ _08928_ VGND VGND VPWR VPWR _08929_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_3_Left_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10860_ net565 net351 _00798_ _00323_ VGND VGND VPWR VPWR _00799_ sky130_fd_sc_hd__and4_1
XFILLER_0_67_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10791_ _00639_ _00638_ VGND VGND VPWR VPWR _00730_ sky130_fd_sc_hd__or2b_1
XFILLER_0_149_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12530_ _02395_ _02459_ _02460_ VGND VGND VPWR VPWR _02469_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12461_ net219 net214 _01910_ _01875_ VGND VGND VPWR VPWR _02400_ sky130_fd_sc_hd__and4_1
XFILLER_0_152_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14200_ _04164_ _04114_ _04177_ VGND VGND VPWR VPWR _04178_ sky130_fd_sc_hd__a21o_1
XFILLER_0_124_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11412_ _01348_ _01349_ _01345_ _01347_ VGND VGND VPWR VPWR _01351_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_35_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15180_ _05253_ _05235_ _05255_ VGND VGND VPWR VPWR _05256_ sky130_fd_sc_hd__a21o_1
X_12392_ _02330_ VGND VGND VPWR VPWR _02331_ sky130_fd_sc_hd__buf_2
X_14131_ _04070_ _04086_ VGND VGND VPWR VPWR _04103_ sky130_fd_sc_hd__or2b_1
X_11343_ _01273_ _01274_ VGND VGND VPWR VPWR _01282_ sky130_fd_sc_hd__xor2_4
X_14062_ _04032_ _04033_ VGND VGND VPWR VPWR _04034_ sky130_fd_sc_hd__nand2_1
X_11274_ _01110_ _00911_ VGND VGND VPWR VPWR _01213_ sky130_fd_sc_hd__and2b_1
X_13013_ net264 _01812_ _02951_ VGND VGND VPWR VPWR _02952_ sky130_fd_sc_hd__and3_1
X_10225_ _07778_ _00163_ _07349_ VGND VGND VPWR VPWR _00164_ sky130_fd_sc_hd__o21a_1
X_18870_ _01929_ _09314_ VGND VGND VPWR VPWR _09315_ sky130_fd_sc_hd__xnor2_1
X_17821_ _08160_ _08040_ VGND VGND VPWR VPWR _08161_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_100_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10156_ _09043_ _09054_ VGND VGND VPWR VPWR _09065_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17752_ net307 _07156_ VGND VGND VPWR VPWR _08085_ sky130_fd_sc_hd__nand2_1
X_14964_ _04969_ _04971_ VGND VGND VPWR VPWR _05019_ sky130_fd_sc_hd__or2_1
X_10087_ _08284_ _08295_ VGND VGND VPWR VPWR _08306_ sky130_fd_sc_hd__nor2_1
X_16703_ _06839_ _06926_ _06930_ VGND VGND VPWR VPWR _06932_ sky130_fd_sc_hd__o21a_1
X_13915_ _02466_ _03883_ VGND VGND VPWR VPWR _03884_ sky130_fd_sc_hd__nor2_1
X_17683_ _08007_ _08008_ VGND VGND VPWR VPWR _08010_ sky130_fd_sc_hd__nand2_1
X_14895_ _04934_ _04937_ VGND VGND VPWR VPWR _04943_ sky130_fd_sc_hd__xor2_1
X_16634_ _06844_ _06851_ _06853_ VGND VGND VPWR VPWR _06856_ sky130_fd_sc_hd__and3_1
X_13846_ net261 _02935_ _03811_ VGND VGND VPWR VPWR _03812_ sky130_fd_sc_hd__and3_1
X_16565_ _06779_ _06714_ VGND VGND VPWR VPWR _06780_ sky130_fd_sc_hd__xor2_1
XFILLER_0_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13777_ _03721_ _03737_ VGND VGND VPWR VPWR _03743_ sky130_fd_sc_hd__nand2_1
X_10989_ _00927_ _00834_ VGND VGND VPWR VPWR _00928_ sky130_fd_sc_hd__xor2_4
XFILLER_0_73_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18304_ _06399_ _06386_ _06336_ net273 VGND VGND VPWR VPWR _08693_ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15516_ net452 net457 net188 net183 VGND VGND VPWR VPWR _05626_ sky130_fd_sc_hd__and4_1
XFILLER_0_45_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12728_ _02575_ _02628_ _02666_ VGND VGND VPWR VPWR _02667_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19284_ clknet_4_7_0_clock _00062_ VGND VGND VPWR VPWR kp\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16496_ _06695_ _06684_ VGND VGND VPWR VPWR _06704_ sky130_fd_sc_hd__or2b_1
XFILLER_0_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18235_ _06131_ _06133_ _08616_ VGND VGND VPWR VPWR _08617_ sky130_fd_sc_hd__nand3_2
X_12659_ net243 _01834_ VGND VGND VPWR VPWR _02598_ sky130_fd_sc_hd__nand2_2
X_15447_ net471 net476 net171 net166 VGND VGND VPWR VPWR _05550_ sky130_fd_sc_hd__and4_1
XFILLER_0_155_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18166_ _08478_ _08538_ _08539_ VGND VGND VPWR VPWR _08541_ sky130_fd_sc_hd__and3b_1
X_15378_ net482 net153 _05405_ _05406_ VGND VGND VPWR VPWR _05474_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_53_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17117_ _07364_ _07353_ VGND VGND VPWR VPWR _07387_ sky130_fd_sc_hd__or2b_1
Xmax_cap102 _08164_ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__buf_1
X_14329_ net438 net137 net136 net443 VGND VGND VPWR VPWR _04320_ sky130_fd_sc_hd__a22oi_1
Xmax_cap113 _04045_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__buf_1
X_18097_ _08463_ _08464_ VGND VGND VPWR VPWR _08465_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_123_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17048_ _07309_ _07297_ VGND VGND VPWR VPWR _07311_ sky130_fd_sc_hd__xor2_2
X_09870_ _04566_ _04577_ _05897_ VGND VGND VPWR VPWR _05919_ sky130_fd_sc_hd__nand3_2
XFILLER_0_110_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18999_ _09195_ _09070_ VGND VGND VPWR VPWR _09457_ sky130_fd_sc_hd__and2b_1
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10010_ net356 _05600_ _05006_ kp\[13\] VGND VGND VPWR VPWR _07459_ sky130_fd_sc_hd__a22oi_1
X_09999_ net402 _07327_ VGND VGND VPWR VPWR _07338_ sky130_fd_sc_hd__and2_2
XPHY_EDGE_ROW_48_Left_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11961_ net208 _01861_ _01899_ VGND VGND VPWR VPWR _01900_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13700_ _03556_ _03607_ VGND VGND VPWR VPWR _03666_ sky130_fd_sc_hd__or2_1
X_10912_ _00847_ _00845_ VGND VGND VPWR VPWR _00851_ sky130_fd_sc_hd__xnor2_2
X_14680_ net464 net133 _04691_ VGND VGND VPWR VPWR _04706_ sky130_fd_sc_hd__and3_1
X_11892_ net221 _01817_ _01830_ _01828_ VGND VGND VPWR VPWR _01831_ sky130_fd_sc_hd__a31o_1
X_13631_ _03565_ _03569_ VGND VGND VPWR VPWR _03590_ sky130_fd_sc_hd__nand2_1
X_10843_ net363 _08196_ _00781_ VGND VGND VPWR VPWR _00782_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13562_ _03519_ _03520_ VGND VGND VPWR VPWR _03521_ sky130_fd_sc_hd__xnor2_1
X_16350_ net312 _01755_ _06316_ VGND VGND VPWR VPWR _06543_ sky130_fd_sc_hd__and3_1
X_10774_ net340 _00615_ _00711_ _00712_ VGND VGND VPWR VPWR _00713_ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12513_ _02449_ _02451_ VGND VGND VPWR VPWR _02452_ sky130_fd_sc_hd__nand2_1
X_15301_ net468 net162 net145 net486 VGND VGND VPWR VPWR _05389_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_94_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16281_ _06466_ VGND VGND VPWR VPWR _06467_ sky130_fd_sc_hd__buf_2
X_13493_ _03447_ _03451_ VGND VGND VPWR VPWR _03452_ sky130_fd_sc_hd__xor2_1
XFILLER_0_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_57_Left_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18020_ _08376_ _08377_ _08379_ VGND VGND VPWR VPWR _08380_ sky130_fd_sc_hd__a21bo_1
X_12444_ _02285_ _02380_ _02382_ VGND VGND VPWR VPWR _02383_ sky130_fd_sc_hd__o21a_1
X_15232_ net464 net162 VGND VGND VPWR VPWR _05313_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15163_ _05235_ _05236_ VGND VGND VPWR VPWR _05238_ sky130_fd_sc_hd__and2_1
X_12375_ net201 _02224_ _02227_ VGND VGND VPWR VPWR _02314_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14114_ _04084_ _04085_ VGND VGND VPWR VPWR _04086_ sky130_fd_sc_hd__and2_1
X_11326_ _01250_ _01251_ _01264_ VGND VGND VPWR VPWR _01265_ sky130_fd_sc_hd__nand3_4
X_15094_ _05147_ _05153_ _05161_ VGND VGND VPWR VPWR _05162_ sky130_fd_sc_hd__o21a_1
X_14045_ _04016_ VGND VGND VPWR VPWR _04017_ sky130_fd_sc_hd__clkbuf_4
X_18922_ _09311_ _09312_ _02148_ VGND VGND VPWR VPWR _09372_ sky130_fd_sc_hd__o21bai_1
X_11257_ _01081_ _01100_ _01101_ VGND VGND VPWR VPWR _01196_ sky130_fd_sc_hd__and3_1
X_10208_ _09571_ VGND VGND VPWR VPWR _09577_ sky130_fd_sc_hd__clkbuf_4
X_18853_ _09294_ _09295_ VGND VGND VPWR VPWR _09297_ sky130_fd_sc_hd__nor2_1
X_11188_ _01124_ _01123_ VGND VGND VPWR VPWR _01127_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_66_Left_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17804_ _08126_ _08142_ VGND VGND VPWR VPWR _08143_ sky130_fd_sc_hd__xnor2_1
X_10139_ _07448_ _08867_ _05600_ VGND VGND VPWR VPWR _08878_ sky130_fd_sc_hd__and3b_1
X_18784_ _09024_ _09031_ _09216_ VGND VGND VPWR VPWR _09221_ sky130_fd_sc_hd__o21ba_1
X_15996_ _06145_ _06153_ VGND VGND VPWR VPWR _06154_ sky130_fd_sc_hd__and2b_1
X_17735_ net331 net314 _06618_ _06992_ VGND VGND VPWR VPWR _08067_ sky130_fd_sc_hd__nand4_2
X_14947_ _04998_ _04999_ VGND VGND VPWR VPWR _05000_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17666_ _07984_ _07985_ _07990_ VGND VGND VPWR VPWR _07991_ sky130_fd_sc_hd__nand3_1
X_14878_ _04862_ _04923_ VGND VGND VPWR VPWR _04924_ sky130_fd_sc_hd__nor2_1
X_16617_ _06752_ _06834_ VGND VGND VPWR VPWR _06837_ sky130_fd_sc_hd__xnor2_1
X_13829_ _03762_ _03792_ _03794_ VGND VGND VPWR VPWR _03795_ sky130_fd_sc_hd__o21ai_2
X_17597_ _07913_ _07914_ VGND VGND VPWR VPWR _07915_ sky130_fd_sc_hd__xor2_1
XFILLER_0_58_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19336_ clknet_4_2_0_clock _00037_ VGND VGND VPWR VPWR kd_2\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16548_ _06759_ _06760_ VGND VGND VPWR VPWR _06761_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_75_Left_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19267_ clknet_4_12_0_clock _00149_ VGND VGND VPWR VPWR prev_d_error\[16\] sky130_fd_sc_hd__dfxtp_1
X_16479_ net293 _06353_ VGND VGND VPWR VPWR _06685_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18218_ i_error\[11\] _08586_ _08589_ i_error\[10\] VGND VGND VPWR VPWR _08598_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_32_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19198_ clknet_4_14_0_clock _00080_ VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18149_ _06934_ _07046_ _08520_ _08521_ VGND VGND VPWR VPWR _08522_ sky130_fd_sc_hd__a31o_1
XFILLER_0_13_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09922_ _05380_ _06480_ VGND VGND VPWR VPWR _06491_ sky130_fd_sc_hd__xor2_1
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_84_Left_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09853_ _05710_ _05721_ VGND VGND VPWR VPWR _05732_ sky130_fd_sc_hd__xor2_2
X_09784_ _04918_ _04962_ VGND VGND VPWR VPWR _04973_ sky130_fd_sc_hd__xor2_4
XFILLER_0_95_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_93_Left_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10490_ _00424_ _00428_ VGND VGND VPWR VPWR _00429_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12160_ _01848_ _01910_ VGND VGND VPWR VPWR _02099_ sky130_fd_sc_hd__or2_1
X_11111_ net392 _05963_ _05974_ _01049_ VGND VGND VPWR VPWR _01050_ sky130_fd_sc_hd__and4_1
X_12091_ _01925_ _02029_ VGND VGND VPWR VPWR _02030_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11042_ _00977_ _00980_ VGND VGND VPWR VPWR _00981_ sky130_fd_sc_hd__xnor2_2
X_15850_ _05981_ _05982_ _05992_ VGND VGND VPWR VPWR _05993_ sky130_fd_sc_hd__o21a_1
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14801_ _04756_ _04838_ VGND VGND VPWR VPWR _04839_ sky130_fd_sc_hd__nor2_1
X_15781_ _05879_ _05894_ VGND VGND VPWR VPWR _05917_ sky130_fd_sc_hd__or2_1
X_12993_ _02931_ VGND VGND VPWR VPWR _02932_ sky130_fd_sc_hd__buf_2
X_17520_ _07662_ _07829_ VGND VGND VPWR VPWR _07830_ sky130_fd_sc_hd__nor2_1
X_14732_ _04754_ _04756_ _04758_ VGND VGND VPWR VPWR _04763_ sky130_fd_sc_hd__or3_1
X_11944_ net203 _01808_ VGND VGND VPWR VPWR _01883_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17451_ _07736_ _07753_ VGND VGND VPWR VPWR _07754_ sky130_fd_sc_hd__xnor2_1
X_14663_ _04617_ _04682_ _04686_ VGND VGND VPWR VPWR _04688_ sky130_fd_sc_hd__or3_1
X_11875_ _01813_ VGND VGND VPWR VPWR _01814_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_86_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16402_ net296 _06335_ _06311_ net300 VGND VGND VPWR VPWR _06600_ sky130_fd_sc_hd__a22oi_1
X_13614_ _03564_ _03570_ _03572_ VGND VGND VPWR VPWR _03573_ sky130_fd_sc_hd__a21oi_1
X_10826_ net405 _05292_ _05303_ VGND VGND VPWR VPWR _00765_ sky130_fd_sc_hd__and3_1
X_17382_ net280 _07183_ net540 net274 VGND VGND VPWR VPWR _07678_ sky130_fd_sc_hd__a22o_1
X_14594_ _04609_ _04611_ VGND VGND VPWR VPWR _04612_ sky130_fd_sc_hd__or2_1
X_19121_ _09099_ _09100_ _09550_ VGND VGND VPWR VPWR _09551_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16333_ _06522_ _06523_ VGND VGND VPWR VPWR _06525_ sky130_fd_sc_hd__and2_1
X_13545_ _03502_ _03503_ VGND VGND VPWR VPWR _03504_ sky130_fd_sc_hd__xor2_1
X_10757_ _00682_ _00695_ VGND VGND VPWR VPWR _00696_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19052_ _09447_ _09485_ _09458_ VGND VGND VPWR VPWR _09506_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13476_ _03430_ _03434_ VGND VGND VPWR VPWR _03435_ sky130_fd_sc_hd__and2b_1
X_16264_ _06446_ _06448_ VGND VGND VPWR VPWR _06449_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10688_ _00529_ _00547_ VGND VGND VPWR VPWR _00627_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18003_ _08359_ _08360_ VGND VGND VPWR VPWR _08362_ sky130_fd_sc_hd__nor2_1
X_12427_ _02362_ _02363_ _02365_ VGND VGND VPWR VPWR _02366_ sky130_fd_sc_hd__o21ba_1
X_15215_ _05293_ _05294_ VGND VGND VPWR VPWR _05295_ sky130_fd_sc_hd__nand2_1
X_16195_ _06366_ _06368_ VGND VGND VPWR VPWR _06373_ sky130_fd_sc_hd__or2_1
X_12358_ _02295_ _02296_ VGND VGND VPWR VPWR _02297_ sky130_fd_sc_hd__xnor2_1
X_15146_ _05217_ _05218_ VGND VGND VPWR VPWR _05219_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11309_ _01247_ _01241_ VGND VGND VPWR VPWR _01248_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15077_ net441 net446 net177 net172 VGND VGND VPWR VPWR _05143_ sky130_fd_sc_hd__and4_1
X_12289_ net201 _02224_ _02227_ VGND VGND VPWR VPWR _02228_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14028_ _03998_ _03999_ net407 net160 VGND VGND VPWR VPWR _04000_ sky130_fd_sc_hd__and4bb_1
X_18905_ _09352_ _09353_ VGND VGND VPWR VPWR _09354_ sky130_fd_sc_hd__or2b_1
X_18836_ _09275_ _09277_ VGND VGND VPWR VPWR _09278_ sky130_fd_sc_hd__xor2_1
XFILLER_0_93_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18767_ _09024_ _09031_ _09201_ VGND VGND VPWR VPWR _09202_ sky130_fd_sc_hd__o21ai_1
X_15979_ _00759_ net533 VGND VGND VPWR VPWR _06135_ sky130_fd_sc_hd__xor2_4
XFILLER_0_89_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17718_ _08044_ _08046_ _08047_ _07966_ VGND VGND VPWR VPWR _08048_ sky130_fd_sc_hd__o211a_4
XFILLER_0_117_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18698_ _06146_ _08620_ _08881_ VGND VGND VPWR VPWR _09126_ sky130_fd_sc_hd__and3_1
XFILLER_0_148_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17649_ _07969_ _07970_ _07971_ VGND VGND VPWR VPWR _07972_ sky130_fd_sc_hd__and3b_1
XFILLER_0_58_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19319_ clknet_4_1_0_clock _00002_ VGND VGND VPWR VPWR kd_1\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout501 net502 VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__clkbuf_2
X_09905_ net344 net341 _05325_ _05424_ VGND VGND VPWR VPWR _06304_ sky130_fd_sc_hd__and4_1
XFILLER_0_10_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09836_ net384 _05072_ _05490_ _05534_ VGND VGND VPWR VPWR _05545_ sky130_fd_sc_hd__a31o_2
X_09767_ _04170_ _04764_ _04775_ VGND VGND VPWR VPWR _04786_ sky130_fd_sc_hd__a21o_4
X_09698_ net42 _03870_ _03903_ net358 VGND VGND VPWR VPWR _00059_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11660_ net399 _00515_ _01597_ _01598_ VGND VGND VPWR VPWR _01599_ sky130_fd_sc_hd__a31o_1
XFILLER_0_83_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10611_ _00528_ _00549_ VGND VGND VPWR VPWR _00550_ sky130_fd_sc_hd__nor2_1
X_11591_ net400 _00243_ _01528_ _01487_ VGND VGND VPWR VPWR _01530_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13330_ _03276_ _03277_ VGND VGND VPWR VPWR _03283_ sky130_fd_sc_hd__or2_1
X_10542_ _00474_ _00479_ _00480_ VGND VGND VPWR VPWR _00481_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_36_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13261_ _03203_ _03212_ _03213_ VGND VGND VPWR VPWR _03214_ sky130_fd_sc_hd__o21a_1
X_10473_ net343 _00324_ _00320_ VGND VGND VPWR VPWR _00412_ sky130_fd_sc_hd__and3_1
X_12212_ net210 _01787_ VGND VGND VPWR VPWR _02151_ sky130_fd_sc_hd__nand2_1
X_15000_ _05055_ _05056_ _05044_ _05049_ VGND VGND VPWR VPWR _05058_ sky130_fd_sc_hd__a211o_1
XFILLER_0_32_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13192_ _03143_ _03144_ VGND VGND VPWR VPWR _03145_ sky130_fd_sc_hd__xor2_1
XFILLER_0_60_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12143_ _01914_ _02081_ VGND VGND VPWR VPWR _02082_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12074_ _02011_ _02012_ VGND VGND VPWR VPWR _02013_ sky130_fd_sc_hd__and2_1
X_16951_ _07201_ _07202_ _07203_ VGND VGND VPWR VPWR _07204_ sky130_fd_sc_hd__o21ba_2
X_15902_ _06048_ _06049_ VGND VGND VPWR VPWR _06050_ sky130_fd_sc_hd__nand2_1
X_11025_ net402 VGND VGND VPWR VPWR _00964_ sky130_fd_sc_hd__inv_2
X_16882_ _07124_ _07123_ VGND VGND VPWR VPWR _07128_ sky130_fd_sc_hd__and2b_1
X_18621_ _09036_ _09039_ VGND VGND VPWR VPWR _09041_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15833_ _05972_ _05973_ VGND VGND VPWR VPWR _05975_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18552_ _06268_ _08884_ _08964_ VGND VGND VPWR VPWR _08965_ sky130_fd_sc_hd__mux2_2
X_15764_ _05872_ _05871_ VGND VGND VPWR VPWR _05899_ sky130_fd_sc_hd__and2b_1
XFILLER_0_59_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12976_ _02914_ VGND VGND VPWR VPWR _02915_ sky130_fd_sc_hd__clkbuf_4
X_17503_ net310 _06801_ _06890_ net307 VGND VGND VPWR VPWR _07812_ sky130_fd_sc_hd__a22o_1
X_14715_ _04636_ _04638_ VGND VGND VPWR VPWR _04745_ sky130_fd_sc_hd__or2_1
XFILLER_0_157_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11927_ _01864_ _01865_ VGND VGND VPWR VPWR _01866_ sky130_fd_sc_hd__or2_1
X_18483_ _08887_ _06266_ _08888_ VGND VGND VPWR VPWR _08890_ sky130_fd_sc_hd__or3_1
X_15695_ _05774_ _05781_ VGND VGND VPWR VPWR _05823_ sky130_fd_sc_hd__and2_1
XFILLER_0_144_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17434_ _07636_ _07651_ _07735_ VGND VGND VPWR VPWR _07736_ sky130_fd_sc_hd__a21o_1
X_14646_ _04667_ _04668_ VGND VGND VPWR VPWR _04669_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11858_ _01796_ _01750_ VGND VGND VPWR VPWR _01797_ sky130_fd_sc_hd__xor2_4
XFILLER_0_83_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17365_ net290 _07182_ _07568_ net287 VGND VGND VPWR VPWR _07660_ sky130_fd_sc_hd__a22o_1
XANTENNA_19 net345 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10809_ _00721_ _00746_ VGND VGND VPWR VPWR _00748_ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14577_ _04487_ _04491_ _04488_ VGND VGND VPWR VPWR _04593_ sky130_fd_sc_hd__o21ba_1
X_11789_ _01723_ _01725_ _01726_ _01727_ VGND VGND VPWR VPWR _01728_ sky130_fd_sc_hd__a211o_1
X_19104_ net499 prev_error\[13\] VGND VGND VPWR VPWR _09541_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16316_ _06488_ _06504_ _06505_ VGND VGND VPWR VPWR _06506_ sky130_fd_sc_hd__a21o_1
X_13528_ _03445_ _03454_ VGND VGND VPWR VPWR _03487_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17296_ net291 _06993_ _07583_ VGND VGND VPWR VPWR _07584_ sky130_fd_sc_hd__and3_1
XFILLER_0_141_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19035_ _09492_ _09493_ net492 VGND VGND VPWR VPWR _00079_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16247_ _01849_ _06290_ _06288_ _06294_ VGND VGND VPWR VPWR _06430_ sky130_fd_sc_hd__a22o_1
X_13459_ _03344_ _03416_ VGND VGND VPWR VPWR _03418_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16178_ net286 _06353_ VGND VGND VPWR VPWR _06354_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15129_ _05198_ _05199_ VGND VGND VPWR VPWR _05200_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09621_ net41 _03091_ _03124_ net152 VGND VGND VPWR VPWR _00020_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18819_ _03921_ _09258_ VGND VGND VPWR VPWR _09259_ sky130_fd_sc_hd__xor2_1
XFILLER_0_78_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout320 net321 VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__clkbuf_4
Xfanout331 net334 VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__clkbuf_4
Xfanout342 kp\[16\] VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__clkbuf_4
Xfanout353 net354 VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__buf_2
Xfanout364 net365 VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__clkbuf_4
Xfanout375 net376 VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__clkbuf_4
Xfanout386 net389 VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__dlymetal6s2s_1
X_09819_ net5 _04731_ net63 VGND VGND VPWR VPWR _05358_ sky130_fd_sc_hd__or3b_1
Xfanout397 net398 VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_21_Left_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12830_ _02676_ _02768_ VGND VGND VPWR VPWR _02769_ sky130_fd_sc_hd__nor2_1
X_12761_ net246 _01807_ _02689_ _02699_ VGND VGND VPWR VPWR _02700_ sky130_fd_sc_hd__a31o_1
XFILLER_0_33_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14500_ _04505_ _04507_ VGND VGND VPWR VPWR _04508_ sky130_fd_sc_hd__nor2_1
X_11712_ _01639_ _01650_ _01550_ VGND VGND VPWR VPWR _01651_ sky130_fd_sc_hd__and3b_1
X_12692_ _02555_ _02557_ VGND VGND VPWR VPWR _02631_ sky130_fd_sc_hd__xor2_1
X_15480_ _05568_ _05583_ _05585_ VGND VGND VPWR VPWR _05586_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14431_ _04409_ _04431_ VGND VGND VPWR VPWR _04432_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11643_ _01540_ _01544_ _01525_ VGND VGND VPWR VPWR _01582_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17150_ _07386_ _07422_ VGND VGND VPWR VPWR _07423_ sky130_fd_sc_hd__xor2_2
X_14362_ _04351_ _04353_ _04355_ VGND VGND VPWR VPWR _04356_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_64_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11574_ net385 _01286_ _00516_ _01512_ VGND VGND VPWR VPWR _01513_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_30_Left_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput17 measurement[6] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
Xinput28 reg_addr[16] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16101_ prev_error\[16\] _04841_ _04852_ VGND VGND VPWR VPWR _06269_ sky130_fd_sc_hd__and3_1
Xinput39 reg_addr[9] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
X_13313_ _03230_ _03265_ _03263_ VGND VGND VPWR VPWR _03266_ sky130_fd_sc_hd__o21a_1
X_10525_ _00462_ _00463_ VGND VGND VPWR VPWR _00464_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_134_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14293_ _04245_ _04248_ _04278_ VGND VGND VPWR VPWR _04281_ sky130_fd_sc_hd__nand3_1
XFILLER_0_52_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17081_ _07345_ _07344_ _07314_ _07310_ VGND VGND VPWR VPWR _07347_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_80_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16032_ _06191_ _06192_ VGND VGND VPWR VPWR _06193_ sky130_fd_sc_hd__nor2_1
X_13244_ _03195_ _03196_ VGND VGND VPWR VPWR _03197_ sky130_fd_sc_hd__nor2_1
X_10456_ _00342_ _00394_ VGND VGND VPWR VPWR _00395_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13175_ _03123_ _03126_ VGND VGND VPWR VPWR _03127_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10387_ _00247_ _00320_ VGND VGND VPWR VPWR _00326_ sky130_fd_sc_hd__xor2_1
X_12126_ _02062_ _02064_ VGND VGND VPWR VPWR _02065_ sky130_fd_sc_hd__or2b_1
X_17983_ _08249_ _08319_ _08322_ VGND VGND VPWR VPWR _08340_ sky130_fd_sc_hd__and3_1
X_16934_ net271 _07183_ _07185_ VGND VGND VPWR VPWR _07186_ sky130_fd_sc_hd__and3_1
X_12057_ _01934_ _01990_ _01995_ VGND VGND VPWR VPWR _01996_ sky130_fd_sc_hd__o21ai_1
X_11008_ _00854_ _00853_ _00830_ VGND VGND VPWR VPWR _00947_ sky130_fd_sc_hd__a21oi_1
X_16865_ _07086_ _07109_ _07106_ VGND VGND VPWR VPWR _07110_ sky130_fd_sc_hd__a21oi_2
X_18604_ _06168_ _09018_ VGND VGND VPWR VPWR _09023_ sky130_fd_sc_hd__nor2_1
X_15816_ _05200_ _05955_ _05198_ VGND VGND VPWR VPWR _05956_ sky130_fd_sc_hd__o21a_1
X_16796_ _07009_ _07033_ VGND VGND VPWR VPWR _07034_ sky130_fd_sc_hd__xor2_1
X_18535_ _08923_ _08945_ _08946_ _08920_ VGND VGND VPWR VPWR _08947_ sky130_fd_sc_hd__a2bb2o_1
X_15747_ _05870_ _05873_ _05879_ VGND VGND VPWR VPWR _05880_ sky130_fd_sc_hd__a21oi_1
X_12959_ _02613_ _02311_ _02818_ _02897_ VGND VGND VPWR VPWR _02898_ sky130_fd_sc_hd__o31a_1
X_18466_ _01698_ _08617_ _06261_ net101 VGND VGND VPWR VPWR _08871_ sky130_fd_sc_hd__o211a_1
X_15678_ _05801_ _05803_ VGND VGND VPWR VPWR _05804_ sky130_fd_sc_hd__nor2_2
XFILLER_0_157_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17417_ _07618_ _07628_ _07716_ VGND VGND VPWR VPWR _07717_ sky130_fd_sc_hd__a21o_1
X_14629_ _04398_ _04407_ VGND VGND VPWR VPWR _04650_ sky130_fd_sc_hd__xnor2_1
X_18397_ i_error\[0\] _08558_ VGND VGND VPWR VPWR _08795_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17348_ net299 _06723_ _07581_ VGND VGND VPWR VPWR _07641_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_16_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17279_ _07563_ _07564_ VGND VGND VPWR VPWR _07565_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19018_ _09456_ _09458_ _09459_ _09477_ VGND VGND VPWR VPWR _09478_ sky130_fd_sc_hd__and4_1
XFILLER_0_140_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09604_ _03058_ VGND VGND VPWR VPWR _03069_ sky130_fd_sc_hd__buf_2
XFILLER_0_3_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10310_ net339 _00245_ _00246_ _00248_ VGND VGND VPWR VPWR _00249_ sky130_fd_sc_hd__a31o_1
XFILLER_0_104_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11290_ _01220_ _01227_ _01228_ VGND VGND VPWR VPWR _01229_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10241_ _00178_ _00179_ VGND VGND VPWR VPWR _00180_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10172_ _07954_ _09230_ VGND VGND VPWR VPWR _09241_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14980_ _04979_ _05004_ _05035_ VGND VGND VPWR VPWR _05036_ sky130_fd_sc_hd__and3_1
Xfanout150 kd_2\[11\] VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_2
Xfanout161 kd_2\[8\] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_2
Xfanout172 net173 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__buf_2
Xfanout183 net185 VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__buf_2
X_13931_ _03899_ _03900_ VGND VGND VPWR VPWR _03901_ sky130_fd_sc_hd__xor2_2
Xfanout194 kd_2\[1\] VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__buf_4
X_16650_ _06398_ _06724_ _06819_ VGND VGND VPWR VPWR _06873_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13862_ net267 _02747_ _03827_ VGND VGND VPWR VPWR _03828_ sky130_fd_sc_hd__and3_1
X_15601_ _05717_ _05718_ VGND VGND VPWR VPWR _05719_ sky130_fd_sc_hd__nor2_1
X_12813_ net202 _02747_ _02749_ _02751_ VGND VGND VPWR VPWR _02752_ sky130_fd_sc_hd__a31o_1
X_16581_ _06729_ _06796_ VGND VGND VPWR VPWR _06797_ sky130_fd_sc_hd__nand2_1
X_13793_ net263 _02543_ _03725_ VGND VGND VPWR VPWR _03759_ sky130_fd_sc_hd__a21oi_1
X_18320_ i_error\[18\] _08709_ VGND VGND VPWR VPWR _08710_ sky130_fd_sc_hd__xnor2_1
X_15532_ net462 net179 _05642_ _05617_ VGND VGND VPWR VPWR _05643_ sky130_fd_sc_hd__o2bb2a_1
X_12744_ _02577_ _02682_ VGND VGND VPWR VPWR _02683_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18251_ net277 _06311_ VGND VGND VPWR VPWR _08634_ sky130_fd_sc_hd__nand2_1
X_15463_ _05555_ _05564_ _05566_ VGND VGND VPWR VPWR _05568_ sky130_fd_sc_hd__a21o_1
X_12675_ _01873_ VGND VGND VPWR VPWR _02614_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17202_ net319 _06463_ _06465_ VGND VGND VPWR VPWR _07480_ sky130_fd_sc_hd__and3_2
X_14414_ _04410_ _04413_ VGND VGND VPWR VPWR _04414_ sky130_fd_sc_hd__nor2_1
X_11626_ _01551_ _01552_ _01564_ VGND VGND VPWR VPWR _01565_ sky130_fd_sc_hd__o21ai_1
X_18182_ _08430_ _08557_ VGND VGND VPWR VPWR _08558_ sky130_fd_sc_hd__nor2_1
X_15394_ _05477_ _05480_ _05491_ VGND VGND VPWR VPWR _05492_ sky130_fd_sc_hd__o21ai_2
X_17133_ _07388_ _07403_ VGND VGND VPWR VPWR _07405_ sky130_fd_sc_hd__xor2_2
XFILLER_0_142_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14345_ _04334_ _04336_ _04326_ _04330_ VGND VGND VPWR VPWR _04338_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_4_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11557_ _01440_ _01482_ _01493_ VGND VGND VPWR VPWR _01496_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10508_ _00442_ _00443_ _00446_ _07338_ VGND VGND VPWR VPWR _00447_ sky130_fd_sc_hd__a31o_2
XFILLER_0_111_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17064_ _07284_ _07288_ VGND VGND VPWR VPWR _07329_ sky130_fd_sc_hd__nand2_1
X_14276_ _04000_ _04261_ VGND VGND VPWR VPWR _04262_ sky130_fd_sc_hd__nor2_1
X_11488_ _01365_ _01422_ _01423_ _01426_ VGND VGND VPWR VPWR _01427_ sky130_fd_sc_hd__o22a_1
X_16015_ _06174_ _01698_ VGND VGND VPWR VPWR _06175_ sky130_fd_sc_hd__and2_1
XFILLER_0_150_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13227_ _03139_ _03175_ VGND VGND VPWR VPWR _03180_ sky130_fd_sc_hd__xnor2_1
X_10439_ _00375_ _00377_ VGND VGND VPWR VPWR _00378_ sky130_fd_sc_hd__nand2_1
X_13158_ _03099_ _03105_ _03107_ VGND VGND VPWR VPWR _03108_ sky130_fd_sc_hd__a21oi_1
X_12109_ _01833_ _01842_ VGND VGND VPWR VPWR _02048_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13089_ net211 _02641_ _02921_ VGND VGND VPWR VPWR _03032_ sky130_fd_sc_hd__a21oi_1
X_17966_ _08319_ _08320_ VGND VGND VPWR VPWR _08321_ sky130_fd_sc_hd__and2_1
X_16917_ net288 net285 _06723_ _06803_ VGND VGND VPWR VPWR _07167_ sky130_fd_sc_hd__and4_1
X_17897_ _08237_ _08238_ _08235_ VGND VGND VPWR VPWR _08245_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16848_ _06994_ _06996_ VGND VGND VPWR VPWR _07091_ sky130_fd_sc_hd__xnor2_1
X_16779_ net324 net320 _06323_ _06540_ VGND VGND VPWR VPWR _07015_ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18518_ _06265_ _08794_ VGND VGND VPWR VPWR _08928_ sky130_fd_sc_hd__or2b_1
XFILLER_0_87_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18449_ _06163_ _06165_ VGND VGND VPWR VPWR _08852_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_141_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclone2 _04181_ net510 _04720_ _04731_ _04753_ VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__a311o_1
XFILLER_0_79_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10790_ net397 _04874_ VGND VGND VPWR VPWR _00729_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12460_ net214 _01910_ _01875_ net219 VGND VGND VPWR VPWR _02399_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11411_ _01345_ _01347_ _01348_ _01349_ VGND VGND VPWR VPWR _01350_ sky130_fd_sc_hd__a211o_2
XFILLER_0_105_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12391_ _02329_ VGND VGND VPWR VPWR _02330_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14130_ _04095_ VGND VGND VPWR VPWR _04102_ sky130_fd_sc_hd__inv_2
X_11342_ _01279_ _01280_ VGND VGND VPWR VPWR _01281_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_104_Left_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14061_ _04004_ _04006_ _04031_ VGND VGND VPWR VPWR _04033_ sky130_fd_sc_hd__or3_1
X_11273_ _01169_ _01211_ VGND VGND VPWR VPWR _01212_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10224_ _09197_ _09208_ VGND VGND VPWR VPWR _00163_ sky130_fd_sc_hd__xnor2_1
X_13012_ _02948_ _02949_ VGND VGND VPWR VPWR _02951_ sky130_fd_sc_hd__xor2_1
X_17820_ _08034_ _08035_ VGND VGND VPWR VPWR _08160_ sky130_fd_sc_hd__xnor2_1
X_10155_ _09021_ _09032_ VGND VGND VPWR VPWR _09054_ sky130_fd_sc_hd__nand2_1
X_17751_ net310 _07155_ _07181_ net307 VGND VGND VPWR VPWR _08084_ sky130_fd_sc_hd__a22o_1
X_14963_ _05012_ _05016_ VGND VGND VPWR VPWR _05018_ sky130_fd_sc_hd__xnor2_1
X_10086_ net354 _06062_ _05325_ net357 VGND VGND VPWR VPWR _08295_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16702_ _06927_ _06929_ VGND VGND VPWR VPWR _06930_ sky130_fd_sc_hd__or2b_1
X_13914_ _02468_ _02568_ _03882_ VGND VGND VPWR VPWR _03883_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_89_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17682_ _08001_ _08006_ VGND VGND VPWR VPWR _08008_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_113_Left_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14894_ _04939_ _04941_ net410 kd_2\[0\] VGND VGND VPWR VPWR _04942_ sky130_fd_sc_hd__and4b_1
X_16633_ _06844_ _06851_ _06853_ VGND VGND VPWR VPWR _06855_ sky130_fd_sc_hd__a21oi_1
X_13845_ net266 _02914_ VGND VGND VPWR VPWR _03811_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16564_ net283 _06438_ VGND VGND VPWR VPWR _06779_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13776_ _03739_ _03741_ VGND VGND VPWR VPWR _03742_ sky130_fd_sc_hd__xor2_1
X_10988_ net392 net510 _06029_ VGND VGND VPWR VPWR _00927_ sky130_fd_sc_hd__and3_2
XFILLER_0_146_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18303_ net273 _06336_ _06386_ _06399_ VGND VGND VPWR VPWR _08692_ sky130_fd_sc_hd__a211oi_1
X_15515_ net452 net188 net183 net457 VGND VGND VPWR VPWR _05625_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_128_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12727_ _02664_ _02665_ VGND VGND VPWR VPWR _02666_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19283_ clknet_4_6_0_clock _00061_ VGND VGND VPWR VPWR kp\[13\] sky130_fd_sc_hd__dfxtp_2
X_16495_ _06696_ _06701_ _06702_ VGND VGND VPWR VPWR _06703_ sky130_fd_sc_hd__o21a_1
XFILLER_0_139_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18234_ _06166_ _06168_ _06170_ VGND VGND VPWR VPWR _08616_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15446_ _05521_ _05522_ _05525_ VGND VGND VPWR VPWR _05549_ sky130_fd_sc_hd__o21ai_1
X_12658_ _02595_ _02596_ VGND VGND VPWR VPWR _02597_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11609_ _01535_ _01537_ _01536_ VGND VGND VPWR VPWR _01548_ sky130_fd_sc_hd__a21o_1
X_18165_ _08538_ _08539_ _08478_ VGND VGND VPWR VPWR _08540_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_108_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15377_ _05471_ _05472_ net480 net157 VGND VGND VPWR VPWR _05473_ sky130_fd_sc_hd__and4bb_1
XPHY_EDGE_ROW_122_Left_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12589_ _02475_ _02504_ _02527_ VGND VGND VPWR VPWR _02528_ sky130_fd_sc_hd__o21a_1
X_17116_ _07383_ _07384_ _07385_ VGND VGND VPWR VPWR _07386_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_40_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14328_ net438 net443 net137 net136 VGND VGND VPWR VPWR _04319_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap103 _01688_ VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__buf_6
XFILLER_0_123_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18096_ _07278_ _07423_ VGND VGND VPWR VPWR _08464_ sky130_fd_sc_hd__xnor2_2
Xmax_cap114 _05165_ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17047_ _07297_ _07309_ VGND VGND VPWR VPWR _07310_ sky130_fd_sc_hd__or2b_1
X_14259_ _03971_ _03976_ VGND VGND VPWR VPWR _04243_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18998_ _09150_ _09455_ VGND VGND VPWR VPWR _09456_ sky130_fd_sc_hd__xnor2_1
X_17949_ _08301_ VGND VGND VPWR VPWR _08302_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09998_ net396 net392 _05512_ _05523_ VGND VGND VPWR VPWR _07327_ sky130_fd_sc_hd__and4_2
X_11960_ _01897_ _01898_ VGND VGND VPWR VPWR _01899_ sky130_fd_sc_hd__nor2_1
X_10911_ _00774_ _00849_ VGND VGND VPWR VPWR _00850_ sky130_fd_sc_hd__nor2_1
X_11891_ _01828_ _01829_ VGND VGND VPWR VPWR _01830_ sky130_fd_sc_hd__nor2_1
X_13630_ _03580_ _03586_ _03588_ VGND VGND VPWR VPWR _03589_ sky130_fd_sc_hd__o21ai_2
X_10842_ net367 _09558_ _09565_ VGND VGND VPWR VPWR _00781_ sky130_fd_sc_hd__and3_1
XFILLER_0_156_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13561_ _03393_ _03449_ _03448_ VGND VGND VPWR VPWR _03520_ sky130_fd_sc_hd__o21a_1
X_10773_ net346 _00409_ _00617_ VGND VGND VPWR VPWR _00712_ sky130_fd_sc_hd__and3_1
XFILLER_0_109_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15300_ _05321_ _05332_ _05331_ VGND VGND VPWR VPWR _05388_ sky130_fd_sc_hd__a21o_1
XFILLER_0_67_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12512_ _02446_ _02450_ VGND VGND VPWR VPWR _02451_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16280_ _06463_ _06465_ VGND VGND VPWR VPWR _06466_ sky130_fd_sc_hd__and2_1
X_13492_ net225 _02935_ _03448_ _03450_ VGND VGND VPWR VPWR _03451_ sky130_fd_sc_hd__a31o_1
XFILLER_0_35_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15231_ _05310_ _05311_ VGND VGND VPWR VPWR _05312_ sky130_fd_sc_hd__nor2_1
X_12443_ net226 _01860_ _01835_ net231 VGND VGND VPWR VPWR _02382_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15162_ _05228_ _05230_ _05234_ VGND VGND VPWR VPWR _05236_ sky130_fd_sc_hd__or3_1
X_12374_ _02230_ _02312_ VGND VGND VPWR VPWR _02313_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14113_ _03902_ _03907_ _04083_ VGND VGND VPWR VPWR _04085_ sky130_fd_sc_hd__or3_1
XFILLER_0_50_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11325_ _01254_ _01262_ _01263_ VGND VGND VPWR VPWR _01264_ sky130_fd_sc_hd__a21o_1
X_15093_ _05158_ _05159_ VGND VGND VPWR VPWR _05161_ sky130_fd_sc_hd__nor2_1
X_18921_ _09250_ _09257_ _09255_ VGND VGND VPWR VPWR _09371_ sky130_fd_sc_hd__a21oi_2
X_14044_ prev_d_error\[18\] VGND VGND VPWR VPWR _04016_ sky130_fd_sc_hd__clkinv_4
X_11256_ _01193_ _01194_ VGND VGND VPWR VPWR _01195_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10207_ _09558_ _09565_ VGND VGND VPWR VPWR _09571_ sky130_fd_sc_hd__and2_1
X_18852_ _09293_ _09292_ VGND VGND VPWR VPWR _09295_ sky130_fd_sc_hd__and2b_1
X_11187_ _01115_ _01117_ _01119_ VGND VGND VPWR VPWR _01126_ sky130_fd_sc_hd__o21ba_1
X_10138_ net356 net354 VGND VGND VPWR VPWR _08867_ sky130_fd_sc_hd__or2_1
X_17803_ _08139_ _08140_ VGND VGND VPWR VPWR _08142_ sky130_fd_sc_hd__xor2_1
X_18783_ _09022_ _09201_ VGND VGND VPWR VPWR _09220_ sky130_fd_sc_hd__and2_1
X_15995_ _06149_ _06152_ VGND VGND VPWR VPWR _06153_ sky130_fd_sc_hd__nor2_1
X_17734_ net331 _06618_ _06992_ net314 VGND VGND VPWR VPWR _08066_ sky130_fd_sc_hd__a22o_1
X_10069_ _08097_ _06194_ _06744_ VGND VGND VPWR VPWR _08108_ sky130_fd_sc_hd__o21ba_1
X_14946_ _04895_ _04997_ VGND VGND VPWR VPWR _04999_ sky130_fd_sc_hd__nand2_1
X_17665_ _07986_ _07989_ VGND VGND VPWR VPWR _07990_ sky130_fd_sc_hd__xor2_1
X_14877_ net426 kd_2\[5\] _04860_ _04922_ VGND VGND VPWR VPWR _04923_ sky130_fd_sc_hd__o2bb2a_1
X_16616_ _06751_ _06835_ VGND VGND VPWR VPWR _06836_ sky130_fd_sc_hd__xnor2_2
X_13828_ net257 _02933_ _02914_ net260 VGND VGND VPWR VPWR _03794_ sky130_fd_sc_hd__a22o_1
X_17596_ _07810_ _07813_ VGND VGND VPWR VPWR _07914_ sky130_fd_sc_hd__xnor2_1
X_19335_ clknet_4_2_0_clock _00036_ VGND VGND VPWR VPWR kd_2\[8\] sky130_fd_sc_hd__dfxtp_1
X_16547_ net306 _06310_ VGND VGND VPWR VPWR _06760_ sky130_fd_sc_hd__nand2_1
X_13759_ _03723_ _03724_ VGND VGND VPWR VPWR _03725_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19266_ clknet_4_3_0_clock _00148_ VGND VGND VPWR VPWR prev_d_error\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16478_ _06682_ _06683_ VGND VGND VPWR VPWR _06684_ sky130_fd_sc_hd__and2_1
XFILLER_0_155_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18217_ _08583_ _08594_ _08593_ VGND VGND VPWR VPWR _08597_ sky130_fd_sc_hd__a21boi_1
X_15429_ _05519_ _05521_ _05429_ VGND VGND VPWR VPWR _05530_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_142_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19197_ clknet_4_14_0_clock _00079_ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18148_ _06933_ _07044_ _06837_ VGND VGND VPWR VPWR _08521_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18079_ _07248_ _08444_ VGND VGND VPWR VPWR _08445_ sky130_fd_sc_hd__xnor2_2
X_09921_ net353 _05325_ VGND VGND VPWR VPWR _06480_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09852_ net360 _05006_ VGND VGND VPWR VPWR _05721_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09783_ _04929_ _04951_ VGND VGND VPWR VPWR _04962_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11110_ net396 _05897_ _06150_ VGND VGND VPWR VPWR _01049_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12090_ _02027_ _02028_ VGND VGND VPWR VPWR _02029_ sky130_fd_sc_hd__and2b_1
XFILLER_0_130_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11041_ _00978_ _00979_ VGND VGND VPWR VPWR _00980_ sky130_fd_sc_hd__xor2_2
XFILLER_0_36_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14800_ net421 net175 _04754_ _04755_ VGND VGND VPWR VPWR _04838_ sky130_fd_sc_hd__o2bb2a_1
X_15780_ _04963_ net188 _05895_ net483 net196 VGND VGND VPWR VPWR _05916_ sky130_fd_sc_hd__o2111a_1
X_12992_ _02930_ VGND VGND VPWR VPWR _02931_ sky130_fd_sc_hd__buf_4
X_14731_ _04760_ _04761_ net409 net190 VGND VGND VPWR VPWR _04762_ sky130_fd_sc_hd__and4b_1
X_11943_ net200 _01861_ VGND VGND VPWR VPWR _01882_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17450_ _07737_ _07752_ VGND VGND VPWR VPWR _07753_ sky130_fd_sc_hd__xnor2_1
X_14662_ _04683_ _04685_ VGND VGND VPWR VPWR _04686_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11874_ _01812_ VGND VGND VPWR VPWR _01813_ sky130_fd_sc_hd__clkbuf_4
X_16401_ net296 _06310_ _06598_ VGND VGND VPWR VPWR _06599_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13613_ _03542_ _03571_ VGND VGND VPWR VPWR _03572_ sky130_fd_sc_hd__or2_1
X_17381_ _07263_ _07665_ VGND VGND VPWR VPWR _07677_ sky130_fd_sc_hd__or2_1
X_10825_ net387 _05314_ _04973_ net405 VGND VGND VPWR VPWR _00764_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14593_ _04594_ _04608_ VGND VGND VPWR VPWR _04611_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19120_ _04126_ VGND VGND VPWR VPWR _09550_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16332_ _06420_ _06510_ _06521_ VGND VGND VPWR VPWR _06523_ sky130_fd_sc_hd__nand3_1
X_13544_ net252 _02329_ VGND VGND VPWR VPWR _03503_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10756_ _00693_ _00694_ VGND VGND VPWR VPWR _00695_ sky130_fd_sc_hd__and2b_1
XFILLER_0_137_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19051_ _04126_ net98 VGND VGND VPWR VPWR _09505_ sky130_fd_sc_hd__and2_1
XFILLER_0_152_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16263_ _06445_ _06426_ VGND VGND VPWR VPWR _06448_ sky130_fd_sc_hd__or2b_1
X_13475_ net252 _02223_ _03094_ _03433_ VGND VGND VPWR VPWR _03434_ sky130_fd_sc_hd__a31o_1
XFILLER_0_82_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10687_ _00599_ _00625_ VGND VGND VPWR VPWR _00626_ sky130_fd_sc_hd__xnor2_2
X_18002_ net314 _02931_ _08188_ VGND VGND VPWR VPWR _08360_ sky130_fd_sc_hd__and3_1
X_15214_ _05201_ _05202_ _05291_ VGND VGND VPWR VPWR _05294_ sky130_fd_sc_hd__a21o_1
X_12426_ _02364_ net111 VGND VGND VPWR VPWR _02365_ sky130_fd_sc_hd__and2_1
X_16194_ _06365_ _06371_ VGND VGND VPWR VPWR _06372_ sky130_fd_sc_hd__and2_2
XFILLER_0_106_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15145_ net462 net157 VGND VGND VPWR VPWR _05218_ sky130_fd_sc_hd__nand2_1
X_12357_ _02214_ _02213_ VGND VGND VPWR VPWR _02296_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11308_ _01242_ _01229_ VGND VGND VPWR VPWR _01247_ sky130_fd_sc_hd__nor2_1
X_15076_ net436 net181 VGND VGND VPWR VPWR _05142_ sky130_fd_sc_hd__nand2_1
X_12288_ _02217_ _02226_ VGND VGND VPWR VPWR _02227_ sky130_fd_sc_hd__nor2_1
X_14027_ net411 net156 net151 net416 VGND VGND VPWR VPWR _03999_ sky130_fd_sc_hd__a22oi_1
X_18904_ _09350_ _09225_ _08968_ VGND VGND VPWR VPWR _09353_ sky130_fd_sc_hd__nand3_1
X_11239_ _04621_ _06579_ _04533_ VGND VGND VPWR VPWR _01178_ sky130_fd_sc_hd__or3b_2
X_18835_ _04158_ _09276_ _06004_ _04216_ VGND VGND VPWR VPWR _09277_ sky130_fd_sc_hd__a2bb2o_1
X_18766_ _09011_ _09020_ VGND VGND VPWR VPWR _09201_ sky130_fd_sc_hd__or2_1
X_15978_ _00563_ _01692_ VGND VGND VPWR VPWR _06134_ sky130_fd_sc_hd__xor2_4
XFILLER_0_89_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14929_ _04976_ _04979_ VGND VGND VPWR VPWR _04980_ sky130_fd_sc_hd__nand2_1
X_17717_ _07961_ _07964_ _07963_ VGND VGND VPWR VPWR _08047_ sky130_fd_sc_hd__o21ai_1
X_18697_ _08796_ _08881_ VGND VGND VPWR VPWR _09125_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17648_ _07882_ _07799_ _07881_ VGND VGND VPWR VPWR _07971_ sky130_fd_sc_hd__nand3_1
XFILLER_0_133_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17579_ net315 _06718_ _06719_ VGND VGND VPWR VPWR _07895_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19318_ clknet_4_1_0_clock _00001_ VGND VGND VPWR VPWR kd_1\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19249_ clknet_4_13_0_clock _00131_ VGND VGND VPWR VPWR i_error\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09904_ net338 _06073_ VGND VGND VPWR VPWR _06293_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout502 net504 VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__clkbuf_4
X_09835_ net406 net389 _05512_ _05523_ VGND VGND VPWR VPWR _05534_ sky130_fd_sc_hd__and4_1
X_09766_ net66 net8 VGND VGND VPWR VPWR _04775_ sky130_fd_sc_hd__and2b_1
XFILLER_0_96_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09697_ net41 _03870_ _03903_ net362 VGND VGND VPWR VPWR _00058_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10610_ _00529_ _00547_ _00548_ VGND VGND VPWR VPWR _00549_ sky130_fd_sc_hd__a21oi_1
X_11590_ net400 _00244_ _01528_ _01487_ VGND VGND VPWR VPWR _01529_ sky130_fd_sc_hd__nand4_1
XFILLER_0_92_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10541_ _00473_ _00470_ VGND VGND VPWR VPWR _00480_ sky130_fd_sc_hd__or2b_1
XFILLER_0_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13260_ _03206_ _03211_ VGND VGND VPWR VPWR _03213_ sky130_fd_sc_hd__or2b_1
XFILLER_0_150_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10472_ net343 _00244_ _00324_ net340 VGND VGND VPWR VPWR _00411_ sky130_fd_sc_hd__a22o_1
X_12211_ _01930_ _02148_ _02149_ VGND VGND VPWR VPWR _02150_ sky130_fd_sc_hd__a21oi_1
X_13191_ net263 _01806_ VGND VGND VPWR VPWR _03144_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12142_ net200 _01910_ _01911_ _01913_ VGND VGND VPWR VPWR _02081_ sky130_fd_sc_hd__a22o_1
X_12073_ _01777_ _01781_ VGND VGND VPWR VPWR _02012_ sky130_fd_sc_hd__xnor2_1
X_16950_ net302 _06620_ _07193_ VGND VGND VPWR VPWR _07203_ sky130_fd_sc_hd__and3_1
X_15901_ _04998_ _05962_ VGND VGND VPWR VPWR _06049_ sky130_fd_sc_hd__xor2_1
X_11024_ net396 _05963_ _05974_ _00927_ VGND VGND VPWR VPWR _00963_ sky130_fd_sc_hd__and4_1
X_16881_ _07049_ _07126_ VGND VGND VPWR VPWR _07127_ sky130_fd_sc_hd__xnor2_2
X_15832_ _05971_ _05969_ _04673_ VGND VGND VPWR VPWR _05973_ sky130_fd_sc_hd__nor3_1
X_18620_ _09036_ _09039_ VGND VGND VPWR VPWR _09040_ sky130_fd_sc_hd__and2b_1
XFILLER_0_154_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15763_ net480 net188 VGND VGND VPWR VPWR _05898_ sky130_fd_sc_hd__nand2_1
X_18551_ _08963_ VGND VGND VPWR VPWR _08964_ sky130_fd_sc_hd__clkbuf_4
X_12975_ _02913_ VGND VGND VPWR VPWR _02914_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14714_ _04740_ _04743_ VGND VGND VPWR VPWR _04744_ sky130_fd_sc_hd__nand2_1
X_17502_ net301 _06992_ VGND VGND VPWR VPWR _07810_ sky130_fd_sc_hd__nand2_1
X_11926_ net200 _01854_ _01863_ VGND VGND VPWR VPWR _01865_ sky130_fd_sc_hd__a21oi_1
X_18482_ net101 _06175_ VGND VGND VPWR VPWR _08888_ sky130_fd_sc_hd__nor2_1
X_15694_ _05788_ _05821_ VGND VGND VPWR VPWR _05822_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17433_ _07638_ _07650_ VGND VGND VPWR VPWR _07735_ sky130_fd_sc_hd__nor2_1
X_14645_ _04536_ _04551_ _04549_ VGND VGND VPWR VPWR _04668_ sky130_fd_sc_hd__a21oi_1
X_11857_ _01702_ _01795_ VGND VGND VPWR VPWR _01796_ sky130_fd_sc_hd__nand2_2
XFILLER_0_157_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17364_ net290 _07570_ VGND VGND VPWR VPWR _07659_ sky130_fd_sc_hd__nand2_1
X_10808_ _00721_ _00746_ VGND VGND VPWR VPWR _00747_ sky130_fd_sc_hd__xor2_1
X_14576_ _04590_ _04591_ VGND VGND VPWR VPWR _04592_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11788_ _01724_ _00322_ VGND VGND VPWR VPWR _01727_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16315_ _06376_ _06503_ VGND VGND VPWR VPWR _06505_ sky130_fd_sc_hd__nor2_1
X_19103_ _09536_ _06073_ _09539_ net488 VGND VGND VPWR VPWR _00107_ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13527_ _03480_ _03484_ _03384_ _03485_ VGND VGND VPWR VPWR _03486_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17295_ _07550_ _07581_ _07582_ VGND VGND VPWR VPWR _07583_ sky130_fd_sc_hd__o21a_1
X_10739_ _00677_ VGND VGND VPWR VPWR _00678_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19034_ _09448_ _09485_ _09470_ VGND VGND VPWR VPWR _09493_ sky130_fd_sc_hd__a21oi_1
X_16246_ _06428_ _06415_ VGND VGND VPWR VPWR _06429_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13458_ _03344_ _03416_ VGND VGND VPWR VPWR _03417_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12409_ _02244_ _02346_ _02306_ _02345_ VGND VGND VPWR VPWR _02348_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_106_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16177_ _06352_ VGND VGND VPWR VPWR _06353_ sky130_fd_sc_hd__buf_2
XFILLER_0_23_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13389_ _03330_ _03329_ _03305_ VGND VGND VPWR VPWR _03343_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15128_ _05104_ _05197_ VGND VGND VPWR VPWR _05199_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15059_ _05111_ _05120_ _05122_ VGND VGND VPWR VPWR _05123_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09620_ net58 _03102_ _03135_ net155 VGND VGND VPWR VPWR _00037_ sky130_fd_sc_hd__a22o_1
X_18818_ _09250_ _09257_ VGND VGND VPWR VPWR _09258_ sky130_fd_sc_hd__xnor2_1
X_18749_ _09166_ _09174_ _09173_ VGND VGND VPWR VPWR _09182_ sky130_fd_sc_hd__a21o_2
XFILLER_0_78_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout310 ki\[6\] VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__buf_4
Xfanout321 ki\[3\] VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout332 net566 VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__clkbuf_4
Xfanout343 kp\[15\] VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__clkbuf_4
Xfanout354 kp\[13\] VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__clkbuf_4
Xfanout365 kp\[10\] VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__clkbuf_4
Xfanout376 kp\[7\] VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__buf_2
X_09818_ net348 _05336_ VGND VGND VPWR VPWR _05347_ sky130_fd_sc_hd__nand2_1
Xfanout387 net388 VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__buf_2
Xfanout398 kp\[2\] VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__buf_4
X_09749_ net61 net3 VGND VGND VPWR VPWR _04588_ sky130_fd_sc_hd__or2b_1
XFILLER_0_96_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12760_ net250 _02698_ _01764_ VGND VGND VPWR VPWR _02699_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11711_ net394 _00812_ _01638_ VGND VGND VPWR VPWR _01650_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12691_ _02608_ _02609_ _02629_ VGND VGND VPWR VPWR _02630_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_84_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14430_ _04408_ _04385_ VGND VGND VPWR VPWR _04431_ sky130_fd_sc_hd__or2b_1
X_11642_ _01525_ _01540_ _01544_ VGND VGND VPWR VPWR _01581_ sky130_fd_sc_hd__and3_1
XFILLER_0_154_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14361_ _04350_ _04354_ VGND VGND VPWR VPWR _04355_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11573_ _01510_ _01511_ VGND VGND VPWR VPWR _01512_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput18 measurement[7] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
X_16100_ _06175_ _06266_ _06267_ VGND VGND VPWR VPWR _06268_ sky130_fd_sc_hd__or3_1
XFILLER_0_92_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13312_ _03263_ _03264_ VGND VGND VPWR VPWR _03265_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput29 reg_addr[17] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10524_ _00269_ _00353_ VGND VGND VPWR VPWR _00463_ sky130_fd_sc_hd__xor2_4
X_17080_ _07310_ _07314_ _07344_ _07345_ VGND VGND VPWR VPWR _07346_ sky130_fd_sc_hd__a211o_1
X_14292_ _04245_ _04248_ _04278_ VGND VGND VPWR VPWR _04279_ sky130_fd_sc_hd__a21o_1
XFILLER_0_150_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16031_ _08636_ _08669_ _06190_ VGND VGND VPWR VPWR _06192_ sky130_fd_sc_hd__nor3_1
X_13243_ _03189_ _03191_ _03194_ VGND VGND VPWR VPWR _03196_ sky130_fd_sc_hd__and3_1
X_10455_ _08097_ _00245_ _00341_ VGND VGND VPWR VPWR _00394_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_149_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13174_ _03071_ _03125_ VGND VGND VPWR VPWR _03126_ sky130_fd_sc_hd__nor2_1
X_10386_ _00324_ VGND VGND VPWR VPWR _00325_ sky130_fd_sc_hd__buf_2
X_12125_ _01900_ _02063_ VGND VGND VPWR VPWR _02064_ sky130_fd_sc_hd__nor2_1
X_17982_ _08337_ VGND VGND VPWR VPWR _08338_ sky130_fd_sc_hd__inv_2
X_16933_ _07158_ _07180_ VGND VGND VPWR VPWR _07185_ sky130_fd_sc_hd__xor2_1
X_12056_ _01993_ _01994_ VGND VGND VPWR VPWR _01995_ sky130_fd_sc_hd__nor2_1
X_11007_ _00854_ _00830_ _00853_ VGND VGND VPWR VPWR _00946_ sky130_fd_sc_hd__and3_1
X_16864_ _07106_ _07108_ VGND VGND VPWR VPWR _07109_ sky130_fd_sc_hd__nor2_1
X_18603_ _09011_ _09020_ VGND VGND VPWR VPWR _09022_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15815_ _05295_ _05954_ _05293_ VGND VGND VPWR VPWR _05955_ sky130_fd_sc_hd__o21a_1
X_16795_ _07011_ _07028_ _07032_ VGND VGND VPWR VPWR _07033_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15746_ _05874_ _05877_ _05878_ VGND VGND VPWR VPWR _05879_ sky130_fd_sc_hd__and3_1
X_18534_ _08921_ VGND VGND VPWR VPWR _08946_ sky130_fd_sc_hd__inv_2
X_12958_ net228 _02221_ _02088_ net233 VGND VGND VPWR VPWR _02897_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11909_ _01847_ VGND VGND VPWR VPWR _01848_ sky130_fd_sc_hd__buf_4
XFILLER_0_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15677_ _05801_ _05802_ net478 net179 VGND VGND VPWR VPWR _05803_ sky130_fd_sc_hd__and4bb_1
X_18465_ _08685_ _08683_ _08684_ VGND VGND VPWR VPWR _08870_ sky130_fd_sc_hd__nand3_2
X_12889_ net211 _02410_ VGND VGND VPWR VPWR _02828_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14628_ _04646_ _04648_ VGND VGND VPWR VPWR _04649_ sky130_fd_sc_hd__xnor2_1
X_17416_ _07619_ _07627_ VGND VGND VPWR VPWR _07716_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18396_ _06149_ _08793_ VGND VGND VPWR VPWR _08794_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17347_ net299 _06802_ VGND VGND VPWR VPWR _07640_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14559_ _04570_ _04572_ VGND VGND VPWR VPWR _04573_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17278_ net290 _07156_ VGND VGND VPWR VPWR _07564_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16229_ _06409_ VGND VGND VPWR VPWR _06410_ sky130_fd_sc_hd__clkbuf_4
X_19017_ _09462_ _09464_ _09465_ _09476_ VGND VGND VPWR VPWR _09477_ sky130_fd_sc_hd__and4_1
XFILLER_0_140_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_143_Right_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09603_ _02992_ _03047_ VGND VGND VPWR VPWR _03058_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10240_ _00176_ _00174_ VGND VGND VPWR VPWR _00179_ sky130_fd_sc_hd__xnor2_1
X_10171_ _07932_ _07943_ VGND VGND VPWR VPWR _09230_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_110_Right_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout140 kd_2\[13\] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_4
Xfanout151 kd_2\[10\] VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_4
Xfanout162 net163 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__buf_2
X_13930_ net448 net116 VGND VGND VPWR VPWR _03900_ sky130_fd_sc_hd__nand2_1
Xfanout173 net174 VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_2
Xfanout184 net185 VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_4
Xfanout195 net196 VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__buf_2
X_13861_ _03792_ _03811_ VGND VGND VPWR VPWR _03827_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15600_ _05713_ _05714_ _05716_ VGND VGND VPWR VPWR _05718_ sky130_fd_sc_hd__and3_1
X_12812_ net204 _02545_ _02750_ VGND VGND VPWR VPWR _02751_ sky130_fd_sc_hd__and3_1
X_16580_ _06727_ _06728_ VGND VGND VPWR VPWR _06796_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13792_ net243 _02934_ _03757_ VGND VGND VPWR VPWR _03758_ sky130_fd_sc_hd__and3_1
XFILLER_0_139_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15531_ _05618_ VGND VGND VPWR VPWR _05642_ sky130_fd_sc_hd__inv_2
X_12743_ _02579_ _02578_ VGND VGND VPWR VPWR _02682_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18250_ net273 _06386_ VGND VGND VPWR VPWR _08633_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15462_ _05485_ _05565_ VGND VGND VPWR VPWR _05566_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12674_ net233 VGND VGND VPWR VPWR _02613_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17201_ _07464_ _07465_ _07476_ _07477_ VGND VGND VPWR VPWR _07479_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14413_ _04410_ _04411_ net435 net146 VGND VGND VPWR VPWR _04413_ sky130_fd_sc_hd__and4bb_1
X_11625_ _01356_ _01550_ VGND VGND VPWR VPWR _01564_ sky130_fd_sc_hd__nand2_1
X_18181_ _08167_ _08168_ _08429_ VGND VGND VPWR VPWR _08557_ sky130_fd_sc_hd__and3_1
X_15393_ _05397_ _05489_ VGND VGND VPWR VPWR _05491_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17132_ _07392_ _07402_ VGND VGND VPWR VPWR _07403_ sky130_fd_sc_hd__xnor2_2
X_14344_ _04326_ _04330_ _04334_ _04336_ VGND VGND VPWR VPWR _04337_ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11556_ _01469_ _01474_ VGND VGND VPWR VPWR _01495_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10507_ _00438_ _00445_ VGND VGND VPWR VPWR _00446_ sky130_fd_sc_hd__or2b_1
X_17063_ _07319_ _07320_ _07326_ VGND VGND VPWR VPWR _07328_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_150_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14275_ net407 net160 _03998_ _03999_ VGND VGND VPWR VPWR _04261_ sky130_fd_sc_hd__o2bb2a_1
X_11487_ _01365_ _01422_ _01425_ VGND VGND VPWR VPWR _01426_ sky130_fd_sc_hd__o21ai_2
X_16014_ _06131_ _06173_ VGND VGND VPWR VPWR _06174_ sky130_fd_sc_hd__and2b_1
X_13226_ _03084_ _03092_ _03176_ VGND VGND VPWR VPWR _03179_ sky130_fd_sc_hd__o21ai_1
X_10438_ _00296_ _00376_ VGND VGND VPWR VPWR _00377_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13157_ _03034_ _03106_ VGND VGND VPWR VPWR _03107_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10369_ _00283_ _00282_ VGND VGND VPWR VPWR _00308_ sky130_fd_sc_hd__and2b_1
X_12108_ _02039_ _02042_ VGND VGND VPWR VPWR _02047_ sky130_fd_sc_hd__or2b_1
X_13088_ _03026_ _03030_ VGND VGND VPWR VPWR _03031_ sky130_fd_sc_hd__xor2_1
X_17965_ net331 _06991_ _07568_ net314 VGND VGND VPWR VPWR _08320_ sky130_fd_sc_hd__a22o_1
X_16916_ net288 _06724_ _07165_ VGND VGND VPWR VPWR _07166_ sky130_fd_sc_hd__a21bo_1
X_12039_ _01975_ _01977_ VGND VGND VPWR VPWR _01978_ sky130_fd_sc_hd__nor2_2
X_17896_ _08232_ _08242_ _08243_ VGND VGND VPWR VPWR _08244_ sky130_fd_sc_hd__o21a_1
X_16847_ net285 _06724_ _06980_ _07089_ VGND VGND VPWR VPWR _07090_ sky130_fd_sc_hd__a31o_1
X_16778_ net329 _06324_ VGND VGND VPWR VPWR _07014_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18517_ _08925_ _08785_ VGND VGND VPWR VPWR _08927_ sky130_fd_sc_hd__and2_1
X_15729_ _05859_ VGND VGND VPWR VPWR _05860_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18448_ _08590_ _08850_ VGND VGND VPWR VPWR _08851_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_91_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18379_ _08772_ _08774_ VGND VGND VPWR VPWR _08775_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_43_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclone3 net562 _04687_ _04698_ VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__o21ai_2
XFILLER_0_79_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11410_ _01277_ _01276_ _01244_ VGND VGND VPWR VPWR _01349_ sky130_fd_sc_hd__a21oi_1
X_12390_ _02326_ _02328_ VGND VGND VPWR VPWR _02329_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_61_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11341_ _01136_ _01206_ VGND VGND VPWR VPWR _01280_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_34_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14060_ _04004_ _04006_ _04031_ VGND VGND VPWR VPWR _04032_ sky130_fd_sc_hd__o21ai_2
X_11272_ _01204_ _01203_ VGND VGND VPWR VPWR _01211_ sky130_fd_sc_hd__or2b_1
XFILLER_0_39_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13011_ _02948_ _02949_ VGND VGND VPWR VPWR _02950_ sky130_fd_sc_hd__nor2_1
X_10223_ _07778_ _07800_ VGND VGND VPWR VPWR _00162_ sky130_fd_sc_hd__xnor2_1
X_10154_ _09021_ _09032_ VGND VGND VPWR VPWR _09043_ sky130_fd_sc_hd__or2_1
X_14962_ _05013_ _05014_ _05015_ VGND VGND VPWR VPWR _05016_ sky130_fd_sc_hd__o21ba_1
X_17750_ _08071_ _08081_ VGND VGND VPWR VPWR _08083_ sky130_fd_sc_hd__xnor2_2
X_10085_ net353 _05325_ _08273_ VGND VGND VPWR VPWR _08284_ sky130_fd_sc_hd__and3_1
X_16701_ _06875_ _06928_ VGND VGND VPWR VPWR _06929_ sky130_fd_sc_hd__nand2_1
X_13913_ _02673_ _03879_ _03880_ VGND VGND VPWR VPWR _03882_ sky130_fd_sc_hd__a21oi_1
X_14893_ net414 net194 net190 net417 VGND VGND VPWR VPWR _04941_ sky130_fd_sc_hd__a22o_1
X_17681_ _08001_ _08006_ VGND VGND VPWR VPWR _08007_ sky130_fd_sc_hd__nand2_1
X_16632_ _06781_ _06852_ VGND VGND VPWR VPWR _06853_ sky130_fd_sc_hd__or2_1
X_13844_ _03793_ _03795_ VGND VGND VPWR VPWR _03810_ sky130_fd_sc_hd__xor2_1
X_16563_ _06772_ _06776_ VGND VGND VPWR VPWR _06778_ sky130_fd_sc_hd__xnor2_1
X_13775_ _03624_ _03740_ _03698_ VGND VGND VPWR VPWR _03741_ sky130_fd_sc_hd__a21oi_1
X_10987_ _00835_ _00838_ VGND VGND VPWR VPWR _00926_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18302_ _08630_ _08645_ _08643_ VGND VGND VPWR VPWR _08690_ sky130_fd_sc_hd__a21oi_1
X_15514_ net450 net192 VGND VGND VPWR VPWR _05624_ sky130_fd_sc_hd__nand2_1
X_12726_ _02575_ _02628_ VGND VGND VPWR VPWR _02665_ sky130_fd_sc_hd__xor2_1
XFILLER_0_84_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19282_ clknet_4_6_0_clock _00060_ VGND VGND VPWR VPWR kp\[12\] sky130_fd_sc_hd__dfxtp_1
X_16494_ _06697_ _06699_ VGND VGND VPWR VPWR _06702_ sky130_fd_sc_hd__or2b_1
XFILLER_0_155_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15445_ _05542_ _05547_ VGND VGND VPWR VPWR _05548_ sky130_fd_sc_hd__nand2_1
X_18233_ _08527_ _08613_ VGND VGND VPWR VPWR _08615_ sky130_fd_sc_hd__xor2_2
XFILLER_0_128_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12657_ _02592_ _02594_ VGND VGND VPWR VPWR _02596_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11608_ _01523_ _01546_ VGND VGND VPWR VPWR _01547_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15376_ net472 net167 net162 net476 VGND VGND VPWR VPWR _05472_ sky130_fd_sc_hd__a22oi_1
X_18164_ _07974_ _08440_ _08491_ _08494_ VGND VGND VPWR VPWR _08539_ sky130_fd_sc_hd__a211o_1
X_12588_ _02525_ _02526_ VGND VGND VPWR VPWR _02527_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17115_ _07381_ _07352_ VGND VGND VPWR VPWR _07385_ sky130_fd_sc_hd__and2b_1
X_14327_ _04306_ _04317_ VGND VGND VPWR VPWR _04318_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11539_ _01388_ _01477_ VGND VGND VPWR VPWR _01478_ sky130_fd_sc_hd__and2b_1
X_18095_ _08450_ _08461_ _08462_ VGND VGND VPWR VPWR _08463_ sky130_fd_sc_hd__a21o_1
Xmax_cap104 _03328_ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_1
Xmax_cap115 _01906_ VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__buf_4
X_17046_ _07303_ _07308_ VGND VGND VPWR VPWR _07309_ sky130_fd_sc_hd__nand2_1
X_14258_ _04239_ _04241_ VGND VGND VPWR VPWR _04242_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13209_ _03121_ _03119_ VGND VGND VPWR VPWR _03162_ sky130_fd_sc_hd__and2b_1
XFILLER_0_111_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14189_ net412 net130 net124 net418 VGND VGND VPWR VPWR _04166_ sky130_fd_sc_hd__a22o_1
X_18997_ _09165_ _09454_ _09162_ VGND VGND VPWR VPWR _09455_ sky130_fd_sc_hd__o21ba_1
X_17948_ _08265_ _08300_ VGND VGND VPWR VPWR _08301_ sky130_fd_sc_hd__nor2_1
X_17879_ net322 _07093_ _07155_ net318 VGND VGND VPWR VPWR _08225_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_45_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09997_ net384 _07294_ _07305_ VGND VGND VPWR VPWR _07316_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_99_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10910_ _00773_ _00772_ VGND VGND VPWR VPWR _00849_ sky130_fd_sc_hd__and2b_1
X_11890_ net230 _01787_ _01799_ net226 VGND VGND VPWR VPWR _01829_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_86_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10841_ net363 _09577_ _08196_ net366 VGND VGND VPWR VPWR _00780_ sky130_fd_sc_hd__a22oi_1
X_13560_ net225 _02934_ VGND VGND VPWR VPWR _03519_ sky130_fd_sc_hd__nand2_1
X_10772_ net346 _00409_ _00617_ VGND VGND VPWR VPWR _00711_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12511_ _02440_ _02445_ VGND VGND VPWR VPWR _02450_ sky130_fd_sc_hd__nor2_1
X_13491_ _03393_ _03449_ VGND VGND VPWR VPWR _03450_ sky130_fd_sc_hd__nor2_1
X_15230_ net468 net486 net158 net139 VGND VGND VPWR VPWR _05311_ sky130_fd_sc_hd__and4_1
X_12442_ _02285_ _02380_ VGND VGND VPWR VPWR _02381_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15161_ _05228_ _05230_ _05234_ VGND VGND VPWR VPWR _05235_ sky130_fd_sc_hd__o21ai_1
X_12373_ _02217_ _02228_ _02229_ VGND VGND VPWR VPWR _02312_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14112_ _03902_ _03907_ _04083_ VGND VGND VPWR VPWR _04084_ sky130_fd_sc_hd__o21ai_1
X_11324_ _01256_ _01261_ VGND VGND VPWR VPWR _01263_ sky130_fd_sc_hd__and2b_1
XFILLER_0_22_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15092_ _05154_ _05155_ _05157_ VGND VGND VPWR VPWR _05159_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14043_ _03997_ _04003_ _04014_ VGND VGND VPWR VPWR _04015_ sky130_fd_sc_hd__a21oi_2
X_18920_ _01929_ _09314_ _09316_ VGND VGND VPWR VPWR _09370_ sky130_fd_sc_hd__o21a_1
X_11255_ _01163_ _01165_ VGND VGND VPWR VPWR _01194_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_31_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10206_ _04412_ _04357_ _09552_ _04478_ VGND VGND VPWR VPWR _09565_ sky130_fd_sc_hd__nand4_4
X_18851_ _09292_ _09293_ VGND VGND VPWR VPWR _09294_ sky130_fd_sc_hd__and2b_1
X_11186_ _01123_ _01124_ VGND VGND VPWR VPWR _01125_ sky130_fd_sc_hd__and2b_1
X_17802_ _08022_ _08023_ VGND VGND VPWR VPWR _08140_ sky130_fd_sc_hd__xnor2_1
X_10137_ _08845_ _07481_ _06887_ VGND VGND VPWR VPWR _08856_ sky130_fd_sc_hd__o21ba_1
X_18782_ _09216_ _09217_ VGND VGND VPWR VPWR _09218_ sky130_fd_sc_hd__or2_1
X_15994_ _06143_ _06151_ _01677_ VGND VGND VPWR VPWR _06152_ sky130_fd_sc_hd__mux2_2
X_17733_ _08057_ _08058_ _08062_ VGND VGND VPWR VPWR _08065_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14945_ _04895_ _04997_ VGND VGND VPWR VPWR _04998_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10068_ _08086_ VGND VGND VPWR VPWR _08097_ sky130_fd_sc_hd__buf_4
X_17664_ _07462_ _07988_ VGND VGND VPWR VPWR _07989_ sky130_fd_sc_hd__xor2_1
X_14876_ _04861_ VGND VGND VPWR VPWR _04922_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16615_ _06752_ _06834_ VGND VGND VPWR VPWR _06835_ sky130_fd_sc_hd__nor2_1
X_13827_ net266 _02746_ VGND VGND VPWR VPWR _03793_ sky130_fd_sc_hd__nand2_1
X_17595_ _07894_ _07896_ _07898_ VGND VGND VPWR VPWR _07913_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_147_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19334_ clknet_4_2_0_clock _00035_ VGND VGND VPWR VPWR kd_2\[7\] sky130_fd_sc_hd__dfxtp_1
X_13758_ net260 _02639_ _02745_ net256 VGND VGND VPWR VPWR _03724_ sky130_fd_sc_hd__a22oi_1
X_16546_ net309 _06316_ _06318_ VGND VGND VPWR VPWR _06759_ sky130_fd_sc_hd__and3_1
X_12709_ net215 _02224_ _02090_ net219 VGND VGND VPWR VPWR _02648_ sky130_fd_sc_hd__a22o_1
X_19265_ clknet_4_3_0_clock _00147_ VGND VGND VPWR VPWR prev_d_error\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13689_ _03653_ VGND VGND VPWR VPWR _03654_ sky130_fd_sc_hd__inv_2
X_16477_ _06675_ _06680_ _06681_ VGND VGND VPWR VPWR _06683_ sky130_fd_sc_hd__or3_1
XFILLER_0_38_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18216_ _08585_ _08587_ _08590_ _08595_ VGND VGND VPWR VPWR _08596_ sky130_fd_sc_hd__or4_4
X_15428_ _05528_ VGND VGND VPWR VPWR _05529_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19196_ clknet_4_14_0_clock _00078_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15359_ _05439_ _05442_ _05451_ VGND VGND VPWR VPWR _05453_ sky130_fd_sc_hd__and3_1
X_18147_ _07154_ _08513_ _08518_ _08519_ VGND VGND VPWR VPWR _08520_ sky130_fd_sc_hd__a31o_2
XFILLER_0_124_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18078_ _07273_ _07271_ VGND VGND VPWR VPWR _08444_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09920_ net348 _06073_ VGND VGND VPWR VPWR _06469_ sky130_fd_sc_hd__nand2_1
X_17029_ net312 _06345_ VGND VGND VPWR VPWR _07290_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09851_ _05083_ _05699_ _05600_ VGND VGND VPWR VPWR _05710_ sky130_fd_sc_hd__and3b_1
XFILLER_0_0_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09782_ _04940_ VGND VGND VPWR VPWR _04951_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_141_Left_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11040_ _00880_ _00879_ VGND VGND VPWR VPWR _00979_ sky130_fd_sc_hd__and2b_1
X_12991_ _02928_ _02929_ VGND VGND VPWR VPWR _02930_ sky130_fd_sc_hd__and2_1
X_11942_ net208 _01808_ _01819_ _01816_ VGND VGND VPWR VPWR _01881_ sky130_fd_sc_hd__a31o_1
X_14730_ net413 net186 _04565_ VGND VGND VPWR VPWR _04761_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14661_ _04683_ _04684_ net475 net125 VGND VGND VPWR VPWR _04685_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_98_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11873_ _01811_ _01748_ VGND VGND VPWR VPWR _01812_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_157_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13612_ _03521_ _03522_ VGND VGND VPWR VPWR _03571_ sky130_fd_sc_hd__nor2_1
X_16400_ net300 _06335_ VGND VGND VPWR VPWR _06598_ sky130_fd_sc_hd__and2_1
X_10824_ _00673_ _00762_ VGND VGND VPWR VPWR _00763_ sky130_fd_sc_hd__xnor2_1
X_14592_ _04594_ _04608_ VGND VGND VPWR VPWR _04609_ sky130_fd_sc_hd__and2_1
X_17380_ net273 _02933_ VGND VGND VPWR VPWR _07676_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13543_ net269 _01873_ VGND VGND VPWR VPWR _03502_ sky130_fd_sc_hd__nand2_1
X_16331_ _06420_ _06510_ _06521_ VGND VGND VPWR VPWR _06522_ sky130_fd_sc_hd__a21o_1
XFILLER_0_67_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10755_ _00680_ _00681_ VGND VGND VPWR VPWR _00694_ sky130_fd_sc_hd__xnor2_1
X_19050_ _09503_ _09504_ net492 VGND VGND VPWR VPWR _00084_ sky130_fd_sc_hd__o21a_1
X_16262_ _06426_ _06445_ VGND VGND VPWR VPWR _06446_ sky130_fd_sc_hd__or2b_1
X_13474_ net249 _03432_ _02331_ VGND VGND VPWR VPWR _03433_ sky130_fd_sc_hd__and3_1
X_10686_ _00601_ _00623_ _00624_ VGND VGND VPWR VPWR _00625_ sky130_fd_sc_hd__o21ba_1
X_15213_ _05201_ _05202_ _05291_ VGND VGND VPWR VPWR _05293_ sky130_fd_sc_hd__nand3_1
XFILLER_0_63_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18001_ net314 _02931_ _08188_ VGND VGND VPWR VPWR _08359_ sky130_fd_sc_hd__a21oi_1
X_12425_ net268 net250 _01759_ VGND VGND VPWR VPWR _02364_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16193_ net303 _06367_ _06369_ _06328_ VGND VGND VPWR VPWR _06371_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15144_ _05214_ _04801_ _05216_ VGND VGND VPWR VPWR _05217_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_152_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12356_ net208 _01875_ VGND VGND VPWR VPWR _02295_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11307_ _01193_ _01194_ VGND VGND VPWR VPWR _01246_ sky130_fd_sc_hd__xor2_4
X_15075_ net441 net178 net172 net446 VGND VGND VPWR VPWR _05141_ sky130_fd_sc_hd__a22oi_2
X_12287_ _02225_ _02210_ _02083_ VGND VGND VPWR VPWR _02226_ sky130_fd_sc_hd__o21a_1
XFILLER_0_121_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14026_ net411 net416 net156 net151 VGND VGND VPWR VPWR _03998_ sky130_fd_sc_hd__and4_1
X_18903_ _09225_ _08968_ _09350_ VGND VGND VPWR VPWR _09352_ sky130_fd_sc_hd__a21oi_1
X_11238_ net402 _05963_ _05974_ VGND VGND VPWR VPWR _01177_ sky130_fd_sc_hd__and3_1
X_18834_ _04216_ _06003_ VGND VGND VPWR VPWR _09276_ sky130_fd_sc_hd__nor2_1
X_11169_ _01106_ _01024_ VGND VGND VPWR VPWR _01108_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18765_ _09044_ _09198_ _09199_ VGND VGND VPWR VPWR _09200_ sky130_fd_sc_hd__a21o_1
X_15977_ _00268_ _06132_ VGND VGND VPWR VPWR _06133_ sky130_fd_sc_hd__xnor2_4
X_17716_ _08038_ _08044_ _08045_ VGND VGND VPWR VPWR _08046_ sky130_fd_sc_hd__nor3_2
XFILLER_0_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14928_ _04976_ _04977_ _04978_ VGND VGND VPWR VPWR _04979_ sky130_fd_sc_hd__nand3_1
X_18696_ _06089_ _09123_ VGND VGND VPWR VPWR _09124_ sky130_fd_sc_hd__nor2_2
XFILLER_0_26_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17647_ _07882_ _07881_ _07799_ VGND VGND VPWR VPWR _07970_ sky130_fd_sc_hd__a21o_1
X_14859_ net449 net159 VGND VGND VPWR VPWR _04903_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17578_ net313 _06802_ VGND VGND VPWR VPWR _07894_ sky130_fd_sc_hd__nand2_1
X_19317_ clknet_4_1_0_clock _00018_ VGND VGND VPWR VPWR kd_1\[9\] sky130_fd_sc_hd__dfxtp_1
X_16529_ _06648_ _06662_ VGND VGND VPWR VPWR _06740_ sky130_fd_sc_hd__xor2_1
XFILLER_0_144_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19248_ clknet_4_15_0_clock _00130_ VGND VGND VPWR VPWR i_error\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19179_ net502 net436 net491 _09586_ VGND VGND VPWR VPWR _00144_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09903_ net338 _06007_ _06106_ _06084_ VGND VGND VPWR VPWR _06282_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout503 net504 VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09834_ _04929_ _05017_ _05501_ VGND VGND VPWR VPWR _05523_ sky130_fd_sc_hd__a21o_4
X_09765_ _04181_ _04709_ _04720_ _04731_ _04753_ VGND VGND VPWR VPWR _04764_ sky130_fd_sc_hd__a311o_4
X_09696_ net58 _03881_ _03914_ net366 VGND VGND VPWR VPWR _00075_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10540_ _00475_ _00476_ _00478_ VGND VGND VPWR VPWR _00479_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_33_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10471_ _00409_ VGND VGND VPWR VPWR _00410_ sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_157_Right_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12210_ net218 _01772_ _01930_ net215 VGND VGND VPWR VPWR _02149_ sky130_fd_sc_hd__a22oi_1
X_13190_ _02998_ _02948_ _02997_ VGND VGND VPWR VPWR _03143_ sky130_fd_sc_hd__o21a_1
X_12141_ _02076_ _02079_ VGND VGND VPWR VPWR _02080_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12072_ _01978_ _01981_ VGND VGND VPWR VPWR _02011_ sky130_fd_sc_hd__nor2_2
XFILLER_0_47_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15900_ _03869_ _06047_ VGND VGND VPWR VPWR _06048_ sky130_fd_sc_hd__and2_1
X_11023_ _00928_ _00961_ VGND VGND VPWR VPWR _00962_ sky130_fd_sc_hd__xnor2_4
X_16880_ _06364_ _06310_ _07050_ VGND VGND VPWR VPWR _07126_ sky130_fd_sc_hd__a21oi_1
X_15831_ _05969_ _04673_ _05971_ VGND VGND VPWR VPWR _05972_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18550_ _08961_ _08962_ VGND VGND VPWR VPWR _08963_ sky130_fd_sc_hd__nand2_2
X_15762_ net474 net196 _05895_ VGND VGND VPWR VPWR _05896_ sky130_fd_sc_hd__and3_1
X_12974_ _01716_ _01717_ VGND VGND VPWR VPWR _02913_ sky130_fd_sc_hd__xor2_4
XFILLER_0_99_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17501_ _06900_ _07808_ net307 VGND VGND VPWR VPWR _07809_ sky130_fd_sc_hd__or3b_1
X_14713_ _04721_ _04741_ VGND VGND VPWR VPWR _04743_ sky130_fd_sc_hd__and2_1
X_11925_ net200 _01854_ _01863_ VGND VGND VPWR VPWR _01864_ sky130_fd_sc_hd__and3_1
X_18481_ net101 _06174_ _01698_ VGND VGND VPWR VPWR _08887_ sky130_fd_sc_hd__and3_1
X_15693_ _05796_ _05818_ _05819_ VGND VGND VPWR VPWR _05821_ sky130_fd_sc_hd__a21oi_1
X_17432_ _07730_ _07731_ _07693_ _07653_ VGND VGND VPWR VPWR _07733_ sky130_fd_sc_hd__o211ai_2
X_14644_ _04664_ _04666_ VGND VGND VPWR VPWR _04667_ sky130_fd_sc_hd__nand2_1
X_11856_ _01701_ _04874_ VGND VGND VPWR VPWR _01795_ sky130_fd_sc_hd__or2_1
XFILLER_0_157_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10807_ _00723_ _00744_ _00745_ VGND VGND VPWR VPWR _00746_ sky130_fd_sc_hd__a21oi_1
X_14575_ _04582_ _04586_ _04589_ VGND VGND VPWR VPWR _04591_ sky130_fd_sc_hd__or3_1
XFILLER_0_27_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17363_ net280 _02933_ VGND VGND VPWR VPWR _07658_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11787_ prev_error\[6\] _00242_ VGND VGND VPWR VPWR _01726_ sky130_fd_sc_hd__and2b_1
XFILLER_0_126_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19102_ net499 prev_error\[12\] VGND VGND VPWR VPWR _09539_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16314_ _06376_ _06503_ VGND VGND VPWR VPWR _06504_ sky130_fd_sc_hd__xor2_1
X_13526_ _03368_ _03383_ _03382_ VGND VGND VPWR VPWR _03485_ sky130_fd_sc_hd__o21a_1
X_10738_ _00673_ _00675_ _00477_ _00676_ VGND VGND VPWR VPWR _00677_ sky130_fd_sc_hd__a2bb2o_1
X_17294_ net299 _06801_ _06890_ net295 VGND VGND VPWR VPWR _07582_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19033_ net563 net92 VGND VGND VPWR VPWR _09492_ sky130_fd_sc_hd__and2_1
X_13457_ _03410_ _03414_ _03415_ VGND VGND VPWR VPWR _03416_ sky130_fd_sc_hd__o21ba_1
X_16245_ net272 _06404_ VGND VGND VPWR VPWR _06428_ sky130_fd_sc_hd__nand2_1
X_10669_ _00519_ _00517_ _00518_ VGND VGND VPWR VPWR _00608_ sky130_fd_sc_hd__and3_1
XFILLER_0_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_124_Right_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12408_ _02306_ _02345_ _02244_ _02346_ VGND VGND VPWR VPWR _02347_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13388_ _03330_ _03305_ _03329_ VGND VGND VPWR VPWR _03342_ sky130_fd_sc_hd__and3_1
X_16176_ _06351_ VGND VGND VPWR VPWR _06352_ sky130_fd_sc_hd__buf_6
X_12339_ _02269_ _02277_ _02275_ VGND VGND VPWR VPWR _02278_ sky130_fd_sc_hd__a21oi_1
X_15127_ _05104_ _05197_ VGND VGND VPWR VPWR _05198_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15058_ _05032_ _05121_ VGND VGND VPWR VPWR _05122_ sky130_fd_sc_hd__nand2_1
X_14009_ _03902_ _03958_ _03979_ VGND VGND VPWR VPWR _03981_ sky130_fd_sc_hd__or3b_1
X_18817_ _09255_ _09256_ VGND VGND VPWR VPWR _09257_ sky130_fd_sc_hd__nor2_2
X_18748_ _06141_ _09180_ VGND VGND VPWR VPWR _09181_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_144_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18679_ _09101_ _09104_ VGND VGND VPWR VPWR _09105_ sky130_fd_sc_hd__or2b_1
XFILLER_0_58_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout300 ki\[9\] VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_111_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout311 ki\[5\] VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout322 net325 VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__buf_2
XFILLER_0_10_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout333 net334 VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__buf_1
Xfanout344 net345 VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__buf_2
Xfanout355 net357 VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__clkbuf_2
Xfanout366 net369 VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__clkbuf_4
X_09817_ _05325_ VGND VGND VPWR VPWR _05336_ sky130_fd_sc_hd__clkbuf_4
Xfanout377 net378 VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__buf_2
Xfanout388 net389 VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__buf_2
Xfanout399 net403 VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__clkbuf_4
X_09748_ net3 net61 VGND VGND VPWR VPWR _04577_ sky130_fd_sc_hd__or2b_1
XFILLER_0_97_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09679_ net48 _03614_ _03647_ net273 VGND VGND VPWR VPWR _00046_ sky130_fd_sc_hd__a22o_1
X_11710_ _01640_ _01641_ VGND VGND VPWR VPWR _01649_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12690_ _02624_ _02610_ VGND VGND VPWR VPWR _02629_ sky130_fd_sc_hd__or2b_1
XFILLER_0_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11641_ _01503_ _01579_ VGND VGND VPWR VPWR _01580_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14360_ _04344_ _04347_ _04349_ VGND VGND VPWR VPWR _04354_ sky130_fd_sc_hd__or3_1
XFILLER_0_65_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11572_ net381 _00614_ VGND VGND VPWR VPWR _01511_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13311_ _03171_ _03262_ _03257_ _03261_ VGND VGND VPWR VPWR _03264_ sky130_fd_sc_hd__a211o_1
Xinput19 measurement[8] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_1
X_10523_ _00359_ _00461_ VGND VGND VPWR VPWR _00462_ sky130_fd_sc_hd__or2_2
X_14291_ _04018_ _04020_ VGND VGND VPWR VPWR _04278_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16030_ _08636_ _08669_ _06190_ VGND VGND VPWR VPWR _06191_ sky130_fd_sc_hd__o21a_1
X_13242_ _03189_ _03191_ _03194_ VGND VGND VPWR VPWR _03195_ sky130_fd_sc_hd__a21oi_1
X_10454_ _00379_ _00392_ VGND VGND VPWR VPWR _00393_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13173_ net202 _02915_ _03070_ VGND VGND VPWR VPWR _03125_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10385_ _00323_ VGND VGND VPWR VPWR _00324_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12124_ net208 _01861_ _01899_ VGND VGND VPWR VPWR _02063_ sky130_fd_sc_hd__a21oi_1
X_17981_ _08331_ _08335_ _08336_ VGND VGND VPWR VPWR _08337_ sky130_fd_sc_hd__o21a_1
X_12055_ net210 _01810_ _01991_ _01992_ VGND VGND VPWR VPWR _01994_ sky130_fd_sc_hd__o2bb2a_1
X_16932_ _07182_ VGND VGND VPWR VPWR _07183_ sky130_fd_sc_hd__clkbuf_4
X_11006_ _00943_ _00944_ VGND VGND VPWR VPWR _00945_ sky130_fd_sc_hd__nand2_1
X_16863_ _07105_ _07092_ _07104_ VGND VGND VPWR VPWR _07108_ sky130_fd_sc_hd__and3_1
X_18602_ _09013_ _09017_ _09019_ VGND VGND VPWR VPWR _09020_ sky130_fd_sc_hd__a21oi_1
X_15814_ _05297_ _05381_ _05953_ VGND VGND VPWR VPWR _05954_ sky130_fd_sc_hd__o21ba_1
X_16794_ _07029_ _07031_ VGND VGND VPWR VPWR _07032_ sky130_fd_sc_hd__or2b_1
XFILLER_0_87_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18533_ _08926_ _08927_ _08941_ _08943_ VGND VGND VPWR VPWR _08945_ sky130_fd_sc_hd__o211a_1
X_15745_ _05870_ _05873_ VGND VGND VPWR VPWR _05878_ sky130_fd_sc_hd__xor2_1
X_12957_ _02613_ _02311_ VGND VGND VPWR VPWR _02896_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11908_ net199 VGND VGND VPWR VPWR _01847_ sky130_fd_sc_hd__inv_2
X_18464_ _08739_ _08744_ net527 _08771_ _08868_ VGND VGND VPWR VPWR _08869_ sky130_fd_sc_hd__o2111ai_1
X_15676_ net469 net188 net183 net473 VGND VGND VPWR VPWR _05802_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12888_ _02825_ _02826_ VGND VGND VPWR VPWR _02827_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17415_ _07645_ _07649_ _07714_ VGND VGND VPWR VPWR _07715_ sky130_fd_sc_hd__a21bo_1
X_14627_ _04647_ _04513_ VGND VGND VPWR VPWR _04648_ sky130_fd_sc_hd__nor2_1
X_18395_ _06146_ _06148_ VGND VGND VPWR VPWR _08793_ sky130_fd_sc_hd__nand2_1
X_11839_ _01757_ _01754_ VGND VGND VPWR VPWR _01778_ sky130_fd_sc_hd__xor2_1
XFILLER_0_56_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17346_ net294 _06891_ VGND VGND VPWR VPWR _07639_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14558_ _04564_ _04571_ VGND VGND VPWR VPWR _04572_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13509_ net266 _01908_ _03467_ VGND VGND VPWR VPWR _03468_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17277_ net287 _07182_ VGND VGND VPWR VPWR _07563_ sky130_fd_sc_hd__nand2_1
X_14489_ net448 net143 VGND VGND VPWR VPWR _04496_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19016_ _09466_ _09470_ _09474_ _09475_ VGND VGND VPWR VPWR _09476_ sky130_fd_sc_hd__and4_1
XFILLER_0_12_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16228_ net514 VGND VGND VPWR VPWR _06409_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_113_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16159_ _01796_ _06272_ _06305_ VGND VGND VPWR VPWR _06333_ sky130_fd_sc_hd__and3b_2
XFILLER_0_140_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09602_ _03003_ _03014_ _03025_ _03036_ VGND VGND VPWR VPWR _03047_ sky130_fd_sc_hd__or4_1
XFILLER_0_79_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10170_ _09197_ _09208_ VGND VGND VPWR VPWR _09219_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout130 net132 VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_4
Xfanout141 net145 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__buf_2
Xfanout152 kd_2\[10\] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__buf_2
Xfanout163 net164 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_2
Xfanout174 kd_2\[6\] VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_2
Xfanout185 net186 VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_4
Xfanout196 net198 VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_2
X_13860_ _03680_ _03814_ VGND VGND VPWR VPWR _03826_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12811_ net207 _02640_ VGND VGND VPWR VPWR _02750_ sky130_fd_sc_hd__and2_1
X_13791_ _03753_ _03756_ VGND VGND VPWR VPWR _03757_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15530_ _05636_ _05638_ _05640_ VGND VGND VPWR VPWR _05641_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_57_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12742_ _02587_ _02588_ VGND VGND VPWR VPWR _02681_ sky130_fd_sc_hd__xor2_1
XFILLER_0_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12673_ _02509_ _02611_ VGND VGND VPWR VPWR _02612_ sky130_fd_sc_hd__and2_1
X_15461_ _05482_ _05484_ VGND VGND VPWR VPWR _05565_ sky130_fd_sc_hd__or2_1
X_17200_ _07464_ _07465_ _07476_ _07477_ VGND VGND VPWR VPWR _07478_ sky130_fd_sc_hd__nand4_1
X_14412_ net438 net142 net137 net443 VGND VGND VPWR VPWR _04411_ sky130_fd_sc_hd__a22oi_1
X_11624_ _01538_ _01548_ _01562_ VGND VGND VPWR VPWR _01563_ sky130_fd_sc_hd__and3_1
X_18180_ _08554_ _08555_ i_error\[2\] VGND VGND VPWR VPWR _08556_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15392_ _05399_ _05398_ VGND VGND VPWR VPWR _05489_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17131_ _07400_ _07401_ VGND VGND VPWR VPWR _07402_ sky130_fd_sc_hd__and2_1
X_14343_ _04331_ _04314_ _04333_ VGND VGND VPWR VPWR _04336_ sky130_fd_sc_hd__nand3_1
X_11555_ _01440_ _01482_ _01493_ VGND VGND VPWR VPWR _01494_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10506_ _04984_ _07327_ _00444_ VGND VGND VPWR VPWR _00445_ sky130_fd_sc_hd__a21oi_4
X_14274_ _04257_ _04259_ net420 net151 VGND VGND VPWR VPWR _04260_ sky130_fd_sc_hd__and4bb_1
X_17062_ _07321_ _07325_ VGND VGND VPWR VPWR _07326_ sky130_fd_sc_hd__xor2_1
X_11486_ net377 _00515_ _01424_ VGND VGND VPWR VPWR _01425_ sky130_fd_sc_hd__a21bo_1
X_13225_ _03089_ _03177_ VGND VGND VPWR VPWR _03178_ sky130_fd_sc_hd__or2_1
X_16013_ _06133_ _06171_ VGND VGND VPWR VPWR _06173_ sky130_fd_sc_hd__and2b_1
XFILLER_0_110_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10437_ _00235_ _00297_ VGND VGND VPWR VPWR _00376_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13156_ _03031_ _03033_ VGND VGND VPWR VPWR _03106_ sky130_fd_sc_hd__nor2_1
X_10368_ _00305_ _00306_ VGND VGND VPWR VPWR _00307_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12107_ _01768_ _02041_ VGND VGND VPWR VPWR _02046_ sky130_fd_sc_hd__or2b_1
X_13087_ net228 _02331_ _02896_ _03029_ VGND VGND VPWR VPWR _03030_ sky130_fd_sc_hd__a31o_1
X_17964_ net331 net314 _06992_ _07568_ VGND VGND VPWR VPWR _08319_ sky130_fd_sc_hd__nand4_2
X_10299_ _04225_ _04269_ _04192_ _04203_ VGND VGND VPWR VPWR _00238_ sky130_fd_sc_hd__o211ai_4
X_16915_ net285 _06803_ VGND VGND VPWR VPWR _07165_ sky130_fd_sc_hd__nand2_1
X_12038_ _01766_ _01976_ VGND VGND VPWR VPWR _01977_ sky130_fd_sc_hd__nand2_1
X_17895_ _08173_ _08182_ VGND VGND VPWR VPWR _08243_ sky130_fd_sc_hd__xor2_1
XFILLER_0_109_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16846_ net282 _06803_ _07088_ VGND VGND VPWR VPWR _07089_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16777_ _06954_ _07012_ VGND VGND VPWR VPWR _07013_ sky130_fd_sc_hd__nand2_1
X_13989_ _03955_ _03960_ _03915_ VGND VGND VPWR VPWR _03961_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18516_ _08819_ _08924_ _08925_ _08785_ VGND VGND VPWR VPWR _08926_ sky130_fd_sc_hd__o2bb2a_1
X_15728_ _05832_ _05836_ VGND VGND VPWR VPWR _05859_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18447_ _08848_ _08849_ VGND VGND VPWR VPWR _08850_ sky130_fd_sc_hd__or2_1
X_15659_ _05737_ _05780_ _05782_ VGND VGND VPWR VPWR _05783_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18378_ _08773_ _08576_ VGND VGND VPWR VPWR _08774_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17329_ net304 _06620_ VGND VGND VPWR VPWR _07620_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11340_ _01212_ _01278_ VGND VGND VPWR VPWR _01279_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11271_ _01135_ _01208_ VGND VGND VPWR VPWR _01210_ sky130_fd_sc_hd__or2_1
X_13010_ net261 _01806_ VGND VGND VPWR VPWR _02949_ sky130_fd_sc_hd__nand2_1
X_10222_ _09472_ _00160_ VGND VGND VPWR VPWR _00161_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_18_Left_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10153_ _07250_ _07580_ _07558_ VGND VGND VPWR VPWR _09032_ sky130_fd_sc_hd__a21oi_1
X_14961_ net453 net459 net158 net154 VGND VGND VPWR VPWR _05015_ sky130_fd_sc_hd__and4_1
XFILLER_0_55_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10084_ net356 net510 _06029_ VGND VGND VPWR VPWR _08273_ sky130_fd_sc_hd__and3_1
X_16700_ _06903_ _06878_ VGND VGND VPWR VPWR _06928_ sky130_fd_sc_hd__or2b_1
X_13912_ _02468_ _02568_ VGND VGND VPWR VPWR _03880_ sky130_fd_sc_hd__xnor2_1
X_17680_ _08003_ _08005_ VGND VGND VPWR VPWR _08006_ sky130_fd_sc_hd__xor2_1
X_14892_ net413 net417 net194 net190 VGND VGND VPWR VPWR _04939_ sky130_fd_sc_hd__and4_1
X_16631_ _06778_ _06780_ VGND VGND VPWR VPWR _06852_ sky130_fd_sc_hd__and2_1
X_13843_ _03786_ _03807_ _03808_ VGND VGND VPWR VPWR _03809_ sky130_fd_sc_hd__or3_1
XFILLER_0_69_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16562_ net293 _06410_ _06773_ _06775_ VGND VGND VPWR VPWR _06776_ sky130_fd_sc_hd__a31o_1
X_13774_ net240 _02934_ VGND VGND VPWR VPWR _03740_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10986_ _00841_ _00842_ _00843_ VGND VGND VPWR VPWR _00925_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_27_Left_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18301_ _06376_ _08661_ _08663_ VGND VGND VPWR VPWR _08689_ sky130_fd_sc_hd__o21ai_1
X_15513_ _05617_ _05619_ _05621_ VGND VGND VPWR VPWR _05623_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_128_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12725_ _02662_ _02663_ VGND VGND VPWR VPWR _02664_ sky130_fd_sc_hd__nor2_1
X_19281_ clknet_4_6_0_clock _00059_ VGND VGND VPWR VPWR kp\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16493_ _06697_ _06699_ VGND VGND VPWR VPWR _06701_ sky130_fd_sc_hd__xor2_2
XFILLER_0_127_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18232_ _08529_ _08534_ _08611_ _08612_ VGND VGND VPWR VPWR _08613_ sky130_fd_sc_hd__a31o_1
XFILLER_0_128_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15444_ _05530_ _05541_ VGND VGND VPWR VPWR _05547_ sky130_fd_sc_hd__nand2_1
X_12656_ _02592_ _02594_ VGND VGND VPWR VPWR _02595_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11607_ _01525_ _01545_ VGND VGND VPWR VPWR _01546_ sky130_fd_sc_hd__xnor2_1
X_18163_ _08496_ _08497_ VGND VGND VPWR VPWR _08538_ sky130_fd_sc_hd__nor2_1
X_12587_ _02475_ _02504_ VGND VGND VPWR VPWR _02526_ sky130_fd_sc_hd__xor2_1
X_15375_ net472 net476 net167 net162 VGND VGND VPWR VPWR _05471_ sky130_fd_sc_hd__and4_1
XFILLER_0_53_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17114_ _07274_ _07276_ VGND VGND VPWR VPWR _07384_ sky130_fd_sc_hd__xnor2_2
X_14326_ _03955_ _04316_ _03915_ VGND VGND VPWR VPWR _04317_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11538_ net362 _00812_ _00818_ net366 VGND VGND VPWR VPWR _01477_ sky130_fd_sc_hd__a22o_1
X_18094_ _08459_ _08458_ VGND VGND VPWR VPWR _08462_ sky130_fd_sc_hd__and2b_1
Xmax_cap105 _03600_ VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__buf_1
XFILLER_0_151_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17045_ _07303_ _07304_ _07306_ _07307_ VGND VGND VPWR VPWR _07308_ sky130_fd_sc_hd__nand4_1
X_14257_ _03991_ _04240_ VGND VGND VPWR VPWR _04241_ sky130_fd_sc_hd__nor2_1
X_11469_ _01312_ _01346_ VGND VGND VPWR VPWR _01408_ sky130_fd_sc_hd__xnor2_4
XPHY_EDGE_ROW_36_Left_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13208_ _03142_ _03160_ VGND VGND VPWR VPWR _03161_ sky130_fd_sc_hd__nor2_1
X_14188_ net412 net418 net130 net124 VGND VGND VPWR VPWR _04165_ sky130_fd_sc_hd__and4_1
XFILLER_0_110_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13139_ _02985_ _03086_ VGND VGND VPWR VPWR _03087_ sky130_fd_sc_hd__nand2_1
X_18996_ _09183_ _09453_ _09189_ VGND VGND VPWR VPWR _09454_ sky130_fd_sc_hd__a21boi_2
X_17947_ _08296_ net110 VGND VGND VPWR VPWR _08300_ sky130_fd_sc_hd__nor2_1
X_17878_ net326 _06992_ VGND VGND VPWR VPWR _08224_ sky130_fd_sc_hd__nand2_1
X_16829_ _06960_ _07069_ VGND VGND VPWR VPWR _07070_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09996_ net384 _05072_ _07294_ VGND VGND VPWR VPWR _07305_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10840_ net359 _00244_ VGND VGND VPWR VPWR _00779_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10771_ _00706_ _00709_ VGND VGND VPWR VPWR _00710_ sky130_fd_sc_hd__nand2_1
X_12510_ _02392_ _02448_ VGND VGND VPWR VPWR _02449_ sky130_fd_sc_hd__nor2_1
X_13490_ net232 _02914_ VGND VGND VPWR VPWR _03449_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12441_ net231 _01860_ VGND VGND VPWR VPWR _02380_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12372_ _02221_ VGND VGND VPWR VPWR _02311_ sky130_fd_sc_hd__inv_2
X_15160_ _05231_ _05233_ VGND VGND VPWR VPWR _05234_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14111_ _04081_ _04082_ VGND VGND VPWR VPWR _04083_ sky130_fd_sc_hd__nor2_1
X_11323_ _01256_ _01261_ VGND VGND VPWR VPWR _01262_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15091_ _05154_ _05155_ _05157_ VGND VGND VPWR VPWR _05158_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_120_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14042_ _04012_ _04013_ VGND VGND VPWR VPWR _04014_ sky130_fd_sc_hd__nand2_1
X_11254_ _01171_ _01191_ VGND VGND VPWR VPWR _01193_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_120_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10205_ _04357_ _09552_ _04478_ _04412_ VGND VGND VPWR VPWR _09558_ sky130_fd_sc_hd__a31o_4
X_18850_ _02149_ _02151_ _02148_ _01930_ VGND VGND VPWR VPWR _09293_ sky130_fd_sc_hd__a2bb2o_1
X_11185_ _01035_ _01036_ VGND VGND VPWR VPWR _01124_ sky130_fd_sc_hd__xnor2_2
X_17801_ _08109_ _08112_ _08138_ VGND VGND VPWR VPWR _08139_ sky130_fd_sc_hd__a21o_1
X_10136_ _06920_ VGND VGND VPWR VPWR _08845_ sky130_fd_sc_hd__inv_2
X_18781_ _09033_ _09200_ VGND VGND VPWR VPWR _09217_ sky130_fd_sc_hd__nor2_1
X_15993_ _01350_ _06143_ VGND VGND VPWR VPWR _06151_ sky130_fd_sc_hd__xor2_1
X_17732_ _08057_ _08058_ _08062_ VGND VGND VPWR VPWR _08063_ sky130_fd_sc_hd__and3_1
X_14944_ _04955_ _04996_ _04993_ VGND VGND VPWR VPWR _04997_ sky130_fd_sc_hd__a21oi_1
X_10067_ net568 VGND VGND VPWR VPWR _08086_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17663_ net315 _06802_ VGND VGND VPWR VPWR _07988_ sky130_fd_sc_hd__nand2_1
X_14875_ _04919_ _04916_ VGND VGND VPWR VPWR _04921_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16614_ _06828_ _06833_ VGND VGND VPWR VPWR _06834_ sky130_fd_sc_hd__nor2_1
X_13826_ net261 _02934_ VGND VGND VPWR VPWR _03792_ sky130_fd_sc_hd__nand2_2
XFILLER_0_58_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17594_ net301 _07095_ _07911_ _07908_ VGND VGND VPWR VPWR _07912_ sky130_fd_sc_hd__a31o_1
XFILLER_0_98_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19333_ clknet_4_2_0_clock _00034_ VGND VGND VPWR VPWR kd_2\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16545_ _06757_ _06365_ VGND VGND VPWR VPWR _06758_ sky130_fd_sc_hd__and2b_1
X_13757_ net260 net256 _02638_ _02745_ VGND VGND VPWR VPWR _03723_ sky130_fd_sc_hd__and4_1
X_10969_ _00804_ _00819_ _00817_ VGND VGND VPWR VPWR _00908_ sky130_fd_sc_hd__o21a_1
X_12708_ net211 _02332_ VGND VGND VPWR VPWR _02647_ sky130_fd_sc_hd__nand2_1
X_19264_ clknet_4_12_0_clock _00146_ VGND VGND VPWR VPWR prev_d_error\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16476_ _06675_ _06680_ _06681_ VGND VGND VPWR VPWR _06682_ sky130_fd_sc_hd__o21ai_1
X_13688_ _03650_ _03651_ _03652_ VGND VGND VPWR VPWR _03653_ sky130_fd_sc_hd__or3_2
XFILLER_0_122_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18215_ _08593_ _08594_ VGND VGND VPWR VPWR _08595_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15427_ _05505_ _05526_ _05447_ _05527_ VGND VGND VPWR VPWR _05528_ sky130_fd_sc_hd__a211o_1
X_12639_ net259 _01785_ _01798_ net254 VGND VGND VPWR VPWR _02578_ sky130_fd_sc_hd__a22oi_1
X_19195_ clknet_4_14_0_clock _00077_ VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18146_ _07153_ _08516_ _07047_ VGND VGND VPWR VPWR _08519_ sky130_fd_sc_hd__a21oi_1
X_15358_ _05439_ _05442_ _05451_ VGND VGND VPWR VPWR _05452_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_44_Left_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14309_ _04157_ _04156_ _04101_ _04097_ VGND VGND VPWR VPWR _04298_ sky130_fd_sc_hd__a211o_1
X_18077_ _07773_ _07777_ _08442_ VGND VGND VPWR VPWR _08443_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_151_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15289_ _05365_ _05373_ _05375_ VGND VGND VPWR VPWR _05376_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17028_ _07284_ _07288_ VGND VGND VPWR VPWR _07289_ sky130_fd_sc_hd__xor2_2
XFILLER_0_21_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09850_ net368 net365 VGND VGND VPWR VPWR _05699_ sky130_fd_sc_hd__or2_1
X_09781_ net68 net10 VGND VGND VPWR VPWR _04940_ sky130_fd_sc_hd__and2b_1
X_18979_ _09403_ _09434_ VGND VGND VPWR VPWR _09435_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_147_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_53_Left_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_138_Right_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_12_0_clock clknet_0_clock VGND VGND VPWR VPWR clknet_4_12_0_clock sky130_fd_sc_hd__clkbuf_8
XFILLER_0_118_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_62_Left_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09979_ _07096_ _07085_ VGND VGND VPWR VPWR _07118_ sky130_fd_sc_hd__and2b_1
X_12990_ prev_error\[0\] _00810_ VGND VGND VPWR VPWR _02929_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11941_ _01857_ _01862_ _01864_ VGND VGND VPWR VPWR _01880_ sky130_fd_sc_hd__o21ba_1
X_14660_ net470 net131 prev_d_error\[18\] VGND VGND VPWR VPWR _04684_ sky130_fd_sc_hd__a21oi_1
X_11872_ prev_error\[15\] _05171_ VGND VGND VPWR VPWR _01811_ sky130_fd_sc_hd__xor2_4
XFILLER_0_39_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13611_ _03565_ _03569_ VGND VGND VPWR VPWR _03570_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10823_ _00477_ _00676_ _00675_ VGND VGND VPWR VPWR _00762_ sky130_fd_sc_hd__a21o_1
X_14591_ _04606_ _04607_ VGND VGND VPWR VPWR _04608_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_105_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16330_ _06519_ _06520_ VGND VGND VPWR VPWR _06521_ sky130_fd_sc_hd__nand2_1
X_13542_ _03500_ _03492_ VGND VGND VPWR VPWR _03501_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10754_ _00684_ _00688_ _00692_ VGND VGND VPWR VPWR _00693_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16261_ _06427_ _06429_ _06444_ VGND VGND VPWR VPWR _06445_ sky130_fd_sc_hd__a21bo_1
X_13473_ _03094_ _03431_ VGND VGND VPWR VPWR _03432_ sky130_fd_sc_hd__xnor2_1
X_10685_ _00611_ _00622_ _00603_ VGND VGND VPWR VPWR _00624_ sky130_fd_sc_hd__o21a_1
X_18000_ _08355_ _08357_ VGND VGND VPWR VPWR _08358_ sky130_fd_sc_hd__and2b_1
XFILLER_0_125_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15212_ _05205_ _05290_ VGND VGND VPWR VPWR _05291_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12424_ net246 _01786_ VGND VGND VPWR VPWR _02363_ sky130_fd_sc_hd__nand2_1
X_16192_ _06368_ VGND VGND VPWR VPWR _06369_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15143_ net467 net153 net135 net485 VGND VGND VPWR VPWR _05216_ sky130_fd_sc_hd__a22oi_2
X_12355_ _02292_ _02293_ VGND VGND VPWR VPWR _02294_ sky130_fd_sc_hd__nor2_1
XFILLER_0_133_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11306_ _01198_ _01201_ _01200_ VGND VGND VPWR VPWR _01245_ sky130_fd_sc_hd__a21o_1
X_12286_ net203 VGND VGND VPWR VPWR _02225_ sky130_fd_sc_hd__inv_2
X_15074_ _05123_ _05135_ _05139_ VGND VGND VPWR VPWR _05140_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_121_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14025_ _03989_ _03991_ _03996_ VGND VGND VPWR VPWR _03997_ sky130_fd_sc_hd__o21ai_1
X_18902_ net101 _09349_ VGND VGND VPWR VPWR _09350_ sky130_fd_sc_hd__xor2_1
X_11237_ _01050_ _01048_ net402 _06062_ VGND VGND VPWR VPWR _01176_ sky130_fd_sc_hd__a2bb2o_1
X_18833_ _09272_ _09273_ VGND VGND VPWR VPWR _09275_ sky130_fd_sc_hd__nor2_1
X_11168_ _01106_ _01024_ VGND VGND VPWR VPWR _01107_ sky130_fd_sc_hd__nor2_1
X_10119_ _08636_ _08647_ VGND VGND VPWR VPWR _08658_ sky130_fd_sc_hd__nor2_1
X_18764_ _09040_ _09042_ _09034_ VGND VGND VPWR VPWR _09199_ sky130_fd_sc_hd__o21a_1
X_11099_ _00948_ _00950_ _00949_ VGND VGND VPWR VPWR _01038_ sky130_fd_sc_hd__a21o_1
X_15976_ _00358_ _01694_ _00356_ VGND VGND VPWR VPWR _06132_ sky130_fd_sc_hd__a21oi_2
X_17715_ _07959_ _07978_ _08043_ VGND VGND VPWR VPWR _08045_ sky130_fd_sc_hd__o21ba_1
X_14927_ _04975_ _04967_ _04972_ VGND VGND VPWR VPWR _04978_ sky130_fd_sc_hd__nand3_1
X_18695_ _06086_ _06088_ VGND VGND VPWR VPWR _09123_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17646_ _07879_ _07967_ _07968_ VGND VGND VPWR VPWR _07969_ sky130_fd_sc_hd__or3_4
X_14858_ _04899_ _04901_ VGND VGND VPWR VPWR _04902_ sky130_fd_sc_hd__or2b_1
XFILLER_0_133_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13809_ _03771_ _03766_ _03770_ VGND VGND VPWR VPWR _03775_ sky130_fd_sc_hd__nor3_1
XFILLER_0_19_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17577_ _07890_ _07892_ VGND VGND VPWR VPWR _07893_ sky130_fd_sc_hd__or2b_1
XFILLER_0_129_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14789_ _04813_ _04824_ _04825_ VGND VGND VPWR VPWR _04826_ sky130_fd_sc_hd__nand3_1
XFILLER_0_58_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19316_ clknet_4_1_0_clock _00017_ VGND VGND VPWR VPWR kd_1\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16528_ _06672_ _06703_ _06738_ VGND VGND VPWR VPWR _06739_ sky130_fd_sc_hd__o21a_1
XFILLER_0_133_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19247_ clknet_4_14_0_clock _00129_ VGND VGND VPWR VPWR i_error\[15\] sky130_fd_sc_hd__dfxtp_1
X_16459_ _06648_ _06662_ _06660_ VGND VGND VPWR VPWR _06663_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_155_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19178_ net501 _09029_ VGND VGND VPWR VPWR _09586_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18129_ _08479_ _08499_ _08480_ VGND VGND VPWR VPWR _08500_ sky130_fd_sc_hd__o21a_1
XFILLER_0_112_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09902_ _06238_ _06260_ VGND VGND VPWR VPWR _06271_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout504 net507 VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09833_ _04929_ _05017_ _05501_ VGND VGND VPWR VPWR _05512_ sky130_fd_sc_hd__nand3_4
XFILLER_0_67_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09764_ _04742_ VGND VGND VPWR VPWR _04753_ sky130_fd_sc_hd__inv_2
X_09695_ net57 _03881_ _03914_ net370 VGND VGND VPWR VPWR _00074_ sky130_fd_sc_hd__a22o_1
Xrebuffer20 net572 VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10470_ _00408_ VGND VGND VPWR VPWR _00409_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_115_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12140_ net208 _01854_ _02078_ VGND VGND VPWR VPWR _02079_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12071_ _01984_ _01986_ VGND VGND VPWR VPWR _02010_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11022_ net401 _05402_ VGND VGND VPWR VPWR _00961_ sky130_fd_sc_hd__nand2_2
X_15830_ _04466_ _05970_ VGND VGND VPWR VPWR _05971_ sky130_fd_sc_hd__and2_1
X_15761_ net480 net192 VGND VGND VPWR VPWR _05895_ sky130_fd_sc_hd__and2_1
X_12973_ _02910_ _02911_ VGND VGND VPWR VPWR _02912_ sky130_fd_sc_hd__and2_1
X_17500_ net310 _06889_ VGND VGND VPWR VPWR _07808_ sky130_fd_sc_hd__nand2_1
X_14712_ _04681_ _04719_ VGND VGND VPWR VPWR _04741_ sky130_fd_sc_hd__nand2_1
X_11924_ _01857_ _01862_ VGND VGND VPWR VPWR _01863_ sky130_fd_sc_hd__xor2_1
X_18480_ net531 _08870_ VGND VGND VPWR VPWR _08886_ sky130_fd_sc_hd__and2_1
X_15692_ _05769_ _05797_ _05817_ VGND VGND VPWR VPWR _05819_ sky130_fd_sc_hd__and3_1
X_17431_ _07693_ _07653_ _07730_ _07731_ VGND VGND VPWR VPWR _07732_ sky130_fd_sc_hd__a211o_1
X_14643_ _04644_ _04662_ _04663_ VGND VGND VPWR VPWR _04666_ sky130_fd_sc_hd__nand3_1
X_11855_ net230 _01779_ _01787_ net226 VGND VGND VPWR VPWR _01794_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_68_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17362_ _07653_ _07654_ _07548_ _07601_ VGND VGND VPWR VPWR _07656_ sky130_fd_sc_hd__a211oi_2
X_10806_ _00743_ _00724_ VGND VGND VPWR VPWR _00745_ sky130_fd_sc_hd__and2b_1
XFILLER_0_138_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14574_ _04582_ _04586_ _04589_ VGND VGND VPWR VPWR _04590_ sky130_fd_sc_hd__o21ai_1
X_11786_ _01724_ _00322_ VGND VGND VPWR VPWR _01725_ sky130_fd_sc_hd__or2_2
X_19101_ _09536_ _06007_ _09538_ net488 VGND VGND VPWR VPWR _00106_ sky130_fd_sc_hd__o211a_1
X_16313_ _06500_ _06501_ VGND VGND VPWR VPWR _06503_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13525_ _03480_ _03482_ _03483_ VGND VGND VPWR VPWR _03484_ sky130_fd_sc_hd__nand3_4
XFILLER_0_153_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17293_ net295 _06801_ VGND VGND VPWR VPWR _07581_ sky130_fd_sc_hd__nand2_1
X_10737_ _00674_ _07008_ VGND VGND VPWR VPWR _00676_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19032_ _09489_ _09490_ net492 VGND VGND VPWR VPWR _00078_ sky130_fd_sc_hd__o21a_1
X_16244_ _06347_ _06354_ _06356_ VGND VGND VPWR VPWR _06427_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_141_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13456_ _03386_ _03409_ net104 _03345_ VGND VGND VPWR VPWR _03415_ sky130_fd_sc_hd__a211oi_1
X_10668_ net347 _00325_ _00606_ VGND VGND VPWR VPWR _00607_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12407_ _02209_ _02243_ _02242_ VGND VGND VPWR VPWR _02346_ sky130_fd_sc_hd__a21o_1
XFILLER_0_112_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16175_ _01811_ _06350_ VGND VGND VPWR VPWR _06351_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_3_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13387_ _03340_ _03335_ VGND VGND VPWR VPWR _03341_ sky130_fd_sc_hd__xnor2_1
X_10599_ net393 _04874_ _04984_ net396 VGND VGND VPWR VPWR _00538_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15126_ _05190_ _05194_ _05196_ VGND VGND VPWR VPWR _05197_ sky130_fd_sc_hd__o21a_1
X_12338_ _02275_ _02276_ VGND VGND VPWR VPWR _02277_ sky130_fd_sc_hd__nor2_1
X_15057_ _05029_ _05031_ VGND VGND VPWR VPWR _05121_ sky130_fd_sc_hd__or2_1
X_12269_ _02067_ _02068_ _02070_ VGND VGND VPWR VPWR _02208_ sky130_fd_sc_hd__a21oi_1
X_14008_ _03902_ _03958_ _03979_ VGND VGND VPWR VPWR _03980_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_128_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18816_ _09254_ _04129_ VGND VGND VPWR VPWR _09256_ sky130_fd_sc_hd__and2b_1
X_15959_ _06036_ _06039_ VGND VGND VPWR VPWR _06113_ sky130_fd_sc_hd__xnor2_2
X_18747_ _09160_ _09159_ VGND VGND VPWR VPWR _09180_ sky130_fd_sc_hd__nor2b_2
X_18678_ _09102_ _09101_ _09103_ VGND VGND VPWR VPWR _09104_ sky130_fd_sc_hd__or3_4
XFILLER_0_53_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17629_ _07861_ _07863_ _07864_ VGND VGND VPWR VPWR _07950_ sky130_fd_sc_hd__nor3_1
XFILLER_0_148_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout301 ki\[8\] VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__clkbuf_4
Xfanout312 ki\[5\] VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__clkbuf_4
Xfanout323 net324 VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__clkbuf_4
Xfanout334 ki\[0\] VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__clkbuf_4
Xfanout345 kp\[15\] VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__clkbuf_2
Xfanout356 net357 VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__buf_4
Xfanout367 net369 VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__clkbuf_2
X_09816_ _05314_ VGND VGND VPWR VPWR _05325_ sky130_fd_sc_hd__clkbuf_4
Xfanout378 kp\[6\] VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__buf_2
Xfanout389 kp\[4\] VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__clkbuf_4
X_09747_ _04544_ _04555_ VGND VGND VPWR VPWR _04566_ sky130_fd_sc_hd__or2_1
X_09678_ net47 _03614_ _03647_ net277 VGND VGND VPWR VPWR _00045_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11640_ _01501_ _01502_ VGND VGND VPWR VPWR _01579_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11571_ _01286_ _01509_ VGND VGND VPWR VPWR _01510_ sky130_fd_sc_hd__xor2_1
XFILLER_0_119_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13310_ _03257_ _03261_ _03171_ _03262_ VGND VGND VPWR VPWR _03263_ sky130_fd_sc_hd__o211ai_2
X_10522_ _00425_ _00459_ _00460_ VGND VGND VPWR VPWR _00461_ sky130_fd_sc_hd__a21boi_1
X_14290_ _04274_ _04276_ VGND VGND VPWR VPWR _04277_ sky130_fd_sc_hd__and2_1
XFILLER_0_123_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13241_ _03192_ _03193_ VGND VGND VPWR VPWR _03194_ sky130_fd_sc_hd__xor2_1
X_10453_ _00389_ _00391_ _00387_ VGND VGND VPWR VPWR _00392_ sky130_fd_sc_hd__o21a_1
XFILLER_0_150_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13172_ _03108_ _03122_ VGND VGND VPWR VPWR _03123_ sky130_fd_sc_hd__or2_1
X_10384_ _00322_ VGND VGND VPWR VPWR _00323_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12123_ _02060_ _02061_ VGND VGND VPWR VPWR _02062_ sky130_fd_sc_hd__nand2_1
X_17980_ _08279_ _08280_ VGND VGND VPWR VPWR _08336_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12054_ _01991_ _01992_ net210 _01810_ VGND VGND VPWR VPWR _01993_ sky130_fd_sc_hd__and4bb_1
X_16931_ _07181_ VGND VGND VPWR VPWR _07182_ sky130_fd_sc_hd__buf_2
X_11005_ _00940_ _00939_ VGND VGND VPWR VPWR _00944_ sky130_fd_sc_hd__xnor2_2
X_16862_ _07092_ _07104_ _07105_ VGND VGND VPWR VPWR _07106_ sky130_fd_sc_hd__a21oi_1
X_15813_ _05465_ _05950_ _05951_ VGND VGND VPWR VPWR _05953_ sky130_fd_sc_hd__a21oi_1
X_18601_ _06168_ _09018_ VGND VGND VPWR VPWR _09019_ sky130_fd_sc_hd__and2_1
X_16793_ _07011_ _07028_ VGND VGND VPWR VPWR _07031_ sky130_fd_sc_hd__xor2_1
XFILLER_0_88_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18532_ _08938_ _08942_ _08937_ VGND VGND VPWR VPWR _08943_ sky130_fd_sc_hd__or3b_1
X_15744_ _05876_ VGND VGND VPWR VPWR _05877_ sky130_fd_sc_hd__inv_2
X_12956_ _02821_ _02894_ VGND VGND VPWR VPWR _02895_ sky130_fd_sc_hd__nor2_1
X_11907_ _01832_ _01843_ _01845_ VGND VGND VPWR VPWR _01846_ sky130_fd_sc_hd__o21a_1
X_18463_ _08830_ _08847_ _08865_ _08866_ _08863_ VGND VGND VPWR VPWR _08868_ sky130_fd_sc_hd__o32ai_2
X_15675_ net469 net473 net188 net183 VGND VGND VPWR VPWR _05801_ sky130_fd_sc_hd__and4_1
XFILLER_0_23_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12887_ _02824_ _02817_ _02821_ VGND VGND VPWR VPWR _02826_ sky130_fd_sc_hd__nor3_1
X_17414_ _07644_ _07643_ VGND VGND VPWR VPWR _07714_ sky130_fd_sc_hd__or2b_1
XFILLER_0_157_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14626_ _04508_ _04504_ VGND VGND VPWR VPWR _04647_ sky130_fd_sc_hd__and2b_1
X_11838_ _01775_ _01776_ VGND VGND VPWR VPWR _01777_ sky130_fd_sc_hd__nand2_2
X_18394_ _08560_ _08791_ VGND VGND VPWR VPWR _08792_ sky130_fd_sc_hd__xor2_2
XFILLER_0_157_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17345_ _07534_ _07543_ _07637_ VGND VGND VPWR VPWR _07638_ sky130_fd_sc_hd__a21oi_1
X_14557_ _04559_ _04561_ _04563_ VGND VGND VPWR VPWR _04571_ sky130_fd_sc_hd__or3_1
XFILLER_0_56_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11769_ _06634_ prev_error\[9\] VGND VGND VPWR VPWR _01708_ sky130_fd_sc_hd__or2b_1
XFILLER_0_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13508_ _03465_ _03466_ VGND VGND VPWR VPWR _03467_ sky130_fd_sc_hd__nor2_1
X_17276_ _07551_ _07556_ _07561_ VGND VGND VPWR VPWR _07562_ sky130_fd_sc_hd__o21a_1
X_14488_ net456 net139 VGND VGND VPWR VPWR _04495_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19015_ _09122_ _09132_ VGND VGND VPWR VPWR _09475_ sky130_fd_sc_hd__xnor2_2
X_16227_ _01742_ _06407_ VGND VGND VPWR VPWR _06408_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_2_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13439_ _03291_ _03290_ VGND VGND VPWR VPWR _03398_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16158_ _06312_ _06330_ VGND VGND VPWR VPWR _06332_ sky130_fd_sc_hd__nand2_1
X_15109_ _05175_ _05177_ VGND VGND VPWR VPWR _05178_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16089_ _06178_ _06193_ _06191_ VGND VGND VPWR VPWR _06256_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09601_ net29 net28 net30 VGND VGND VPWR VPWR _03036_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout120 net122 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__buf_2
Xfanout131 net132 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout142 net145 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_2
Xfanout153 net154 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__buf_2
Xfanout164 kd_2\[8\] VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_2
Xfanout175 kd_2\[5\] VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__buf_2
Xfanout186 kd_2\[3\] VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__buf_2
Xfanout197 net198 VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_4
X_12810_ _02225_ _02748_ _02635_ VGND VGND VPWR VPWR _02749_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13790_ _01763_ _03065_ _03755_ VGND VGND VPWR VPWR _03756_ sky130_fd_sc_hd__or3b_1
X_12741_ _02627_ _02679_ VGND VGND VPWR VPWR _02680_ sky130_fd_sc_hd__nand2_1
X_15460_ _05561_ _05563_ VGND VGND VPWR VPWR _05564_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12672_ net222 _01874_ _02508_ VGND VGND VPWR VPWR _02611_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14411_ net438 net443 net142 kd_2\[13\] VGND VGND VPWR VPWR _04410_ sky130_fd_sc_hd__and4_1
XFILLER_0_155_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11623_ _01553_ _01560_ _01561_ VGND VGND VPWR VPWR _01562_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15391_ _05476_ _05485_ _05487_ VGND VGND VPWR VPWR _05488_ sky130_fd_sc_hd__a21o_1
X_17130_ _07373_ _07394_ _07399_ VGND VGND VPWR VPWR _07401_ sky130_fd_sc_hd__or3_1
XFILLER_0_53_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14342_ _04331_ _04314_ _04333_ VGND VGND VPWR VPWR _04334_ sky130_fd_sc_hd__a21o_1
X_11554_ _01483_ _01491_ _01492_ VGND VGND VPWR VPWR _01493_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_108_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17061_ _07323_ _07324_ VGND VGND VPWR VPWR _07325_ sky130_fd_sc_hd__or2b_1
X_10505_ net396 _05512_ _05523_ _04984_ net392 VGND VGND VPWR VPWR _00444_ sky130_fd_sc_hd__a32oi_4
X_14273_ net425 net146 net141 net430 VGND VGND VPWR VPWR _04259_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_123_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11485_ net374 _00613_ VGND VGND VPWR VPWR _01424_ sky130_fd_sc_hd__nand2_1
X_16012_ _06169_ _06170_ VGND VGND VPWR VPWR _06171_ sky130_fd_sc_hd__nor2_1
X_13224_ _03084_ _03092_ _03176_ VGND VGND VPWR VPWR _03177_ sky130_fd_sc_hd__or3_2
X_10436_ _00369_ _00374_ VGND VGND VPWR VPWR _00375_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13155_ _03103_ _03104_ VGND VGND VPWR VPWR _03105_ sky130_fd_sc_hd__or2b_1
X_10367_ _07316_ _00301_ VGND VGND VPWR VPWR _00306_ sky130_fd_sc_hd__xor2_1
X_12106_ _02035_ _02044_ VGND VGND VPWR VPWR _02045_ sky130_fd_sc_hd__nor2_1
X_13086_ net224 _02408_ _03028_ VGND VGND VPWR VPWR _03029_ sky130_fd_sc_hd__and3_1
X_17963_ _08311_ _08313_ _08309_ VGND VGND VPWR VPWR _08318_ sky130_fd_sc_hd__o21a_1
XFILLER_0_109_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10298_ _00230_ _00236_ VGND VGND VPWR VPWR _00237_ sky130_fd_sc_hd__and2b_1
XFILLER_0_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16914_ _07097_ _07158_ _07163_ VGND VGND VPWR VPWR _07164_ sky130_fd_sc_hd__o21a_1
X_12037_ net246 _01764_ _01765_ VGND VGND VPWR VPWR _01976_ sky130_fd_sc_hd__a21bo_1
X_17894_ _08239_ _08241_ VGND VGND VPWR VPWR _08242_ sky130_fd_sc_hd__and2b_1
X_16845_ _06980_ _07087_ VGND VGND VPWR VPWR _07088_ sky130_fd_sc_hd__xnor2_1
X_16776_ _06951_ _06952_ VGND VGND VPWR VPWR _07012_ sky130_fd_sc_hd__or2_1
X_13988_ _03958_ _03959_ VGND VGND VPWR VPWR _03960_ sky130_fd_sc_hd__nor2_1
X_15727_ _05837_ _05857_ _05855_ VGND VGND VPWR VPWR _05858_ sky130_fd_sc_hd__o21ai_1
X_18515_ _06265_ _08787_ VGND VGND VPWR VPWR _08925_ sky130_fd_sc_hd__nor2_1
X_12939_ _02802_ _02877_ VGND VGND VPWR VPWR _02878_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15658_ _05774_ _05781_ VGND VGND VPWR VPWR _05782_ sky130_fd_sc_hd__nor2_1
X_18446_ _08542_ _08579_ _08584_ _08593_ _08831_ VGND VGND VPWR VPWR _08849_ sky130_fd_sc_hd__o311a_1
XFILLER_0_118_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14609_ _04603_ _04627_ VGND VGND VPWR VPWR _04628_ sky130_fd_sc_hd__and2b_1
X_18377_ i_error\[6\] _08574_ _08575_ VGND VGND VPWR VPWR _08773_ sky130_fd_sc_hd__and3_1
XFILLER_0_157_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15589_ _05703_ _05704_ _05705_ VGND VGND VPWR VPWR _05706_ sky130_fd_sc_hd__o21ba_1
X_17328_ _07527_ _07528_ VGND VGND VPWR VPWR _07619_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_44_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17259_ _07537_ _07542_ VGND VGND VPWR VPWR _07543_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11270_ _01135_ _01208_ VGND VGND VPWR VPWR _01209_ sky130_fd_sc_hd__and2_2
XFILLER_0_30_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10221_ _09483_ _00159_ _00157_ VGND VGND VPWR VPWR _00160_ sky130_fd_sc_hd__o21a_1
X_10152_ _08823_ _09010_ VGND VGND VPWR VPWR _09021_ sky130_fd_sc_hd__xnor2_1
X_14960_ net453 net158 net154 net459 VGND VGND VPWR VPWR _05014_ sky130_fd_sc_hd__a22oi_2
X_10083_ _08218_ _08251_ _08229_ VGND VGND VPWR VPWR _08262_ sky130_fd_sc_hd__o21ba_1
X_13911_ _02770_ _03876_ _03878_ VGND VGND VPWR VPWR _03879_ sky130_fd_sc_hd__a21o_1
X_14891_ _04934_ _04937_ VGND VGND VPWR VPWR _04938_ sky130_fd_sc_hd__nand2_1
X_16630_ _06849_ _06850_ VGND VGND VPWR VPWR _06851_ sky130_fd_sc_hd__or2b_1
X_13842_ _03758_ _03782_ VGND VGND VPWR VPWR _03808_ sky130_fd_sc_hd__xor2_2
XFILLER_0_69_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16561_ _06687_ _06774_ VGND VGND VPWR VPWR _06775_ sky130_fd_sc_hd__nor2_1
X_13773_ _01763_ _03731_ _03729_ VGND VGND VPWR VPWR _03739_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_85_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10985_ _00882_ _00923_ VGND VGND VPWR VPWR _00924_ sky130_fd_sc_hd__nor2_1
X_15512_ _05569_ _05620_ VGND VGND VPWR VPWR _05621_ sky130_fd_sc_hd__xnor2_1
X_18300_ _08678_ _08679_ _08687_ VGND VGND VPWR VPWR _08688_ sky130_fd_sc_hd__a21bo_1
X_12724_ _02632_ _02661_ VGND VGND VPWR VPWR _02663_ sky130_fd_sc_hd__and2_1
X_19280_ clknet_4_6_0_clock _00058_ VGND VGND VPWR VPWR kp\[10\] sky130_fd_sc_hd__dfxtp_2
X_16492_ _06649_ _06698_ _06548_ VGND VGND VPWR VPWR _06699_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18231_ i_error\[15\] _08528_ VGND VGND VPWR VPWR _08612_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15443_ _05469_ _05470_ _05544_ VGND VGND VPWR VPWR _05546_ sky130_fd_sc_hd__o21a_1
X_12655_ _02593_ _02485_ VGND VGND VPWR VPWR _02594_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11606_ _01540_ _01544_ VGND VGND VPWR VPWR _01545_ sky130_fd_sc_hd__nand2_1
X_18162_ i_error\[13\] _08535_ VGND VGND VPWR VPWR _08536_ sky130_fd_sc_hd__and2_1
X_15374_ _05463_ _05458_ _05461_ VGND VGND VPWR VPWR _05470_ sky130_fd_sc_hd__nor3_1
X_12586_ _02523_ _02524_ VGND VGND VPWR VPWR _02525_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17113_ _07352_ _07381_ VGND VGND VPWR VPWR _07383_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_136_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14325_ _04314_ _04315_ VGND VGND VPWR VPWR _04316_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11537_ _01469_ _01474_ _01475_ VGND VGND VPWR VPWR _01476_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_108_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18093_ _08458_ _08459_ VGND VGND VPWR VPWR _08461_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_151_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap106 _06553_ VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__buf_1
X_17044_ _07220_ _07222_ _07219_ VGND VGND VPWR VPWR _07307_ sky130_fd_sc_hd__a21o_1
X_14256_ net420 net146 _03989_ _03990_ VGND VGND VPWR VPWR _04240_ sky130_fd_sc_hd__o2bb2a_1
X_11468_ _01354_ _01406_ VGND VGND VPWR VPWR _01407_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13207_ _03156_ _03159_ VGND VGND VPWR VPWR _03160_ sky130_fd_sc_hd__and2_1
X_10419_ _00356_ _00357_ VGND VGND VPWR VPWR _00358_ sky130_fd_sc_hd__nor2_2
X_14187_ _04106_ _04109_ _04111_ VGND VGND VPWR VPWR _04164_ sky130_fd_sc_hd__or3_1
X_11399_ _01300_ _01309_ VGND VGND VPWR VPWR _01338_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13138_ _02986_ _03085_ VGND VGND VPWR VPWR _03086_ sky130_fd_sc_hd__nor2_1
X_18995_ _09136_ _09179_ VGND VGND VPWR VPWR _09453_ sky130_fd_sc_hd__and2b_1
X_13069_ _03007_ _03009_ VGND VGND VPWR VPWR _03010_ sky130_fd_sc_hd__xnor2_1
X_17946_ _08297_ _08296_ _08298_ VGND VGND VPWR VPWR _08299_ sky130_fd_sc_hd__nor3_1
XPHY_EDGE_ROW_119_Right_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17877_ _08158_ _08169_ _08222_ VGND VGND VPWR VPWR _08223_ sky130_fd_sc_hd__nand3_1
XFILLER_0_45_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16828_ net297 _06431_ _06434_ VGND VGND VPWR VPWR _07069_ sky130_fd_sc_hd__and3_2
XFILLER_0_45_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16759_ _06992_ VGND VGND VPWR VPWR _06993_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18429_ _08775_ _08781_ _08789_ _08822_ _08829_ VGND VGND VPWR VPWR _08830_ sky130_fd_sc_hd__o221a_1
XFILLER_0_119_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09995_ _07283_ VGND VGND VPWR VPWR _07294_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_86_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10770_ _00707_ _00708_ VGND VGND VPWR VPWR _00709_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12440_ _02288_ _02378_ VGND VGND VPWR VPWR _02379_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12371_ _02307_ _02309_ VGND VGND VPWR VPWR _02310_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14110_ _04075_ _04079_ VGND VGND VPWR VPWR _04082_ sky130_fd_sc_hd__nor2_1
X_11322_ _01258_ _01260_ VGND VGND VPWR VPWR _01261_ sky130_fd_sc_hd__nand2_1
X_15090_ _05049_ _05156_ VGND VGND VPWR VPWR _05157_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14041_ _03992_ _03994_ _04011_ VGND VGND VPWR VPWR _04013_ sky130_fd_sc_hd__or3_1
X_11253_ _01171_ _01191_ VGND VGND VPWR VPWR _01192_ sky130_fd_sc_hd__or2b_1
X_10204_ _04192_ _04313_ _04346_ _04379_ VGND VGND VPWR VPWR _09552_ sky130_fd_sc_hd__a211o_2
XFILLER_0_101_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11184_ _01104_ _01122_ VGND VGND VPWR VPWR _01123_ sky130_fd_sc_hd__nor2_1
X_17800_ _08106_ _08113_ VGND VGND VPWR VPWR _08138_ sky130_fd_sc_hd__and2_1
X_10135_ _07272_ _07349_ VGND VGND VPWR VPWR _08834_ sky130_fd_sc_hd__nor2_1
X_18780_ _09033_ _09200_ VGND VGND VPWR VPWR _09216_ sky130_fd_sc_hd__and2_1
X_15992_ _06146_ _06148_ VGND VGND VPWR VPWR _06149_ sky130_fd_sc_hd__or2_1
X_10066_ _07976_ _07998_ _08020_ VGND VGND VPWR VPWR _08075_ sky130_fd_sc_hd__a21o_1
X_14943_ _04993_ _04994_ VGND VGND VPWR VPWR _04996_ sky130_fd_sc_hd__nor2_1
X_17731_ net326 _06801_ _08060_ _08061_ VGND VGND VPWR VPWR _08062_ sky130_fd_sc_hd__a31o_1
X_14874_ _04916_ _04919_ VGND VGND VPWR VPWR _04920_ sky130_fd_sc_hd__and2b_1
XFILLER_0_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17662_ net313 _06890_ VGND VGND VPWR VPWR _07986_ sky130_fd_sc_hd__nand2_1
X_16613_ _06829_ _06831_ VGND VGND VPWR VPWR _06833_ sky130_fd_sc_hd__and2b_1
X_13825_ _03764_ _03790_ VGND VGND VPWR VPWR _03791_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17593_ _07908_ _07909_ VGND VGND VPWR VPWR _07911_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19332_ clknet_4_3_0_clock _00033_ VGND VGND VPWR VPWR kd_2\[5\] sky130_fd_sc_hd__dfxtp_1
X_16544_ _06754_ _06756_ VGND VGND VPWR VPWR _06757_ sky130_fd_sc_hd__xnor2_1
X_13756_ net263 _02408_ _03675_ VGND VGND VPWR VPWR _03722_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10968_ net337 _00811_ VGND VGND VPWR VPWR _00907_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12707_ net218 net215 _02224_ _02091_ VGND VGND VPWR VPWR _02646_ sky130_fd_sc_hd__nand4_1
X_19263_ clknet_4_3_0_clock _00145_ VGND VGND VPWR VPWR prev_d_error\[12\] sky130_fd_sc_hd__dfxtp_1
X_16475_ _06606_ _06607_ VGND VGND VPWR VPWR _06681_ sky130_fd_sc_hd__xor2_1
XFILLER_0_45_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13687_ _03633_ _03649_ VGND VGND VPWR VPWR _03652_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10899_ _00836_ _00837_ VGND VGND VPWR VPWR _00838_ sky130_fd_sc_hd__xor2_1
XFILLER_0_122_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15426_ _05442_ _05443_ _05445_ VGND VGND VPWR VPWR _05527_ sky130_fd_sc_hd__a21oi_1
X_18214_ i_error\[9\] _08591_ VGND VGND VPWR VPWR _08594_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12638_ net264 net111 VGND VGND VPWR VPWR _02577_ sky130_fd_sc_hd__nand2_1
X_19194_ clknet_4_12_0_clock _00076_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18145_ _08516_ _08517_ VGND VGND VPWR VPWR _08518_ sky130_fd_sc_hd__and2_2
XFILLER_0_136_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15357_ _05275_ _05450_ VGND VGND VPWR VPWR _05451_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12569_ _02380_ _02507_ VGND VGND VPWR VPWR _02508_ sky130_fd_sc_hd__xor2_1
XFILLER_0_81_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14308_ _04289_ _04294_ _04296_ VGND VGND VPWR VPWR _04297_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18076_ _07775_ _07776_ VGND VGND VPWR VPWR _08442_ sky130_fd_sc_hd__or2b_1
XFILLER_0_41_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15288_ _05372_ _05362_ _05370_ VGND VGND VPWR VPWR _05375_ sky130_fd_sc_hd__nand3_1
XFILLER_0_124_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17027_ _07285_ _07287_ VGND VGND VPWR VPWR _07288_ sky130_fd_sc_hd__xnor2_2
X_14239_ net448 net123 _04220_ VGND VGND VPWR VPWR _04221_ sky130_fd_sc_hd__and3_1
XFILLER_0_150_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09780_ net10 net68 VGND VGND VPWR VPWR _04929_ sky130_fd_sc_hd__or2b_2
XFILLER_0_147_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18978_ _09425_ _09433_ VGND VGND VPWR VPWR _09434_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_0_Left_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17929_ _08271_ _08269_ VGND VGND VPWR VPWR _08280_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09978_ _07085_ _07096_ VGND VGND VPWR VPWR _07107_ sky130_fd_sc_hd__and2b_1
X_11940_ _01868_ _01878_ VGND VGND VPWR VPWR _01879_ sky130_fd_sc_hd__and2b_1
X_11871_ _01799_ VGND VGND VPWR VPWR _01810_ sky130_fd_sc_hd__buf_2
XFILLER_0_79_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13610_ net237 _02915_ _03567_ _03568_ VGND VGND VPWR VPWR _03569_ sky130_fd_sc_hd__a31oi_1
X_10822_ _00720_ _00747_ VGND VGND VPWR VPWR _00761_ sky130_fd_sc_hd__xnor2_1
X_14590_ _03913_ _04605_ _04603_ VGND VGND VPWR VPWR _04607_ sky130_fd_sc_hd__nor3_1
XFILLER_0_39_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13541_ _03458_ _03462_ VGND VGND VPWR VPWR _03500_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10753_ _00689_ _00691_ VGND VGND VPWR VPWR _00692_ sky130_fd_sc_hd__and2b_1
XFILLER_0_137_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16260_ _06442_ _06443_ VGND VGND VPWR VPWR _06444_ sky130_fd_sc_hd__nand2_1
X_13472_ net251 _02222_ VGND VGND VPWR VPWR _03431_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10684_ _00603_ _00611_ _00622_ VGND VGND VPWR VPWR _00623_ sky130_fd_sc_hd__nor3_1
XFILLER_0_152_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15211_ _05286_ _05289_ VGND VGND VPWR VPWR _05290_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12423_ net250 net111 _01761_ VGND VGND VPWR VPWR _02362_ sky130_fd_sc_hd__a21oi_1
X_16191_ net303 _06324_ _06367_ VGND VGND VPWR VPWR _06368_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15142_ net484 net153 VGND VGND VPWR VPWR _05214_ sky130_fd_sc_hd__nand2_1
X_12354_ _02291_ _02284_ _02288_ VGND VGND VPWR VPWR _02293_ sky130_fd_sc_hd__nor3_1
XFILLER_0_106_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11305_ _01214_ _01243_ VGND VGND VPWR VPWR _01244_ sky130_fd_sc_hd__and2b_1
X_15073_ _05136_ _05137_ VGND VGND VPWR VPWR _05139_ sky130_fd_sc_hd__or2_1
X_12285_ _02223_ VGND VGND VPWR VPWR _02224_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14024_ _03994_ _03995_ VGND VGND VPWR VPWR _03996_ sky130_fd_sc_hd__nor2_1
X_18901_ _09345_ _09348_ VGND VGND VPWR VPWR _09349_ sky130_fd_sc_hd__xor2_1
X_11236_ _01050_ _01047_ _01048_ VGND VGND VPWR VPWR _01175_ sky130_fd_sc_hd__or3_1
XFILLER_0_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18832_ _09270_ _09271_ _04213_ VGND VGND VPWR VPWR _09273_ sky130_fd_sc_hd__a21oi_1
X_11167_ net351 _00815_ VGND VGND VPWR VPWR _01106_ sky130_fd_sc_hd__nand2_1
X_10118_ _08625_ _08614_ VGND VGND VPWR VPWR _08647_ sky130_fd_sc_hd__and2b_1
X_18763_ _09058_ _09196_ _09056_ VGND VGND VPWR VPWR _09198_ sky130_fd_sc_hd__o21ai_2
X_15975_ _00186_ _01696_ VGND VGND VPWR VPWR _06131_ sky130_fd_sc_hd__xor2_4
X_11098_ _01035_ _01036_ VGND VGND VPWR VPWR _01037_ sky130_fd_sc_hd__and2b_1
XFILLER_0_26_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17714_ _07959_ _07978_ _08043_ VGND VGND VPWR VPWR _08044_ sky130_fd_sc_hd__nor3b_2
X_10049_ _07866_ _07877_ VGND VGND VPWR VPWR _07888_ sky130_fd_sc_hd__nor2_1
X_14926_ _04908_ _04906_ VGND VGND VPWR VPWR _04977_ sky130_fd_sc_hd__xnor2_1
X_18694_ _09108_ _09121_ VGND VGND VPWR VPWR _09122_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_78_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17645_ _07876_ _07878_ _07839_ VGND VGND VPWR VPWR _07968_ sky130_fd_sc_hd__a21oi_1
X_14857_ _04821_ _04900_ VGND VGND VPWR VPWR _04901_ sky130_fd_sc_hd__xor2_1
XFILLER_0_26_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13808_ _03758_ _03773_ VGND VGND VPWR VPWR _03774_ sky130_fd_sc_hd__or2_1
X_14788_ _04812_ _04800_ _04810_ VGND VGND VPWR VPWR _04825_ sky130_fd_sc_hd__nand3_1
X_17576_ _07891_ _07842_ VGND VGND VPWR VPWR _07892_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19315_ clknet_4_1_0_clock _00016_ VGND VGND VPWR VPWR kd_1\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16527_ _06736_ _06737_ VGND VGND VPWR VPWR _06738_ sky130_fd_sc_hd__or2b_1
X_13739_ _03690_ _03703_ _03653_ _03704_ VGND VGND VPWR VPWR _03705_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19246_ clknet_4_12_0_clock _00128_ VGND VGND VPWR VPWR i_error\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16458_ _06660_ _06661_ VGND VGND VPWR VPWR _06662_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15409_ _05506_ _05507_ net437 net197 VGND VGND VPWR VPWR _05508_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_6_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19177_ net502 net439 net490 _09585_ VGND VGND VPWR VPWR _00143_ sky130_fd_sc_hd__o211a_1
X_16389_ _06584_ _06585_ VGND VGND VPWR VPWR _06586_ sky130_fd_sc_hd__nor2_1
X_18128_ _08465_ _08477_ VGND VGND VPWR VPWR _08499_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18059_ _08417_ _08419_ _08420_ _08421_ _08422_ VGND VGND VPWR VPWR _08423_ sky130_fd_sc_hd__a32o_1
XFILLER_0_41_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09901_ _06128_ _06249_ VGND VGND VPWR VPWR _06260_ sky130_fd_sc_hd__and2b_1
XFILLER_0_112_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7 _04654_ VGND VGND VPWR VPWR net562 sky130_fd_sc_hd__buf_6
Xfanout505 net506 VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__clkbuf_4
X_09832_ net69 net11 VGND VGND VPWR VPWR _05501_ sky130_fd_sc_hd__xor2_2
X_09763_ net65 net7 VGND VGND VPWR VPWR _04742_ sky130_fd_sc_hd__xnor2_1
X_09694_ net56 _03881_ _03914_ net558 VGND VGND VPWR VPWR _00073_ sky130_fd_sc_hd__a22o_1
Xrebuffer10 _08437_ VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__clkbuf_1
Xrebuffer21 _08754_ VGND VGND VPWR VPWR net528 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12070_ _01971_ _02008_ VGND VGND VPWR VPWR _02009_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11021_ _00932_ _00933_ _00934_ VGND VGND VPWR VPWR _00960_ sky130_fd_sc_hd__o21ai_2
X_15760_ _05874_ _05877_ _05878_ VGND VGND VPWR VPWR _05894_ sky130_fd_sc_hd__a21oi_1
X_12972_ _02893_ _02908_ _02909_ VGND VGND VPWR VPWR _02911_ sky130_fd_sc_hd__or3_1
X_11923_ net203 _01861_ VGND VGND VPWR VPWR _01862_ sky130_fd_sc_hd__nand2_1
X_14711_ _04738_ _04739_ VGND VGND VPWR VPWR _04740_ sky130_fd_sc_hd__and2_1
X_15691_ _05769_ _05797_ _05817_ VGND VGND VPWR VPWR _05818_ sky130_fd_sc_hd__a21o_1
XFILLER_0_157_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14642_ _04644_ _04662_ _04663_ VGND VGND VPWR VPWR _04664_ sky130_fd_sc_hd__a21o_1
X_17430_ _07711_ _07713_ _07729_ VGND VGND VPWR VPWR _07731_ sky130_fd_sc_hd__o21a_1
X_11854_ net230 net226 _01779_ _01787_ VGND VGND VPWR VPWR _01793_ sky130_fd_sc_hd__and4_1
XFILLER_0_68_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10805_ _00724_ _00743_ VGND VGND VPWR VPWR _00744_ sky130_fd_sc_hd__xnor2_4
X_14573_ _04388_ _04587_ VGND VGND VPWR VPWR _04589_ sky130_fd_sc_hd__nor2_1
X_17361_ _07548_ _07601_ _07653_ _07654_ VGND VGND VPWR VPWR _07655_ sky130_fd_sc_hd__o211a_2
X_11785_ prev_error\[5\] VGND VGND VPWR VPWR _01724_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19100_ net499 prev_error\[11\] VGND VGND VPWR VPWR _09538_ sky130_fd_sc_hd__or2_1
X_13524_ _03479_ _03472_ _03477_ VGND VGND VPWR VPWR _03483_ sky130_fd_sc_hd__or3_2
X_16312_ _06499_ _06490_ _06494_ VGND VGND VPWR VPWR _06501_ sky130_fd_sc_hd__nand3_1
X_17292_ _07504_ _07511_ VGND VGND VPWR VPWR _07579_ sky130_fd_sc_hd__nand2_1
X_10736_ net379 _06062_ _08735_ _00674_ VGND VGND VPWR VPWR _00675_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_126_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19031_ _09448_ _09485_ _09474_ VGND VGND VPWR VPWR _09490_ sky130_fd_sc_hd__a21oi_1
X_16243_ _06416_ _06424_ VGND VGND VPWR VPWR _06426_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_152_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13455_ _03411_ _03413_ VGND VGND VPWR VPWR _03414_ sky130_fd_sc_hd__xnor2_1
X_10667_ _00604_ _00605_ VGND VGND VPWR VPWR _00606_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12406_ _02306_ _02343_ _02344_ VGND VGND VPWR VPWR _02345_ sky130_fd_sc_hd__nor3_1
X_16174_ _06299_ _06343_ _06349_ VGND VGND VPWR VPWR _06350_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_152_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13386_ _01848_ _03220_ VGND VGND VPWR VPWR _03340_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10598_ net396 net392 _04874_ _04984_ VGND VGND VPWR VPWR _00537_ sky130_fd_sc_hd__nand4_1
X_15125_ _05097_ _05195_ VGND VGND VPWR VPWR _05196_ sky130_fd_sc_hd__and2_1
X_12337_ _02270_ _02274_ _02273_ VGND VGND VPWR VPWR _02276_ sky130_fd_sc_hd__nor3_1
XFILLER_0_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_81_Left_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15056_ _05113_ _05119_ VGND VGND VPWR VPWR _05120_ sky130_fd_sc_hd__nand2_1
X_12268_ _02206_ VGND VGND VPWR VPWR _02207_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14007_ _03936_ _03978_ VGND VGND VPWR VPWR _03979_ sky130_fd_sc_hd__or2_1
X_11219_ _01153_ _01156_ _01157_ VGND VGND VPWR VPWR _01158_ sky130_fd_sc_hd__o21a_1
X_12199_ _02123_ _02124_ _02137_ VGND VGND VPWR VPWR _02138_ sky130_fd_sc_hd__a21o_1
Xoutput90 net90 VGND VGND VPWR VPWR out_clocked[1] sky130_fd_sc_hd__buf_2
X_18815_ _03902_ _03907_ _09254_ VGND VGND VPWR VPWR _09255_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18746_ _09177_ _09178_ VGND VGND VPWR VPWR _09179_ sky130_fd_sc_hd__xnor2_2
X_15958_ _06050_ _06110_ _06111_ VGND VGND VPWR VPWR _06112_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14909_ _04796_ VGND VGND VPWR VPWR _04958_ sky130_fd_sc_hd__inv_2
X_18677_ net511 _09100_ _09095_ VGND VGND VPWR VPWR _09103_ sky130_fd_sc_hd__a21oi_1
X_15889_ _03876_ _06035_ VGND VGND VPWR VPWR _06036_ sky130_fd_sc_hd__and2_2
XPHY_EDGE_ROW_90_Left_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17628_ _07924_ _07948_ VGND VGND VPWR VPWR _07949_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17559_ _07872_ VGND VGND VPWR VPWR _07873_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19229_ clknet_4_5_0_clock _00111_ VGND VGND VPWR VPWR prev_error\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout302 net304 VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__clkbuf_4
Xfanout313 ki\[5\] VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout324 net325 VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__clkbuf_4
Xfanout335 kp\[18\] VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__buf_2
Xfanout346 net347 VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__buf_2
Xfanout357 kp\[12\] VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__clkbuf_4
X_09815_ _05292_ _05303_ VGND VGND VPWR VPWR _05314_ sky130_fd_sc_hd__and2_2
Xfanout368 net369 VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__clkbuf_4
Xfanout379 net380 VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09746_ net62 net4 VGND VGND VPWR VPWR _04555_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_129_Left_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09677_ net46 _03614_ _03647_ net280 VGND VGND VPWR VPWR _00044_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11570_ net385 _00515_ VGND VGND VPWR VPWR _01509_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10521_ _00427_ _00458_ VGND VGND VPWR VPWR _00460_ sky130_fd_sc_hd__or2b_1
XFILLER_0_134_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_138_Left_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13240_ net236 _02223_ VGND VGND VPWR VPWR _03193_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10452_ _00332_ _00390_ VGND VGND VPWR VPWR _00391_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_33_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13171_ _03119_ _03121_ VGND VGND VPWR VPWR _03122_ sky130_fd_sc_hd__and2b_1
XFILLER_0_0_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10383_ _04324_ _00321_ VGND VGND VPWR VPWR _00322_ sky130_fd_sc_hd__xor2_4
X_12122_ _02059_ _02053_ _02057_ VGND VGND VPWR VPWR _02061_ sky130_fd_sc_hd__nand3_1
XFILLER_0_20_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12053_ net218 _01930_ _01941_ VGND VGND VPWR VPWR _01992_ sky130_fd_sc_hd__and3_1
X_16930_ _02744_ _06276_ VGND VGND VPWR VPWR _07181_ sky130_fd_sc_hd__xor2_4
X_11004_ _00896_ _00942_ VGND VGND VPWR VPWR _00943_ sky130_fd_sc_hd__nor2_1
X_16861_ _06999_ _06988_ VGND VGND VPWR VPWR _07105_ sky130_fd_sc_hd__xor2_1
X_18600_ _09013_ _09017_ VGND VGND VPWR VPWR _09018_ sky130_fd_sc_hd__xor2_1
X_15812_ _05297_ _05381_ VGND VGND VPWR VPWR _05951_ sky130_fd_sc_hd__xnor2_1
X_16792_ _06972_ _06970_ VGND VGND VPWR VPWR _07029_ sky130_fd_sc_hd__xor2_1
X_18531_ _08927_ _08934_ _08926_ VGND VGND VPWR VPWR _08942_ sky130_fd_sc_hd__or3b_1
XFILLER_0_99_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15743_ net466 net483 net195 net179 VGND VGND VPWR VPWR _05876_ sky130_fd_sc_hd__and4_1
X_12955_ _02818_ _02820_ VGND VGND VPWR VPWR _02894_ sky130_fd_sc_hd__and2_1
X_11906_ _01825_ _01844_ VGND VGND VPWR VPWR _01845_ sky130_fd_sc_hd__nor2_1
X_18462_ _08854_ _08844_ _08864_ VGND VGND VPWR VPWR _08866_ sky130_fd_sc_hd__o21a_1
X_15674_ net478 net176 _05738_ _05739_ VGND VGND VPWR VPWR _05800_ sky130_fd_sc_hd__o2bb2a_1
X_12886_ _02817_ _02821_ _02824_ VGND VGND VPWR VPWR _02825_ sky130_fd_sc_hd__o21a_1
XFILLER_0_87_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17413_ _07709_ _07710_ _07694_ _07630_ VGND VGND VPWR VPWR _07713_ sky130_fd_sc_hd__o211a_1
X_14625_ _04644_ _04645_ VGND VGND VPWR VPWR _04646_ sky130_fd_sc_hd__nand2_1
X_11837_ _01768_ _01774_ VGND VGND VPWR VPWR _01776_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18393_ _08563_ _08562_ VGND VGND VPWR VPWR _08791_ sky130_fd_sc_hd__or2b_1
XFILLER_0_135_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14556_ _04567_ _04569_ VGND VGND VPWR VPWR _04570_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17344_ _07542_ _07537_ VGND VGND VPWR VPWR _07637_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11768_ _06194_ prev_error\[10\] VGND VGND VPWR VPWR _01707_ sky130_fd_sc_hd__and2b_1
XFILLER_0_16_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13507_ net258 _02222_ _02089_ net262 VGND VGND VPWR VPWR _03466_ sky130_fd_sc_hd__a22oi_1
X_10719_ _00565_ _00653_ _00657_ VGND VGND VPWR VPWR _00658_ sky130_fd_sc_hd__o21a_1
XFILLER_0_125_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14487_ _04483_ _04486_ _04493_ VGND VGND VPWR VPWR _04494_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17275_ _07557_ _07560_ VGND VGND VPWR VPWR _07561_ sky130_fd_sc_hd__or2b_1
X_11699_ _01637_ VGND VGND VPWR VPWR _01638_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19014_ _09471_ _09473_ VGND VGND VPWR VPWR _09474_ sky130_fd_sc_hd__xor2_2
X_13438_ net224 _02914_ _03396_ VGND VGND VPWR VPWR _03397_ sky130_fd_sc_hd__and3_1
X_16226_ _06298_ _06297_ _01738_ _07008_ VGND VGND VPWR VPWR _06407_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_153_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer1 _09136_ VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__buf_1
XFILLER_0_140_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16157_ _06312_ _06330_ VGND VGND VPWR VPWR _06331_ sky130_fd_sc_hd__or2_1
X_13369_ _03319_ _03313_ _03318_ VGND VGND VPWR VPWR _03322_ sky130_fd_sc_hd__or3_2
XFILLER_0_51_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15108_ _05075_ _05176_ VGND VGND VPWR VPWR _05177_ sky130_fd_sc_hd__nor2_1
X_16088_ _06251_ _06254_ VGND VGND VPWR VPWR _06255_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15039_ _05000_ _05099_ VGND VGND VPWR VPWR _05101_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09600_ net25 net24 net27 net26 VGND VGND VPWR VPWR _03025_ sky130_fd_sc_hd__or4_1
XFILLER_0_155_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18729_ _09158_ _09155_ _09156_ VGND VGND VPWR VPWR _09160_ sky130_fd_sc_hd__and3_1
XFILLER_0_149_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout121 net122 VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_4
Xfanout132 kd_2\[15\] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__buf_4
Xfanout143 net144 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__buf_2
Xfanout154 kd_2\[10\] VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_2
Xfanout165 net169 VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__buf_2
Xfanout176 net178 VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__buf_2
Xfanout187 net188 VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__buf_2
Xfanout198 kd_2\[0\] VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__buf_2
X_09729_ net75 net17 VGND VGND VPWR VPWR _04368_ sky130_fd_sc_hd__or2b_1
XFILLER_0_97_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12740_ _02625_ _02626_ VGND VGND VPWR VPWR _02679_ sky130_fd_sc_hd__or2_1
XFILLER_0_139_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12671_ _02608_ _02609_ VGND VGND VPWR VPWR _02610_ sky130_fd_sc_hd__xor2_1
XFILLER_0_49_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14410_ _04385_ _04408_ VGND VGND VPWR VPWR _04409_ sky130_fd_sc_hd__or2b_1
XFILLER_0_154_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11622_ _01555_ _01559_ VGND VGND VPWR VPWR _01561_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15390_ _05416_ _05486_ VGND VGND VPWR VPWR _05487_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_146_Left_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14341_ _04242_ _04332_ VGND VGND VPWR VPWR _04333_ sky130_fd_sc_hd__or2_1
X_11553_ _01484_ _01486_ _01490_ VGND VGND VPWR VPWR _01492_ sky130_fd_sc_hd__nand3_1
XFILLER_0_37_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10504_ net539 _07327_ VGND VGND VPWR VPWR _00443_ sky130_fd_sc_hd__nand2_1
X_17060_ net334 _01755_ _06314_ _07322_ VGND VGND VPWR VPWR _07324_ sky130_fd_sc_hd__a31o_1
X_14272_ net425 net430 net146 net141 VGND VGND VPWR VPWR _04257_ sky130_fd_sc_hd__and4_1
X_11484_ net370 _00815_ VGND VGND VPWR VPWR _01423_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16011_ _00358_ _01694_ VGND VGND VPWR VPWR _06170_ sky130_fd_sc_hd__xor2_4
XFILLER_0_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13223_ _03139_ _03175_ _03173_ VGND VGND VPWR VPWR _03176_ sky130_fd_sc_hd__a21oi_1
X_10435_ _00372_ _00373_ VGND VGND VPWR VPWR _00374_ sky130_fd_sc_hd__or2b_1
XFILLER_0_60_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13154_ _03097_ _03098_ VGND VGND VPWR VPWR _03104_ sky130_fd_sc_hd__xor2_1
XFILLER_0_103_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10366_ _07338_ _00304_ VGND VGND VPWR VPWR _00305_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12105_ _02011_ _02043_ _01978_ VGND VGND VPWR VPWR _02044_ sky130_fd_sc_hd__a21oi_1
X_13085_ _03027_ _02896_ VGND VGND VPWR VPWR _03028_ sky130_fd_sc_hd__xnor2_1
X_17962_ _08309_ _08314_ _08315_ VGND VGND VPWR VPWR _08316_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_155_Left_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10297_ _00232_ _00235_ VGND VGND VPWR VPWR _00236_ sky130_fd_sc_hd__or2_1
X_16913_ _07159_ _07161_ VGND VGND VPWR VPWR _07163_ sky130_fd_sc_hd__or2b_1
X_12036_ _01973_ _01974_ VGND VGND VPWR VPWR _01975_ sky130_fd_sc_hd__or2_1
X_17893_ _08231_ _08228_ VGND VGND VPWR VPWR _08241_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16844_ net285 _06723_ VGND VGND VPWR VPWR _07087_ sky130_fd_sc_hd__nand2_1
X_16775_ _06917_ _07010_ VGND VGND VPWR VPWR _07011_ sky130_fd_sc_hd__nand2_1
X_13987_ _03905_ _03957_ VGND VGND VPWR VPWR _03959_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18514_ _06265_ _08817_ VGND VGND VPWR VPWR _08924_ sky130_fd_sc_hd__or2_1
X_15726_ _05855_ _05856_ VGND VGND VPWR VPWR _05857_ sky130_fd_sc_hd__nand2_1
X_12938_ net240 _01853_ _02801_ VGND VGND VPWR VPWR _02877_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18445_ _08594_ VGND VGND VPWR VPWR _08848_ sky130_fd_sc_hd__inv_2
X_15657_ _05737_ _05780_ VGND VGND VPWR VPWR _05781_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12869_ _02793_ _02806_ _02709_ _02807_ VGND VGND VPWR VPWR _02808_ sky130_fd_sc_hd__a211o_1
XFILLER_0_87_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14608_ _04596_ _04602_ VGND VGND VPWR VPWR _04627_ sky130_fd_sc_hd__nand2_1
X_18376_ _08544_ _08571_ VGND VGND VPWR VPWR _08772_ sky130_fd_sc_hd__or2_1
X_15588_ net455 net457 net191 net187 VGND VGND VPWR VPWR _05705_ sky130_fd_sc_hd__and4_1
XFILLER_0_7_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17327_ net302 _06724_ _07541_ _07539_ VGND VGND VPWR VPWR _07618_ sky130_fd_sc_hd__a31o_1
X_14539_ _04549_ _04550_ VGND VGND VPWR VPWR _04551_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17258_ _07538_ _07541_ VGND VGND VPWR VPWR _07542_ sky130_fd_sc_hd__xor2_2
XFILLER_0_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16209_ net286 _06336_ _06311_ net289 VGND VGND VPWR VPWR _06388_ sky130_fd_sc_hd__a22oi_1
X_17189_ net323 net319 _06408_ _06401_ VGND VGND VPWR VPWR _07466_ sky130_fd_sc_hd__nand4_1
XFILLER_0_141_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10220_ _00157_ _00158_ VGND VGND VPWR VPWR _00159_ sky130_fd_sc_hd__nand2_1
X_10151_ _08988_ _08999_ VGND VGND VPWR VPWR _09010_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10082_ _08229_ _08240_ VGND VGND VPWR VPWR _08251_ sky130_fd_sc_hd__or2_1
X_13910_ _02673_ _03877_ VGND VGND VPWR VPWR _03878_ sky130_fd_sc_hd__nand2_1
X_14890_ _04935_ _04936_ VGND VGND VPWR VPWR _04937_ sky130_fd_sc_hd__xnor2_1
X_13841_ _03788_ _03806_ VGND VGND VPWR VPWR _03807_ sky130_fd_sc_hd__or2b_1
X_16560_ net300 _06345_ VGND VGND VPWR VPWR _06774_ sky130_fd_sc_hd__nand2_1
X_13772_ _03721_ _03737_ VGND VGND VPWR VPWR _03738_ sky130_fd_sc_hd__or2_2
X_10984_ _00878_ _00881_ VGND VGND VPWR VPWR _00923_ sky130_fd_sc_hd__and2_1
X_15511_ _05571_ _05570_ VGND VGND VPWR VPWR _05620_ sky130_fd_sc_hd__nor2_1
X_12723_ _02632_ _02661_ VGND VGND VPWR VPWR _02662_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16491_ _06677_ _06679_ VGND VGND VPWR VPWR _06698_ sky130_fd_sc_hd__xor2_1
X_18230_ _08536_ _08608_ _08609_ _08610_ VGND VGND VPWR VPWR _08611_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_155_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12654_ net234 _01835_ VGND VGND VPWR VPWR _02593_ sky130_fd_sc_hd__nand2_1
X_15442_ _05539_ _05542_ _05461_ _05543_ VGND VGND VPWR VPWR _05544_ sky130_fd_sc_hd__a211o_2
XFILLER_0_38_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11605_ _01540_ _01542_ _01543_ VGND VGND VPWR VPWR _01544_ sky130_fd_sc_hd__nand3_2
XFILLER_0_143_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18161_ _07046_ _08520_ VGND VGND VPWR VPWR _08535_ sky130_fd_sc_hd__xor2_4
X_12585_ _02522_ _02517_ VGND VGND VPWR VPWR _02524_ sky130_fd_sc_hd__and2b_1
X_15373_ _05464_ VGND VGND VPWR VPWR _05469_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17112_ _07365_ _07380_ VGND VGND VPWR VPWR _07381_ sky130_fd_sc_hd__xnor2_2
X_14324_ _04307_ _04309_ _04312_ VGND VGND VPWR VPWR _04315_ sky130_fd_sc_hd__or3_1
XFILLER_0_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11536_ _01467_ _01468_ VGND VGND VPWR VPWR _01475_ sky130_fd_sc_hd__nand2_1
X_18092_ _07383_ _07384_ VGND VGND VPWR VPWR _08459_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_25_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14255_ _04237_ _04234_ VGND VGND VPWR VPWR _04239_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap107 _03539_ VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_2
X_17043_ _07219_ _07220_ _07222_ VGND VGND VPWR VPWR _07306_ sky130_fd_sc_hd__nand3_1
X_11467_ _01401_ _01405_ VGND VGND VPWR VPWR _01406_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13206_ _03156_ _03157_ _03158_ VGND VGND VPWR VPWR _03159_ sky130_fd_sc_hd__nand3_1
X_10418_ _00354_ _00355_ VGND VGND VPWR VPWR _00357_ sky130_fd_sc_hd__and2_1
X_14186_ _04129_ _04139_ _04141_ VGND VGND VPWR VPWR _04163_ sky130_fd_sc_hd__o21bai_2
X_11398_ _01331_ _01335_ _01268_ _01336_ VGND VGND VPWR VPWR _01337_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_29_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13137_ _03081_ _03084_ VGND VGND VPWR VPWR _03085_ sky130_fd_sc_hd__nor2_1
X_10349_ _00286_ _00287_ VGND VGND VPWR VPWR _00288_ sky130_fd_sc_hd__nand2_1
X_18994_ _09058_ _09196_ VGND VGND VPWR VPWR _09452_ sky130_fd_sc_hd__xnor2_1
X_13068_ _03008_ _02889_ VGND VGND VPWR VPWR _03009_ sky130_fd_sc_hd__xnor2_1
X_17945_ _08293_ _08294_ _08283_ _08292_ VGND VGND VPWR VPWR _08298_ sky130_fd_sc_hd__a211oi_1
X_12019_ net205 _01817_ VGND VGND VPWR VPWR _01958_ sky130_fd_sc_hd__nand2_1
X_17876_ _08220_ _08221_ VGND VGND VPWR VPWR _08222_ sky130_fd_sc_hd__nor2_1
X_16827_ _07067_ _06962_ VGND VGND VPWR VPWR _07068_ sky130_fd_sc_hd__xor2_1
XFILLER_0_45_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16758_ _06991_ VGND VGND VPWR VPWR _06992_ sky130_fd_sc_hd__buf_4
XFILLER_0_49_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15709_ net469 net473 net191 net187 VGND VGND VPWR VPWR _05838_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16689_ _06910_ _06913_ VGND VGND VPWR VPWR _06916_ sky130_fd_sc_hd__xor2_1
X_18428_ _08826_ _08828_ VGND VGND VPWR VPWR _08829_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18359_ _08596_ _08600_ _08607_ VGND VGND VPWR VPWR _08753_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09994_ _05534_ _05490_ _05061_ VGND VGND VPWR VPWR _07283_ sky130_fd_sc_hd__and3b_1
XFILLER_0_99_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12370_ _02308_ _02232_ VGND VGND VPWR VPWR _02309_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11321_ net402 _06172_ _01258_ _01259_ VGND VGND VPWR VPWR _01260_ sky130_fd_sc_hd__nand4_2
X_14040_ _03992_ _03994_ _04011_ VGND VGND VPWR VPWR _04012_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_133_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11252_ _01059_ _01172_ _01186_ _01190_ VGND VGND VPWR VPWR _01191_ sky130_fd_sc_hd__a31o_2
X_10203_ net341 _06634_ _09540_ VGND VGND VPWR VPWR _09546_ sky130_fd_sc_hd__and3_1
X_11183_ _01104_ _01105_ _01121_ VGND VGND VPWR VPWR _01122_ sky130_fd_sc_hd__nor3b_1
X_10134_ _08801_ _08812_ VGND VGND VPWR VPWR _08823_ sky130_fd_sc_hd__and2_1
X_15991_ _06147_ _01675_ VGND VGND VPWR VPWR _06148_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_100_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17730_ _08054_ _08059_ VGND VGND VPWR VPWR _08061_ sky130_fd_sc_hd__nor2_1
X_10065_ _07811_ _07822_ _08053_ VGND VGND VPWR VPWR _08064_ sky130_fd_sc_hd__a21o_1
X_14942_ _04992_ _04987_ _04990_ VGND VGND VPWR VPWR _04994_ sky130_fd_sc_hd__and3_1
X_17661_ _07889_ _07983_ _07982_ VGND VGND VPWR VPWR _07985_ sky130_fd_sc_hd__a21o_1
X_14873_ _04832_ _04917_ VGND VGND VPWR VPWR _04919_ sky130_fd_sc_hd__nor2_1
X_16612_ _06734_ _06792_ _06793_ _06830_ VGND VGND VPWR VPWR _06831_ sky130_fd_sc_hd__o31ai_2
X_13824_ net263 _02641_ _03763_ VGND VGND VPWR VPWR _03790_ sky130_fd_sc_hd__a21oi_1
X_17592_ _07808_ _07907_ VGND VGND VPWR VPWR _07909_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19331_ clknet_4_3_0_clock _00032_ VGND VGND VPWR VPWR kd_2\[4\] sky130_fd_sc_hd__dfxtp_1
X_16543_ _06366_ _06320_ _06676_ VGND VGND VPWR VPWR _06756_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_156_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13755_ _03687_ _03720_ VGND VGND VPWR VPWR _03721_ sky130_fd_sc_hd__or2_1
X_10967_ net346 _00615_ _00905_ VGND VGND VPWR VPWR _00906_ sky130_fd_sc_hd__and3_1
X_12706_ _02547_ _02635_ _02644_ VGND VGND VPWR VPWR _02645_ sky130_fd_sc_hd__o21bai_2
X_19262_ clknet_4_11_0_clock _00144_ VGND VGND VPWR VPWR prev_d_error\[11\] sky130_fd_sc_hd__dfxtp_1
X_16474_ _06677_ _06679_ VGND VGND VPWR VPWR _06680_ sky130_fd_sc_hd__and2_1
X_13686_ _03622_ _03627_ VGND VGND VPWR VPWR _03651_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10898_ net397 _04764_ _05369_ VGND VGND VPWR VPWR _00837_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18213_ i_error\[9\] _08591_ VGND VGND VPWR VPWR _08593_ sky130_fd_sc_hd__nand2_1
X_15425_ _05521_ _05522_ _05525_ VGND VGND VPWR VPWR _05526_ sky130_fd_sc_hd__or3_2
XFILLER_0_54_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12637_ _02490_ _02503_ VGND VGND VPWR VPWR _02576_ sky130_fd_sc_hd__xnor2_2
X_19193_ _09550_ _09438_ _09594_ net491 VGND VGND VPWR VPWR _00151_ sky130_fd_sc_hd__o211a_1
X_18144_ _08507_ _08514_ VGND VGND VPWR VPWR _08517_ sky130_fd_sc_hd__or2_1
X_12568_ net227 _01852_ VGND VGND VPWR VPWR _02507_ sky130_fd_sc_hd__nand2_1
X_15356_ net419 net198 _05274_ VGND VGND VPWR VPWR _05450_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_152_Right_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14307_ _04101_ _04295_ VGND VGND VPWR VPWR _04296_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11519_ _01456_ _01457_ VGND VGND VPWR VPWR _01458_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18075_ _07974_ _08440_ VGND VGND VPWR VPWR _08441_ sky130_fd_sc_hd__nand2_1
X_12499_ _02271_ _02272_ VGND VGND VPWR VPWR _02438_ sky130_fd_sc_hd__nor2_1
X_15287_ _05373_ VGND VGND VPWR VPWR _05374_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17026_ _07119_ _07286_ VGND VGND VPWR VPWR _07287_ sky130_fd_sc_hd__xor2_2
X_14238_ _04218_ _04219_ VGND VGND VPWR VPWR _04220_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14169_ _04127_ _04143_ VGND VGND VPWR VPWR _04144_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18977_ _09426_ _09432_ VGND VGND VPWR VPWR _09433_ sky130_fd_sc_hd__xnor2_1
X_17928_ _08277_ _08278_ VGND VGND VPWR VPWR _08279_ sky130_fd_sc_hd__xor2_1
X_17859_ _08083_ _08098_ VGND VGND VPWR VPWR _08203_ sky130_fd_sc_hd__xor2_2
XFILLER_0_89_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_101_Left_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09977_ net348 _05193_ _06821_ _06832_ VGND VGND VPWR VPWR _07096_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_110_Left_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_6_0_clock clknet_0_clock VGND VGND VPWR VPWR clknet_4_6_0_clock sky130_fd_sc_hd__clkbuf_8
X_11870_ net208 _01808_ VGND VGND VPWR VPWR _01809_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10821_ _00752_ _00750_ VGND VGND VPWR VPWR _00760_ sky130_fd_sc_hd__xor2_1
XFILLER_0_138_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13540_ _03496_ _03498_ VGND VGND VPWR VPWR _03499_ sky130_fd_sc_hd__or2b_1
X_10752_ _00607_ _00690_ VGND VGND VPWR VPWR _00691_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13471_ _03428_ _03429_ VGND VGND VPWR VPWR _03430_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10683_ _00619_ _00621_ VGND VGND VPWR VPWR _00622_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12422_ _02294_ _02297_ VGND VGND VPWR VPWR _02361_ sky130_fd_sc_hd__xnor2_1
X_15210_ _05268_ _05280_ _05288_ VGND VGND VPWR VPWR _05289_ sky130_fd_sc_hd__o21a_1
X_16190_ net309 ki\[7\] _06366_ VGND VGND VPWR VPWR _06367_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_51_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12353_ _02284_ _02288_ _02291_ VGND VGND VPWR VPWR _02292_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15141_ _05208_ _05210_ _05212_ VGND VGND VPWR VPWR _05213_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11304_ _01229_ _01241_ _01242_ VGND VGND VPWR VPWR _01243_ sky130_fd_sc_hd__o21bai_2
X_15072_ _05034_ _05033_ _05018_ VGND VGND VPWR VPWR _05137_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12284_ _02222_ VGND VGND VPWR VPWR _02223_ sky130_fd_sc_hd__clkbuf_4
X_14023_ net407 net156 _03992_ _03993_ VGND VGND VPWR VPWR _03995_ sky130_fd_sc_hd__o2bb2a_1
X_18900_ _08890_ _09347_ _08964_ VGND VGND VPWR VPWR _09348_ sky130_fd_sc_hd__mux2_2
X_11235_ _01141_ _01173_ VGND VGND VPWR VPWR _01174_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_121_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18831_ _04213_ _09270_ _09271_ VGND VGND VPWR VPWR _09272_ sky130_fd_sc_hd__and3_1
X_11166_ _01013_ _01103_ _01081_ _01102_ VGND VGND VPWR VPWR _01105_ sky130_fd_sc_hd__o211a_1
X_10117_ _08614_ _08625_ VGND VGND VPWR VPWR _08636_ sky130_fd_sc_hd__and2b_1
X_18762_ _09070_ _09194_ _09195_ VGND VGND VPWR VPWR _09196_ sky130_fd_sc_hd__a21oi_4
X_15974_ _06127_ _06129_ VGND VGND VPWR VPWR _06130_ sky130_fd_sc_hd__nor2_1
X_11097_ _01015_ _01014_ VGND VGND VPWR VPWR _01036_ sky130_fd_sc_hd__xnor2_2
X_17713_ _08036_ _08040_ _08041_ VGND VGND VPWR VPWR _08043_ sky130_fd_sc_hd__a21bo_1
X_10048_ net364 _05171_ _04885_ net368 VGND VGND VPWR VPWR _07877_ sky130_fd_sc_hd__a22oi_1
X_14925_ _04967_ _04972_ _04975_ VGND VGND VPWR VPWR _04976_ sky130_fd_sc_hd__a21o_1
X_18693_ _09117_ _09116_ VGND VGND VPWR VPWR _09121_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17644_ _07961_ _07966_ VGND VGND VPWR VPWR _07967_ sky130_fd_sc_hd__and2b_1
X_14856_ net461 net143 _04702_ _04822_ VGND VGND VPWR VPWR _04900_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13807_ net243 _02934_ _03757_ VGND VGND VPWR VPWR _03773_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17575_ net328 _06435_ VGND VGND VPWR VPWR _07891_ sky130_fd_sc_hd__nand2_1
X_14787_ _04818_ _04823_ VGND VGND VPWR VPWR _04824_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11999_ _01936_ _01937_ VGND VGND VPWR VPWR _01938_ sky130_fd_sc_hd__or2_1
X_19314_ clknet_4_1_0_clock _00015_ VGND VGND VPWR VPWR kd_1\[6\] sky130_fd_sc_hd__dfxtp_1
X_16526_ _06672_ _06703_ VGND VGND VPWR VPWR _06737_ sky130_fd_sc_hd__xor2_1
X_13738_ _03650_ _03652_ _03651_ VGND VGND VPWR VPWR _03704_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19245_ clknet_4_14_0_clock _00127_ VGND VGND VPWR VPWR i_error\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16457_ _06659_ _06653_ _06658_ VGND VGND VPWR VPWR _06661_ sky130_fd_sc_hd__nor3_1
X_13669_ _03582_ _03584_ VGND VGND VPWR VPWR _03632_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15408_ net441 net193 net189 net446 VGND VGND VPWR VPWR _05507_ sky130_fd_sc_hd__a22oi_1
X_19176_ net502 _09036_ VGND VGND VPWR VPWR _09585_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16388_ _06549_ _06583_ _06582_ VGND VGND VPWR VPWR _06585_ sky130_fd_sc_hd__and3_1
XFILLER_0_143_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18127_ _08496_ _08497_ _08478_ _08481_ VGND VGND VPWR VPWR _08498_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15339_ _05429_ _05430_ VGND VGND VPWR VPWR _05431_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18058_ _08302_ _08308_ VGND VGND VPWR VPWR _08422_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09900_ _05391_ _05952_ _06117_ VGND VGND VPWR VPWR _06249_ sky130_fd_sc_hd__or3b_1
XFILLER_0_10_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17009_ _07253_ _07257_ _07259_ VGND VGND VPWR VPWR _07268_ sky130_fd_sc_hd__or3_1
XFILLER_0_111_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout506 net507 VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__buf_2
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09831_ net406 net389 VGND VGND VPWR VPWR _05490_ sky130_fd_sc_hd__or2_1
X_09762_ net64 net6 VGND VGND VPWR VPWR _04731_ sky130_fd_sc_hd__and2b_2
X_09693_ net55 _03881_ _03914_ net378 VGND VGND VPWR VPWR _00072_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer11 _08549_ VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__clkbuf_1
Xrebuffer22 net528 VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11020_ _00957_ _00958_ VGND VGND VPWR VPWR _00959_ sky130_fd_sc_hd__and2_2
XFILLER_0_99_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12971_ _02893_ _02908_ _02909_ VGND VGND VPWR VPWR _02910_ sky130_fd_sc_hd__o21ai_1
X_14710_ _04736_ _04737_ _04728_ _04733_ VGND VGND VPWR VPWR _04739_ sky130_fd_sc_hd__a211o_1
X_11922_ _01860_ VGND VGND VPWR VPWR _01861_ sky130_fd_sc_hd__buf_2
X_15690_ _05752_ _05799_ _05811_ _05813_ _05816_ VGND VGND VPWR VPWR _05817_ sky130_fd_sc_hd__a32o_1
X_14641_ _04442_ _04461_ VGND VGND VPWR VPWR _04663_ sky130_fd_sc_hd__xnor2_1
X_11853_ _01788_ _01791_ VGND VGND VPWR VPWR _01792_ sky130_fd_sc_hd__xor2_1
X_17360_ _07632_ _07633_ _07652_ VGND VGND VPWR VPWR _07654_ sky130_fd_sc_hd__o21ai_1
X_10804_ _00725_ _00741_ _00742_ VGND VGND VPWR VPWR _00743_ sky130_fd_sc_hd__a21boi_4
X_14572_ net448 net135 _04386_ _04387_ VGND VGND VPWR VPWR _04587_ sky130_fd_sc_hd__o2bb2a_1
X_11784_ _01712_ _01713_ _01721_ _01722_ VGND VGND VPWR VPWR _01723_ sky130_fd_sc_hd__a31o_2
XFILLER_0_95_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16311_ _06490_ _06494_ _06499_ VGND VGND VPWR VPWR _06500_ sky130_fd_sc_hd__a21o_1
X_13523_ _03441_ _03481_ VGND VGND VPWR VPWR _03482_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17291_ _07505_ _07510_ VGND VGND VPWR VPWR _07578_ sky130_fd_sc_hd__nand2_1
X_10735_ net383 VGND VGND VPWR VPWR _00674_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19030_ net563 net91 VGND VGND VPWR VPWR _09489_ sky130_fd_sc_hd__and2_1
X_16242_ _06417_ _06423_ VGND VGND VPWR VPWR _06424_ sky130_fd_sc_hd__xor2_1
XFILLER_0_153_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13454_ _03225_ _03412_ VGND VGND VPWR VPWR _03413_ sky130_fd_sc_hd__or2_1
X_10666_ net351 _00245_ _00503_ VGND VGND VPWR VPWR _00605_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12405_ _02206_ _02305_ _02279_ _02304_ VGND VGND VPWR VPWR _02344_ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13385_ _03270_ _03338_ VGND VGND VPWR VPWR _03339_ sky130_fd_sc_hd__nor2_1
X_16173_ prev_error\[14\] net509 _05369_ VGND VGND VPWR VPWR _06349_ sky130_fd_sc_hd__and3_1
X_10597_ _00438_ _00445_ VGND VGND VPWR VPWR _00536_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_23_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15124_ _05093_ _05087_ _05096_ VGND VGND VPWR VPWR _05195_ sky130_fd_sc_hd__nand3_1
X_12336_ _02270_ _02273_ _02274_ VGND VGND VPWR VPWR _02275_ sky130_fd_sc_hd__o21a_1
XFILLER_0_105_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12267_ _02203_ _02205_ VGND VGND VPWR VPWR _02206_ sky130_fd_sc_hd__nor2_2
X_15055_ _05117_ _05118_ VGND VGND VPWR VPWR _05119_ sky130_fd_sc_hd__xnor2_1
X_14006_ _03930_ _03935_ VGND VGND VPWR VPWR _03978_ sky130_fd_sc_hd__nor2_1
X_11218_ _01090_ _01093_ VGND VGND VPWR VPWR _01157_ sky130_fd_sc_hd__xor2_1
X_12198_ _02126_ _02136_ VGND VGND VPWR VPWR _02137_ sky130_fd_sc_hd__xnor2_1
Xoutput80 net80 VGND VGND VPWR VPWR out_clocked[0] sky130_fd_sc_hd__buf_2
XFILLER_0_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput91 net91 VGND VGND VPWR VPWR out_clocked[2] sky130_fd_sc_hd__buf_2
X_18814_ _04138_ _09253_ VGND VGND VPWR VPWR _09254_ sky130_fd_sc_hd__xor2_1
X_11149_ net358 _00410_ VGND VGND VPWR VPWR _01088_ sky130_fd_sc_hd__nand2_1
X_18745_ _06099_ _09088_ _09091_ _09092_ _06145_ VGND VGND VPWR VPWR _09178_ sky130_fd_sc_hd__a32o_1
X_15957_ _06043_ _06045_ VGND VGND VPWR VPWR _06111_ sky130_fd_sc_hd__xnor2_1
X_14908_ _04813_ _04825_ _04824_ VGND VGND VPWR VPWR _04957_ sky130_fd_sc_hd__a21o_1
X_18676_ _06152_ VGND VGND VPWR VPWR _09102_ sky130_fd_sc_hd__inv_2
X_15888_ _03875_ _02873_ _03873_ VGND VGND VPWR VPWR _06035_ sky130_fd_sc_hd__nand3_1
XFILLER_0_144_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17627_ _07940_ _07947_ VGND VGND VPWR VPWR _07948_ sky130_fd_sc_hd__xnor2_2
X_14839_ _04858_ _04880_ VGND VGND VPWR VPWR _04881_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_53_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17558_ _07868_ _07869_ _07871_ VGND VGND VPWR VPWR _07872_ sky130_fd_sc_hd__or3_4
XFILLER_0_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16509_ _06273_ _02087_ _06287_ VGND VGND VPWR VPWR _06718_ sky130_fd_sc_hd__nand3_2
XFILLER_0_85_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17489_ _07768_ _07795_ VGND VGND VPWR VPWR _07796_ sky130_fd_sc_hd__xor2_2
X_19228_ clknet_4_5_0_clock _00110_ VGND VGND VPWR VPWR prev_error\[15\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_143_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19159_ net501 net482 net490 _09574_ VGND VGND VPWR VPWR _00134_ sky130_fd_sc_hd__o211a_1
XFILLER_0_143_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout303 net304 VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__buf_2
Xfanout314 ki\[4\] VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__clkbuf_4
Xfanout325 ki\[2\] VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__buf_2
Xfanout336 kp\[18\] VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__clkbuf_2
Xfanout347 kp\[14\] VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__buf_2
X_09814_ _05281_ _04731_ _04181_ _04709_ VGND VGND VPWR VPWR _05303_ sky130_fd_sc_hd__o211ai_4
Xfanout358 kp\[11\] VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__clkbuf_4
Xfanout369 kp\[9\] VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__clkbuf_4
X_09745_ net4 net62 VGND VGND VPWR VPWR _04544_ sky130_fd_sc_hd__and2b_1
XFILLER_0_97_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09676_ net45 _03614_ _03647_ net281 VGND VGND VPWR VPWR _00043_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10520_ _00427_ _00458_ VGND VGND VPWR VPWR _00459_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_91_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10451_ _00334_ _00333_ VGND VGND VPWR VPWR _00390_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13170_ _03108_ _03120_ VGND VGND VPWR VPWR _03121_ sky130_fd_sc_hd__nor2_1
X_10382_ _04280_ _00238_ _04335_ _04445_ VGND VGND VPWR VPWR _00321_ sky130_fd_sc_hd__a31o_1
XFILLER_0_60_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12121_ _02053_ _02057_ _02059_ VGND VGND VPWR VPWR _02060_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12052_ net218 _01930_ _01941_ VGND VGND VPWR VPWR _01991_ sky130_fd_sc_hd__a21oi_1
X_11003_ _00895_ _00893_ VGND VGND VPWR VPWR _00942_ sky130_fd_sc_hd__and2b_1
X_16860_ _07101_ _07103_ VGND VGND VPWR VPWR _07104_ sky130_fd_sc_hd__nand2_1
X_15811_ _05467_ _05949_ VGND VGND VPWR VPWR _05950_ sky130_fd_sc_hd__or2_1
X_16791_ _07013_ _07027_ _07025_ VGND VGND VPWR VPWR _07028_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18530_ _08931_ _08932_ _08940_ VGND VGND VPWR VPWR _08941_ sky130_fd_sc_hd__a21o_1
X_15742_ net466 net195 net179 net483 VGND VGND VPWR VPWR _05874_ sky130_fd_sc_hd__a22o_1
X_12954_ _02884_ _02891_ _02892_ VGND VGND VPWR VPWR _02893_ sky130_fd_sc_hd__a21oi_2
X_11905_ _01783_ _01823_ VGND VGND VPWR VPWR _01844_ sky130_fd_sc_hd__nor2_1
X_18461_ _08854_ _08863_ _08864_ VGND VGND VPWR VPWR _08865_ sky130_fd_sc_hd__or3b_1
X_15673_ _05749_ _05751_ VGND VGND VPWR VPWR _05799_ sky130_fd_sc_hd__or2_1
X_12885_ _02822_ _02823_ VGND VGND VPWR VPWR _02824_ sky130_fd_sc_hd__xnor2_1
X_17412_ _07694_ _07630_ _07709_ _07710_ VGND VGND VPWR VPWR _07711_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_157_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14624_ _04590_ _04640_ _04642_ VGND VGND VPWR VPWR _04645_ sky130_fd_sc_hd__nand3_1
X_11836_ _01768_ _01774_ VGND VGND VPWR VPWR _01775_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18392_ _08785_ _08788_ _08781_ _08775_ VGND VGND VPWR VPWR _08789_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17343_ _07588_ _07595_ _07634_ VGND VGND VPWR VPWR _07636_ sky130_fd_sc_hd__a21o_1
X_14555_ _04567_ _04568_ net409 net186 VGND VGND VPWR VPWR _04569_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11767_ prev_error\[12\] _06051_ VGND VGND VPWR VPWR _01706_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_55_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13506_ net262 net258 _02222_ _02089_ VGND VGND VPWR VPWR _03465_ sky130_fd_sc_hd__and4_1
XFILLER_0_15_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17274_ _07551_ _07556_ _07559_ VGND VGND VPWR VPWR _07560_ sky130_fd_sc_hd__o21a_1
X_10718_ _00654_ _00656_ VGND VGND VPWR VPWR _00657_ sky130_fd_sc_hd__or2b_1
XFILLER_0_126_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14486_ _04487_ _04492_ VGND VGND VPWR VPWR _04493_ sky130_fd_sc_hd__xnor2_1
X_11698_ net399 _00815_ VGND VGND VPWR VPWR _01637_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19013_ _09122_ _09132_ VGND VGND VPWR VPWR _09473_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16225_ net280 _06346_ VGND VGND VPWR VPWR _06406_ sky130_fd_sc_hd__nand2_1
X_13437_ _03394_ _03395_ VGND VGND VPWR VPWR _03396_ sky130_fd_sc_hd__nor2_1
Xrebuffer2 _01688_ VGND VGND VPWR VPWR net569 sky130_fd_sc_hd__buf_6
X_10649_ _00582_ _00587_ VGND VGND VPWR VPWR _00588_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16156_ _06327_ _06329_ VGND VGND VPWR VPWR _06330_ sky130_fd_sc_hd__nand2_1
X_13368_ _03284_ _03282_ VGND VGND VPWR VPWR _03321_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_23_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15107_ net414 net197 net193 net419 VGND VGND VPWR VPWR _05176_ sky130_fd_sc_hd__a22oi_1
X_12319_ net246 net111 VGND VGND VPWR VPWR _02258_ sky130_fd_sc_hd__nand2_1
X_16087_ net345 _05512_ _05523_ _06252_ _06253_ VGND VGND VPWR VPWR _06254_ sky130_fd_sc_hd__a41o_1
X_13299_ _03201_ _03214_ VGND VGND VPWR VPWR _03252_ sky130_fd_sc_hd__nand2_1
X_15038_ _05000_ _05099_ VGND VGND VPWR VPWR _05100_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16989_ _07210_ _07244_ _07245_ VGND VGND VPWR VPWR _07246_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_79_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18728_ _09155_ _09156_ _09158_ VGND VGND VPWR VPWR _09159_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18659_ _09080_ _09081_ _09074_ VGND VGND VPWR VPWR _09083_ sky130_fd_sc_hd__a21o_1
XFILLER_0_148_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout122 kd_2\[17\] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_4
Xfanout133 net135 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_4
Xfanout144 net145 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_4
Xfanout155 net156 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_4
Xfanout166 net168 VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__buf_2
Xfanout177 net178 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__buf_2
Xfanout188 kd_2\[2\] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__buf_2
Xfanout199 kd_1\[18\] VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09728_ net17 net75 VGND VGND VPWR VPWR _04357_ sky130_fd_sc_hd__nand2b_2
X_09659_ _03603_ net487 VGND VGND VPWR VPWR _03636_ sky130_fd_sc_hd__and2b_1
X_12670_ _02511_ _02515_ VGND VGND VPWR VPWR _02609_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11621_ _01555_ _01559_ VGND VGND VPWR VPWR _01560_ sky130_fd_sc_hd__xor2_1
XFILLER_0_108_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14340_ _04239_ _04241_ VGND VGND VPWR VPWR _04332_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11552_ _01484_ _01486_ _01490_ VGND VGND VPWR VPWR _01491_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10503_ net401 _00438_ _00441_ VGND VGND VPWR VPWR _00442_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14271_ _04230_ _04254_ _03986_ _04255_ VGND VGND VPWR VPWR _04256_ sky130_fd_sc_hd__a211oi_2
X_11483_ net377 _00613_ VGND VGND VPWR VPWR _01422_ sky130_fd_sc_hd__nand2_1
X_16010_ _06166_ _06168_ VGND VGND VPWR VPWR _06169_ sky130_fd_sc_hd__and2_1
X_10434_ _00368_ _00361_ VGND VGND VPWR VPWR _00373_ sky130_fd_sc_hd__xnor2_2
X_13222_ _03173_ _03174_ VGND VGND VPWR VPWR _03175_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10365_ _00301_ _00303_ VGND VGND VPWR VPWR _00304_ sky130_fd_sc_hd__and2_1
X_13153_ net236 _02223_ _03100_ _03101_ VGND VGND VPWR VPWR _03103_ sky130_fd_sc_hd__a31oi_2
X_12104_ _02039_ _02042_ VGND VGND VPWR VPWR _02043_ sky130_fd_sc_hd__xnor2_1
X_13084_ net228 _02330_ VGND VGND VPWR VPWR _03027_ sky130_fd_sc_hd__nand2_1
X_17961_ _08220_ _08221_ VGND VGND VPWR VPWR _08315_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10296_ net350 _06645_ _00234_ VGND VGND VPWR VPWR _00235_ sky130_fd_sc_hd__and3_1
X_16912_ _07097_ _07158_ _07160_ VGND VGND VPWR VPWR _07161_ sky130_fd_sc_hd__o21a_1
X_12035_ net259 net254 _01759_ VGND VGND VPWR VPWR _01974_ sky130_fd_sc_hd__nand3_1
X_17892_ _08237_ _08238_ VGND VGND VPWR VPWR _08239_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16843_ _06398_ _06993_ VGND VGND VPWR VPWR _07086_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16774_ _06915_ _06916_ VGND VGND VPWR VPWR _07010_ sky130_fd_sc_hd__nand2_1
X_13986_ _03905_ _03957_ VGND VGND VPWR VPWR _03958_ sky130_fd_sc_hd__nor2_1
X_18513_ _08775_ _08918_ _08920_ _08921_ VGND VGND VPWR VPWR _08923_ sky130_fd_sc_hd__a211o_1
X_15725_ _05854_ _05846_ _05851_ VGND VGND VPWR VPWR _05856_ sky130_fd_sc_hd__nand3_1
XFILLER_0_125_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12937_ _02835_ _02864_ _02863_ VGND VGND VPWR VPWR _02876_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18444_ _08844_ _08846_ VGND VGND VPWR VPWR _08847_ sky130_fd_sc_hd__nand2_1
X_15656_ _05772_ _05779_ VGND VGND VPWR VPWR _05780_ sky130_fd_sc_hd__or2b_1
X_12868_ _02696_ _02708_ _02707_ VGND VGND VPWR VPWR _02807_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_146_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14607_ _04623_ _04625_ VGND VGND VPWR VPWR _04626_ sky130_fd_sc_hd__and2_1
X_18375_ _08750_ _08748_ _08759_ _08769_ _08770_ VGND VGND VPWR VPWR _08771_ sky130_fd_sc_hd__a2111oi_1
X_11819_ prev_error\[18\] VGND VGND VPWR VPWR _01758_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15587_ net452 net191 net187 net457 VGND VGND VPWR VPWR _05704_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_7_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12799_ net216 _02223_ _02737_ VGND VGND VPWR VPWR _02738_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17326_ _07614_ _07615_ _07604_ VGND VGND VPWR VPWR _07617_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_141_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14538_ _04548_ _04539_ _04546_ VGND VGND VPWR VPWR _04550_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17257_ _07539_ _07540_ VGND VGND VPWR VPWR _07541_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14469_ _04472_ _04473_ VGND VGND VPWR VPWR _04474_ sky130_fd_sc_hd__and2b_1
X_16208_ net283 _06386_ VGND VGND VPWR VPWR _06387_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17188_ net311 _06468_ _07461_ _07463_ VGND VGND VPWR VPWR _07465_ sky130_fd_sc_hd__a22o_1
X_16139_ _06310_ VGND VGND VPWR VPWR _06311_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone7 _01742_ _06407_ VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__xnor2_4
XFILLER_0_149_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10150_ _08834_ _08977_ _07525_ VGND VGND VPWR VPWR _08999_ sky130_fd_sc_hd__nor3_1
X_10081_ net341 _06645_ _06557_ VGND VGND VPWR VPWR _08240_ sky130_fd_sc_hd__a21oi_1
X_13840_ _03770_ _03789_ _03802_ _03805_ VGND VGND VPWR VPWR _03806_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_69_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13771_ _03676_ _03722_ _03727_ _03736_ VGND VGND VPWR VPWR _03737_ sky130_fd_sc_hd__o31a_1
XFILLER_0_58_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10983_ _00828_ _00856_ VGND VGND VPWR VPWR _00922_ sky130_fd_sc_hd__xnor2_4
X_15510_ _05617_ net180 net463 _05618_ VGND VGND VPWR VPWR _05619_ sky130_fd_sc_hd__and4b_1
XFILLER_0_69_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12722_ _02634_ _02658_ _02660_ VGND VGND VPWR VPWR _02661_ sky130_fd_sc_hd__a21oi_1
X_16490_ _06649_ _06650_ VGND VGND VPWR VPWR _06697_ sky130_fd_sc_hd__xnor2_2
X_15441_ _05459_ _05460_ _05452_ VGND VGND VPWR VPWR _05543_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_133_Right_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12653_ _02364_ _01799_ _02585_ _02586_ VGND VGND VPWR VPWR _02592_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_0_139_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11604_ _01526_ _01527_ _01539_ VGND VGND VPWR VPWR _01543_ sky130_fd_sc_hd__a21o_1
X_18160_ i_error\[14\] _08533_ VGND VGND VPWR VPWR _08534_ sky130_fd_sc_hd__nand2_1
X_15372_ _05465_ _05466_ VGND VGND VPWR VPWR _05467_ sky130_fd_sc_hd__nand2_1
X_12584_ _02517_ _02522_ VGND VGND VPWR VPWR _02523_ sky130_fd_sc_hd__and2b_1
XFILLER_0_154_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17111_ _07366_ _07379_ VGND VGND VPWR VPWR _07380_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14323_ _04307_ _04309_ _04312_ VGND VGND VPWR VPWR _04314_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_135_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11535_ _01424_ _01470_ _01471_ _01473_ VGND VGND VPWR VPWR _01474_ sky130_fd_sc_hd__o22a_1
X_18091_ _08454_ _08457_ VGND VGND VPWR VPWR _08458_ sky130_fd_sc_hd__nand2_1
X_17042_ _07282_ _07302_ _07301_ VGND VGND VPWR VPWR _07304_ sky130_fd_sc_hd__a21o_1
X_14254_ _04234_ _04237_ VGND VGND VPWR VPWR _04238_ sky130_fd_sc_hd__and2b_1
XFILLER_0_52_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap108 _03703_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__buf_1
XFILLER_0_151_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11466_ _01402_ _01403_ _01401_ _01404_ VGND VGND VPWR VPWR _01405_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_1_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13205_ _03149_ _03154_ _03155_ VGND VGND VPWR VPWR _03158_ sky130_fd_sc_hd__or3_1
X_10417_ _00354_ _00355_ VGND VGND VPWR VPWR _00356_ sky130_fd_sc_hd__nor2_1
X_14185_ _04104_ _04120_ VGND VGND VPWR VPWR _04162_ sky130_fd_sc_hd__nand2_1
X_11397_ _01265_ _01267_ _01266_ VGND VGND VPWR VPWR _01336_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13136_ _03051_ _03082_ _03083_ VGND VGND VPWR VPWR _03084_ sky130_fd_sc_hd__a21boi_1
X_10348_ _00278_ _00284_ _00285_ VGND VGND VPWR VPWR _00287_ sky130_fd_sc_hd__or3_1
X_18993_ _09198_ _09449_ VGND VGND VPWR VPWR _09451_ sky130_fd_sc_hd__xnor2_1
X_13067_ net236 _01909_ VGND VGND VPWR VPWR _03008_ sky130_fd_sc_hd__nand2_1
X_17944_ _08286_ _08289_ VGND VGND VPWR VPWR _08297_ sky130_fd_sc_hd__nand2_1
X_10279_ _00204_ _00217_ VGND VGND VPWR VPWR _00218_ sky130_fd_sc_hd__xor2_1
X_12018_ net200 _01836_ VGND VGND VPWR VPWR _01957_ sky130_fd_sc_hd__nand2_1
X_17875_ _08129_ _08146_ VGND VGND VPWR VPWR _08221_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16826_ net294 _06437_ VGND VGND VPWR VPWR _07067_ sky130_fd_sc_hd__nand2_1
X_16757_ _02406_ _06283_ VGND VGND VPWR VPWR _06991_ sky130_fd_sc_hd__xor2_4
X_13969_ _03940_ _03923_ VGND VGND VPWR VPWR _03941_ sky130_fd_sc_hd__nor2_1
X_15708_ _05832_ _05836_ VGND VGND VPWR VPWR _05837_ sky130_fd_sc_hd__xnor2_1
X_16688_ _06850_ _06849_ VGND VGND VPWR VPWR _06915_ sky130_fd_sc_hd__xor2_1
XFILLER_0_152_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15639_ _05757_ _05759_ VGND VGND VPWR VPWR _05761_ sky130_fd_sc_hd__nor2_1
X_18427_ _08827_ _08743_ VGND VGND VPWR VPWR _08828_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Left_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18358_ i_error\[12\] _08606_ VGND VGND VPWR VPWR _08752_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17309_ _07578_ _07579_ _07596_ VGND VGND VPWR VPWR _07598_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18289_ _08674_ _08624_ _08626_ VGND VGND VPWR VPWR _08676_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09993_ _05655_ _07261_ VGND VGND VPWR VPWR _07272_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_23_Left_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_32_Left_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11320_ net396 _01178_ _01179_ net392 _08185_ VGND VGND VPWR VPWR _01259_ sky130_fd_sc_hd__a32o_1
XFILLER_0_16_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_2_0_clock clknet_0_clock VGND VGND VPWR VPWR clknet_4_2_0_clock sky130_fd_sc_hd__clkbuf_8
XFILLER_0_132_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11251_ _01187_ _01188_ _01189_ VGND VGND VPWR VPWR _01190_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10202_ net345 _08196_ VGND VGND VPWR VPWR _09540_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11182_ _01119_ _01120_ VGND VGND VPWR VPWR _01121_ sky130_fd_sc_hd__nor2_1
X_10133_ _08768_ _08790_ VGND VGND VPWR VPWR _08812_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15990_ _01676_ _01410_ VGND VGND VPWR VPWR _06147_ sky130_fd_sc_hd__or2b_2
X_10064_ _08020_ _08031_ _08042_ VGND VGND VPWR VPWR _08053_ sky130_fd_sc_hd__nor3_1
X_14941_ _04987_ _04990_ _04992_ VGND VGND VPWR VPWR _04993_ sky130_fd_sc_hd__a21oi_1
X_17660_ _07889_ _07982_ _07983_ VGND VGND VPWR VPWR _07984_ sky130_fd_sc_hd__nand3_1
X_14872_ net439 net163 _04829_ _04831_ VGND VGND VPWR VPWR _04917_ sky130_fd_sc_hd__o2bb2a_1
X_16611_ _06822_ _06795_ VGND VGND VPWR VPWR _06830_ sky130_fd_sc_hd__or2b_1
X_13823_ _03768_ _03769_ VGND VGND VPWR VPWR _03789_ sky130_fd_sc_hd__and2_1
X_17591_ _07808_ _07907_ VGND VGND VPWR VPWR _07908_ sky130_fd_sc_hd__nor2_1
X_19330_ clknet_4_3_0_clock _00031_ VGND VGND VPWR VPWR kd_2\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16542_ net303 _06311_ VGND VGND VPWR VPWR _06754_ sky130_fd_sc_hd__nand2_1
X_13754_ _03684_ _03686_ VGND VGND VPWR VPWR _03720_ sky130_fd_sc_hd__nor2_1
X_10966_ _00902_ _00904_ VGND VGND VPWR VPWR _00905_ sky130_fd_sc_hd__and2b_1
XFILLER_0_85_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12705_ kd_1\[17\] _02641_ _02643_ VGND VGND VPWR VPWR _02644_ sky130_fd_sc_hd__and3_1
X_19261_ clknet_4_10_0_clock _00143_ VGND VGND VPWR VPWR prev_d_error\[10\] sky130_fd_sc_hd__dfxtp_1
X_16473_ _06365_ _06674_ VGND VGND VPWR VPWR _06679_ sky130_fd_sc_hd__xor2_1
X_13685_ _03633_ _03649_ VGND VGND VPWR VPWR _03650_ sky130_fd_sc_hd__and2_1
XFILLER_0_155_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10897_ net393 _05292_ _05303_ VGND VGND VPWR VPWR _00836_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18212_ _07460_ _08501_ VGND VGND VPWR VPWR _08591_ sky130_fd_sc_hd__xor2_1
X_15424_ _05505_ _05524_ VGND VGND VPWR VPWR _05525_ sky130_fd_sc_hd__nand2_1
X_12636_ _02527_ _02574_ VGND VGND VPWR VPWR _02575_ sky130_fd_sc_hd__nand2_2
X_19192_ prev_d_error\[18\] net501 VGND VGND VPWR VPWR _09594_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18143_ _08507_ _08514_ VGND VGND VPWR VPWR _08516_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15355_ _05387_ _05448_ VGND VGND VPWR VPWR _05449_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12567_ _02384_ _02505_ VGND VGND VPWR VPWR _02506_ sky130_fd_sc_hd__or2_1
X_14306_ _04099_ _04100_ _04098_ _04041_ VGND VGND VPWR VPWR _04295_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_81_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11518_ _01455_ _01448_ _01453_ VGND VGND VPWR VPWR _01457_ sky130_fd_sc_hd__or3_1
X_18074_ _07972_ _07975_ _08437_ _08439_ VGND VGND VPWR VPWR _08440_ sky130_fd_sc_hd__nand4bb_4
X_15286_ _05362_ _05370_ _05372_ VGND VGND VPWR VPWR _05373_ sky130_fd_sc_hd__a21o_1
X_12498_ _02426_ _02436_ VGND VGND VPWR VPWR _02437_ sky130_fd_sc_hd__and2_1
XFILLER_0_151_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17025_ net320 _06335_ VGND VGND VPWR VPWR _07286_ sky130_fd_sc_hd__nand2_1
X_14237_ net451 net120 net116 net456 VGND VGND VPWR VPWR _04219_ sky130_fd_sc_hd__a22oi_1
X_11449_ net366 net362 _00811_ _00818_ VGND VGND VPWR VPWR _01388_ sky130_fd_sc_hd__and4_1
X_14168_ _04141_ _04142_ VGND VGND VPWR VPWR _04143_ sky130_fd_sc_hd__or2_1
X_13119_ _02931_ VGND VGND VPWR VPWR _03065_ sky130_fd_sc_hd__clkinv_4
X_14099_ net422 net130 VGND VGND VPWR VPWR _04071_ sky130_fd_sc_hd__nand2_1
X_18976_ _09427_ _09431_ VGND VGND VPWR VPWR _09432_ sky130_fd_sc_hd__xnor2_1
X_17927_ net313 _07568_ VGND VGND VPWR VPWR _08278_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17858_ _08187_ _08201_ VGND VGND VPWR VPWR _08202_ sky130_fd_sc_hd__and2b_1
XFILLER_0_89_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16809_ _07039_ _07037_ VGND VGND VPWR VPWR _07048_ sky130_fd_sc_hd__xor2_1
X_17789_ _08124_ _08125_ VGND VGND VPWR VPWR _08126_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09976_ _07030_ _07074_ VGND VGND VPWR VPWR _07085_ sky130_fd_sc_hd__xor2_1
X_10820_ _00757_ _00758_ VGND VGND VPWR VPWR _00759_ sky130_fd_sc_hd__and2_2
XFILLER_0_67_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10751_ net347 _00325_ _00606_ VGND VGND VPWR VPWR _00690_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13470_ _03371_ _03279_ _03370_ VGND VGND VPWR VPWR _03429_ sky130_fd_sc_hd__o21ai_1
X_10682_ _00611_ _00620_ VGND VGND VPWR VPWR _00621_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12421_ _02345_ _02359_ VGND VGND VPWR VPWR _02360_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15140_ _05108_ _05211_ VGND VGND VPWR VPWR _05212_ sky130_fd_sc_hd__nor2_1
X_12352_ _02289_ _02290_ VGND VGND VPWR VPWR _02291_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11303_ _01220_ _01227_ _01228_ VGND VGND VPWR VPWR _01242_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_132_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15071_ _05034_ _05018_ _05033_ VGND VGND VPWR VPWR _05136_ sky130_fd_sc_hd__and3_1
X_12283_ _02221_ VGND VGND VPWR VPWR _02222_ sky130_fd_sc_hd__buf_2
XFILLER_0_133_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14022_ _03992_ _03993_ net407 net156 VGND VGND VPWR VPWR _03994_ sky130_fd_sc_hd__and4bb_1
X_11234_ net383 _08196_ VGND VGND VPWR VPWR _01173_ sky130_fd_sc_hd__nand2_1
X_18830_ _04209_ _09226_ _09269_ VGND VGND VPWR VPWR _09271_ sky130_fd_sc_hd__or3_2
X_11165_ _01081_ _01102_ _01013_ _01103_ VGND VGND VPWR VPWR _01104_ sky130_fd_sc_hd__a211oi_2
X_10116_ _07437_ _07459_ _07448_ _05677_ VGND VGND VPWR VPWR _08625_ sky130_fd_sc_hd__a2bb2o_1
X_15973_ _06008_ _06126_ VGND VGND VPWR VPWR _06129_ sky130_fd_sc_hd__nor2_2
X_18761_ _09067_ _09069_ _09060_ VGND VGND VPWR VPWR _09195_ sky130_fd_sc_hd__o21a_1
X_11096_ _01023_ _01034_ VGND VGND VPWR VPWR _01035_ sky130_fd_sc_hd__xnor2_2
X_14924_ _04810_ _04974_ VGND VGND VPWR VPWR _04975_ sky130_fd_sc_hd__nand2_1
X_17712_ _08034_ _08035_ VGND VGND VPWR VPWR _08041_ sky130_fd_sc_hd__nand2_1
X_10047_ net364 _04874_ _07855_ VGND VGND VPWR VPWR _07866_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18692_ _09104_ _09107_ _09118_ VGND VGND VPWR VPWR _09119_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14855_ _04820_ _04897_ _04898_ VGND VGND VPWR VPWR _04899_ sky130_fd_sc_hd__o21ba_1
X_17643_ _07963_ _07961_ _07964_ VGND VGND VPWR VPWR _07966_ sky130_fd_sc_hd__or3_4
X_13806_ _03766_ _03770_ _03771_ VGND VGND VPWR VPWR _03772_ sky130_fd_sc_hd__o21a_1
X_17574_ _07886_ _07889_ VGND VGND VPWR VPWR _07890_ sky130_fd_sc_hd__nand2_1
X_14786_ _04495_ _04820_ _04821_ _04822_ VGND VGND VPWR VPWR _04823_ sky130_fd_sc_hd__o22a_1
X_11998_ _01933_ _01934_ _01935_ VGND VGND VPWR VPWR _01937_ sky130_fd_sc_hd__o21a_1
XFILLER_0_147_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16525_ _06709_ _06735_ VGND VGND VPWR VPWR _06736_ sky130_fd_sc_hd__xor2_1
X_19313_ clknet_4_1_0_clock _00014_ VGND VGND VPWR VPWR kd_1\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13737_ _03690_ _03701_ _03702_ VGND VGND VPWR VPWR _03703_ sky130_fd_sc_hd__nor3_1
XFILLER_0_86_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10949_ _00887_ _00781_ VGND VGND VPWR VPWR _00888_ sky130_fd_sc_hd__xor2_1
X_19244_ clknet_4_12_0_clock _00126_ VGND VGND VPWR VPWR i_error\[12\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_85_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16456_ _06653_ _06658_ _06659_ VGND VGND VPWR VPWR _06660_ sky130_fd_sc_hd__o21a_1
XFILLER_0_156_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13668_ _03628_ _03630_ VGND VGND VPWR VPWR _03631_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15407_ net441 net446 net193 net189 VGND VGND VPWR VPWR _05506_ sky130_fd_sc_hd__and4_1
X_12619_ _02416_ _02533_ _02554_ _02555_ _02557_ VGND VGND VPWR VPWR _02558_ sky130_fd_sc_hd__a32oi_2
X_19175_ net502 net445 net490 _09584_ VGND VGND VPWR VPWR _00142_ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16387_ _06549_ _06582_ _06583_ VGND VGND VPWR VPWR _06584_ sky130_fd_sc_hd__a21oi_1
X_13599_ net252 _02409_ _01908_ net269 VGND VGND VPWR VPWR _03558_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_42_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18126_ _08484_ _08490_ _08492_ VGND VGND VPWR VPWR _08497_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15338_ net428 net197 net194 net432 VGND VGND VPWR VPWR _05430_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_130_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18057_ _08410_ _08413_ _08406_ VGND VGND VPWR VPWR _08421_ sky130_fd_sc_hd__a21o_1
X_15269_ _05252_ _05353_ VGND VGND VPWR VPWR _05354_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17008_ _07158_ _07262_ _07266_ VGND VGND VPWR VPWR _07267_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09830_ _05248_ _05468_ VGND VGND VPWR VPWR _05479_ sky130_fd_sc_hd__nand2_1
Xfanout507 net1 VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09761_ net6 net64 VGND VGND VPWR VPWR _04720_ sky130_fd_sc_hd__or2b_2
X_18959_ _09411_ _09412_ VGND VGND VPWR VPWR _09413_ sky130_fd_sc_hd__xor2_1
X_09692_ net54 _03881_ _03914_ net382 VGND VGND VPWR VPWR _00071_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer12 _08753_ VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__buf_1
Xrebuffer23 _08686_ VGND VGND VPWR VPWR net530 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09959_ net361 _05699_ VGND VGND VPWR VPWR _06898_ sky130_fd_sc_hd__or2_1
X_12970_ _02841_ _02861_ VGND VGND VPWR VPWR _02909_ sky130_fd_sc_hd__xor2_1
X_11921_ _01859_ VGND VGND VPWR VPWR _01860_ sky130_fd_sc_hd__clkbuf_4
X_14640_ _04646_ _04648_ VGND VGND VPWR VPWR _04662_ sky130_fd_sc_hd__or2_1
X_11852_ _01789_ _01779_ _01790_ VGND VGND VPWR VPWR _01791_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_157_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10803_ _00726_ _00727_ _00740_ VGND VGND VPWR VPWR _00742_ sky130_fd_sc_hd__or3_2
X_14571_ _04584_ _04585_ VGND VGND VPWR VPWR _04586_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11783_ _01711_ _00406_ _00407_ VGND VGND VPWR VPWR _01722_ sky130_fd_sc_hd__and3_1
XFILLER_0_83_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16310_ _06495_ _06498_ VGND VGND VPWR VPWR _06499_ sky130_fd_sc_hd__xnor2_1
X_13522_ _03436_ _03440_ VGND VGND VPWR VPWR _03481_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17290_ _07555_ _07562_ _07576_ VGND VGND VPWR VPWR _07577_ sky130_fd_sc_hd__o21bai_1
X_10734_ net375 _05996_ VGND VGND VPWR VPWR _00673_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16241_ _06418_ _06422_ VGND VGND VPWR VPWR _06423_ sky130_fd_sc_hd__xnor2_1
X_13453_ net207 _03220_ _03224_ VGND VGND VPWR VPWR _03412_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10665_ net352 _00245_ _00503_ VGND VGND VPWR VPWR _00604_ sky130_fd_sc_hd__and3_1
XFILLER_0_137_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12404_ _02341_ _02342_ VGND VGND VPWR VPWR _02343_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16172_ net289 _06335_ VGND VGND VPWR VPWR _06347_ sky130_fd_sc_hd__nand2_1
X_13384_ _03271_ _03334_ _03337_ VGND VGND VPWR VPWR _03338_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_88_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10596_ _00469_ _00534_ VGND VGND VPWR VPWR _00535_ sky130_fd_sc_hd__xnor2_4
X_15123_ _05181_ _05186_ _05192_ VGND VGND VPWR VPWR _05194_ sky130_fd_sc_hd__o21ba_1
X_12335_ _01977_ _02271_ VGND VGND VPWR VPWR _02274_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15054_ net463 net153 VGND VGND VPWR VPWR _05118_ sky130_fd_sc_hd__nand2_1
X_12266_ _02186_ _02204_ VGND VGND VPWR VPWR _02205_ sky130_fd_sc_hd__nand2_1
X_14005_ _03971_ _03976_ VGND VGND VPWR VPWR _03977_ sky130_fd_sc_hd__and2_1
X_11217_ net358 _00614_ _01155_ VGND VGND VPWR VPWR _01156_ sky130_fd_sc_hd__and3_1
X_12197_ _02134_ _02135_ VGND VGND VPWR VPWR _02136_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput81 net81 VGND VGND VPWR VPWR out_clocked[10] sky130_fd_sc_hd__buf_2
X_18813_ _04190_ _09251_ VGND VGND VPWR VPWR _09253_ sky130_fd_sc_hd__xor2_1
Xoutput92 net92 VGND VGND VPWR VPWR out_clocked[3] sky130_fd_sc_hd__buf_2
X_11148_ _01028_ _01086_ VGND VGND VPWR VPWR _01087_ sky130_fd_sc_hd__nand2_1
X_18744_ _09166_ _09176_ VGND VGND VPWR VPWR _09177_ sky130_fd_sc_hd__xnor2_2
X_15956_ _06056_ _06108_ _06109_ VGND VGND VPWR VPWR _06110_ sky130_fd_sc_hd__a21o_1
X_11079_ _01010_ _00998_ VGND VGND VPWR VPWR _01018_ sky130_fd_sc_hd__and2b_1
X_14907_ _04847_ _04848_ _04850_ VGND VGND VPWR VPWR _04956_ sky130_fd_sc_hd__a21oi_1
X_15887_ _06031_ _06033_ VGND VGND VPWR VPWR _06034_ sky130_fd_sc_hd__nand2_1
X_18675_ _09095_ _09099_ _09100_ VGND VGND VPWR VPWR _09101_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17626_ _07945_ _07946_ VGND VGND VPWR VPWR _07947_ sky130_fd_sc_hd__nor2_1
X_14838_ _04859_ _04879_ _04877_ VGND VGND VPWR VPWR _04880_ sky130_fd_sc_hd__a21oi_1
X_14769_ _04802_ _04803_ VGND VGND VPWR VPWR _04804_ sky130_fd_sc_hd__or2_1
X_17557_ _07839_ _07870_ VGND VGND VPWR VPWR _07871_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16508_ _06625_ _06716_ VGND VGND VPWR VPWR _06717_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17488_ _07781_ _07794_ VGND VGND VPWR VPWR _07795_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19227_ clknet_4_5_0_clock _00109_ VGND VGND VPWR VPWR prev_error\[14\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_144_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16439_ _06617_ _06639_ VGND VGND VPWR VPWR _06641_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19158_ net502 _09111_ VGND VGND VPWR VPWR _09574_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18109_ _08465_ _08477_ VGND VGND VPWR VPWR _08478_ sky130_fd_sc_hd__xor2_2
XFILLER_0_124_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19089_ net499 prev_error\[6\] VGND VGND VPWR VPWR _09531_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout304 ki\[8\] VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__buf_2
Xfanout315 net317 VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__clkbuf_4
Xfanout326 net327 VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__buf_2
Xfanout337 kp\[17\] VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__clkbuf_4
X_09813_ _04181_ _04709_ _05281_ _04731_ VGND VGND VPWR VPWR _05292_ sky130_fd_sc_hd__a211o_2
Xfanout348 net350 VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__clkbuf_4
Xfanout359 kp\[11\] VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__dlymetal6s2s_1
X_09744_ _04511_ _04522_ VGND VGND VPWR VPWR _04533_ sky130_fd_sc_hd__or2b_2
XFILLER_0_69_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09675_ net44 _03614_ _03647_ net287 VGND VGND VPWR VPWR _00042_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_6_Left_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10450_ _00387_ _00388_ VGND VGND VPWR VPWR _00389_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10381_ net340 _00243_ VGND VGND VPWR VPWR _00320_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12120_ _02058_ _01830_ VGND VGND VPWR VPWR _02059_ sky130_fd_sc_hd__xor2_1
XFILLER_0_130_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12051_ _01772_ _01988_ _01989_ VGND VGND VPWR VPWR _01990_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11002_ _00939_ _00940_ VGND VGND VPWR VPWR _00941_ sky130_fd_sc_hd__or2b_1
X_15810_ _05546_ _05947_ _05948_ VGND VGND VPWR VPWR _05949_ sky130_fd_sc_hd__o21ba_1
X_16790_ _07025_ _07026_ VGND VGND VPWR VPWR _07027_ sky130_fd_sc_hd__nand2_1
X_15741_ net480 net187 _05871_ _05872_ VGND VGND VPWR VPWR _05873_ sky130_fd_sc_hd__a31o_1
X_12953_ _02827_ _02829_ VGND VGND VPWR VPWR _02892_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11904_ _01833_ _01842_ VGND VGND VPWR VPWR _01843_ sky130_fd_sc_hd__and2_1
X_15672_ _05756_ _05768_ _05767_ VGND VGND VPWR VPWR _05797_ sky130_fd_sc_hd__a21o_1
X_18460_ _08858_ _08862_ _08853_ _08851_ VGND VGND VPWR VPWR _08864_ sky130_fd_sc_hd__o2bb2a_1
X_12884_ _02722_ _02721_ VGND VGND VPWR VPWR _02823_ sky130_fd_sc_hd__and2b_1
XFILLER_0_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14623_ _04590_ _04640_ _04642_ VGND VGND VPWR VPWR _04644_ sky130_fd_sc_hd__a21o_1
X_17411_ _07697_ _07698_ _07708_ VGND VGND VPWR VPWR _07710_ sky130_fd_sc_hd__o21ba_1
X_11835_ _01771_ _01773_ VGND VGND VPWR VPWR _01774_ sky130_fd_sc_hd__or2_1
X_18391_ _08787_ _08743_ VGND VGND VPWR VPWR _08788_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17342_ _07587_ _07586_ VGND VGND VPWR VPWR _07634_ sky130_fd_sc_hd__and2b_1
X_14554_ net413 net182 net175 net417 VGND VGND VPWR VPWR _04568_ sky130_fd_sc_hd__a22oi_1
X_11766_ _05908_ _05919_ _01704_ VGND VGND VPWR VPWR _01705_ sky130_fd_sc_hd__a21o_2
XFILLER_0_138_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13505_ _03409_ _03463_ VGND VGND VPWR VPWR _03464_ sky130_fd_sc_hd__nand2_2
XFILLER_0_82_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17273_ net298 _06992_ _07093_ net295 VGND VGND VPWR VPWR _07559_ sky130_fd_sc_hd__a22o_1
X_10717_ _00597_ _00655_ VGND VGND VPWR VPWR _00656_ sky130_fd_sc_hd__nand2_2
XFILLER_0_153_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14485_ _04488_ _04491_ VGND VGND VPWR VPWR _04492_ sky130_fd_sc_hd__nor2_1
X_11697_ _01635_ _01620_ VGND VGND VPWR VPWR _01636_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19012_ _09133_ _09119_ VGND VGND VPWR VPWR _09471_ sky130_fd_sc_hd__and2b_1
X_16224_ _06399_ _06404_ VGND VGND VPWR VPWR _06405_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13436_ _03392_ _03393_ VGND VGND VPWR VPWR _03395_ sky130_fd_sc_hd__and2_1
X_10648_ _00583_ _00586_ _00584_ VGND VGND VPWR VPWR _00587_ sky130_fd_sc_hd__o21ba_1
Xrebuffer3 _08432_ VGND VGND VPWR VPWR net570 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16155_ net299 _06328_ _06320_ net296 VGND VGND VPWR VPWR _06329_ sky130_fd_sc_hd__a22o_1
X_13367_ _03313_ _03318_ _03319_ VGND VGND VPWR VPWR _03320_ sky130_fd_sc_hd__o21ai_4
X_10579_ net340 _00410_ _00325_ net343 VGND VGND VPWR VPWR _00518_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15106_ net423 net193 _05174_ _05172_ VGND VGND VPWR VPWR _05175_ sky130_fd_sc_hd__a31o_1
X_12318_ _02011_ _02184_ VGND VGND VPWR VPWR _02257_ sky130_fd_sc_hd__xnor2_1
X_16086_ net345 _05600_ _06252_ VGND VGND VPWR VPWR _06253_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13298_ _03246_ _03249_ _03159_ _03250_ VGND VGND VPWR VPWR _03251_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_48_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15037_ _05092_ _05097_ _05098_ VGND VGND VPWR VPWR _05099_ sky130_fd_sc_hd__a21oi_2
X_12249_ _02062_ _02064_ VGND VGND VPWR VPWR _02188_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16988_ _07224_ _07231_ _07243_ VGND VGND VPWR VPWR _07245_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_147_Right_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18727_ _06103_ _09157_ VGND VGND VPWR VPWR _09158_ sky130_fd_sc_hd__and2_1
X_15939_ _06083_ _06090_ VGND VGND VPWR VPWR _06091_ sky130_fd_sc_hd__and2_1
XFILLER_0_155_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18658_ _09074_ _09080_ _09081_ VGND VGND VPWR VPWR _09082_ sky130_fd_sc_hd__nand3_1
XFILLER_0_94_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17609_ _07925_ _07926_ VGND VGND VPWR VPWR _07928_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18589_ _06170_ _09005_ VGND VGND VPWR VPWR _09006_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout123 net126 VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__buf_2
Xfanout134 net135 VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__buf_2
Xfanout145 kd_2\[12\] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__buf_2
Xfanout156 net159 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_4
Xfanout167 net168 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_2
Xfanout178 kd_2\[5\] VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_4
Xfanout189 net190 VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_114_Right_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09727_ _04324_ _04335_ VGND VGND VPWR VPWR _04346_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09658_ _03614_ VGND VGND VPWR VPWR _03625_ sky130_fd_sc_hd__buf_2
XFILLER_0_97_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11620_ _01556_ _01558_ VGND VGND VPWR VPWR _01559_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11551_ net400 _00244_ _01487_ _01489_ VGND VGND VPWR VPWR _01490_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10502_ _00439_ _00440_ _05039_ _05050_ _07327_ VGND VGND VPWR VPWR _00441_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14270_ _03983_ _03984_ _03985_ VGND VGND VPWR VPWR _04255_ sky130_fd_sc_hd__o21a_1
X_11482_ _01416_ _01419_ VGND VGND VPWR VPWR _01421_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13221_ _03141_ _03172_ VGND VGND VPWR VPWR _03174_ sky130_fd_sc_hd__and2_1
X_10433_ net372 _05336_ _00370_ _00371_ VGND VGND VPWR VPWR _00372_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_116_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13152_ net244 net239 _02089_ _01907_ VGND VGND VPWR VPWR _03101_ sky130_fd_sc_hd__and4_1
X_10364_ _07294_ _00302_ VGND VGND VPWR VPWR _00303_ sky130_fd_sc_hd__xnor2_1
X_12103_ _01768_ _02041_ VGND VGND VPWR VPWR _02042_ sky130_fd_sc_hd__xnor2_1
X_13083_ _02899_ _03024_ VGND VGND VPWR VPWR _03026_ sky130_fd_sc_hd__nor2_1
X_17960_ _08311_ _08313_ VGND VGND VPWR VPWR _08314_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10295_ _00232_ _00233_ VGND VGND VPWR VPWR _00234_ sky130_fd_sc_hd__nor2_1
X_16911_ net278 _06993_ _07095_ net274 VGND VGND VPWR VPWR _07160_ sky130_fd_sc_hd__a22o_1
X_12034_ net264 VGND VGND VPWR VPWR _01973_ sky130_fd_sc_hd__inv_2
X_17891_ net313 _07182_ VGND VGND VPWR VPWR _08238_ sky130_fd_sc_hd__nand2_1
X_16842_ _07066_ _07081_ _07083_ VGND VGND VPWR VPWR _07084_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_69_Left_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16773_ _06907_ _07007_ VGND VGND VPWR VPWR _07009_ sky130_fd_sc_hd__xnor2_1
X_13985_ _03898_ _03956_ _03897_ VGND VGND VPWR VPWR _03957_ sky130_fd_sc_hd__o21ba_1
X_18512_ _08919_ _08826_ VGND VGND VPWR VPWR _08921_ sky130_fd_sc_hd__nor2_1
X_12936_ _02872_ _02874_ VGND VGND VPWR VPWR _02875_ sky130_fd_sc_hd__nor2_1
X_15724_ _05846_ _05851_ _05854_ VGND VGND VPWR VPWR _05855_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18443_ _08843_ _08841_ _08828_ _08826_ VGND VGND VPWR VPWR _08846_ sky130_fd_sc_hd__o2bb2a_1
X_15655_ _05772_ _05777_ _05778_ VGND VGND VPWR VPWR _05779_ sky130_fd_sc_hd__or3_1
X_12867_ _02804_ _02805_ VGND VGND VPWR VPWR _02806_ sky130_fd_sc_hd__or2_1
X_14606_ _04620_ _04624_ VGND VGND VPWR VPWR _04625_ sky130_fd_sc_hd__nor2_1
X_11818_ _01755_ _01756_ VGND VGND VPWR VPWR _01757_ sky130_fd_sc_hd__nand2_4
X_15586_ net450 net195 VGND VGND VPWR VPWR _05703_ sky130_fd_sc_hd__nand2_1
X_18374_ _08764_ _08762_ VGND VGND VPWR VPWR _08770_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12798_ net220 _02331_ VGND VGND VPWR VPWR _02737_ sky130_fd_sc_hd__and2_1
XFILLER_0_141_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14537_ _04539_ _04546_ _04548_ VGND VGND VPWR VPWR _04549_ sky130_fd_sc_hd__a21oi_1
X_17325_ _07604_ _07614_ _07615_ VGND VGND VPWR VPWR _07616_ sky130_fd_sc_hd__and3_1
X_11749_ _01134_ _01209_ _01681_ _01685_ _01687_ VGND VGND VPWR VPWR _01688_ sky130_fd_sc_hd__o41ai_4
XFILLER_0_44_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_78_Left_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14468_ _04441_ _04462_ _04439_ VGND VGND VPWR VPWR _04473_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17256_ net308 _06467_ _06619_ net305 VGND VGND VPWR VPWR _07540_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_154_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13419_ _03356_ _03360_ _03375_ VGND VGND VPWR VPWR _03376_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16207_ _06353_ VGND VGND VPWR VPWR _06386_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17187_ net311 _06468_ _07461_ _07463_ VGND VGND VPWR VPWR _07464_ sky130_fd_sc_hd__nand4_2
X_14399_ _04395_ _04386_ _04388_ VGND VGND VPWR VPWR _04397_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16138_ _06309_ VGND VGND VPWR VPWR _06310_ sky130_fd_sc_hd__buf_2
XFILLER_0_12_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16069_ _06232_ _06233_ VGND VGND VPWR VPWR _06234_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_87_Left_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_96_Left_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10080_ net341 _06645_ _06557_ VGND VGND VPWR VPWR _08229_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13770_ _03733_ _03735_ VGND VGND VPWR VPWR _03736_ sky130_fd_sc_hd__nand2_1
X_10982_ _00826_ _00897_ _00898_ _00920_ VGND VGND VPWR VPWR _00921_ sky130_fd_sc_hd__o31ai_4
X_12721_ _02546_ _02659_ kd_1\[18\] VGND VGND VPWR VPWR _02660_ sky130_fd_sc_hd__and3b_1
X_15440_ _05530_ _05541_ VGND VGND VPWR VPWR _05542_ sky130_fd_sc_hd__or2_1
X_12652_ _02583_ _02589_ _02590_ VGND VGND VPWR VPWR _02591_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11603_ _01517_ _01541_ VGND VGND VPWR VPWR _01542_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15371_ _05383_ _05464_ VGND VGND VPWR VPWR _05466_ sky130_fd_sc_hd__nand2_1
X_12583_ _02520_ _02521_ VGND VGND VPWR VPWR _02522_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17110_ _07368_ _07378_ VGND VGND VPWR VPWR _07379_ sky130_fd_sc_hd__xnor2_2
X_14322_ _03896_ _04311_ VGND VGND VPWR VPWR _04312_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11534_ _01422_ _01472_ VGND VGND VPWR VPWR _01473_ sky130_fd_sc_hd__and2_1
X_18090_ _08454_ _08455_ _08456_ VGND VGND VPWR VPWR _08457_ sky130_fd_sc_hd__nand3_1
XFILLER_0_136_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17041_ _07282_ _07301_ _07302_ VGND VGND VPWR VPWR _07303_ sky130_fd_sc_hd__nand3_1
XFILLER_0_123_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14253_ _03965_ _04235_ VGND VGND VPWR VPWR _04237_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11465_ _01341_ _01400_ _01387_ _01399_ VGND VGND VPWR VPWR _01404_ sky130_fd_sc_hd__a211oi_1
Xmax_cap109 _01122_ VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__buf_1
XFILLER_0_33_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13204_ _03104_ _03103_ VGND VGND VPWR VPWR _03157_ sky130_fd_sc_hd__xnor2_1
X_10416_ _00264_ _00263_ VGND VGND VPWR VPWR _00355_ sky130_fd_sc_hd__xor2_1
X_14184_ _04122_ _04160_ VGND VGND VPWR VPWR _04161_ sky130_fd_sc_hd__nand2_1
X_11396_ _01333_ _01334_ VGND VGND VPWR VPWR _01335_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13135_ _03079_ _03076_ VGND VGND VPWR VPWR _03083_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10347_ _00278_ _00284_ _00285_ VGND VGND VPWR VPWR _00286_ sky130_fd_sc_hd__o21ai_1
X_18992_ _09199_ _09044_ VGND VGND VPWR VPWR _09449_ sky130_fd_sc_hd__and2b_1
XFILLER_0_29_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13066_ net247 _01852_ _02990_ _03006_ VGND VGND VPWR VPWR _03007_ sky130_fd_sc_hd__a31o_1
X_17943_ _08283_ _08292_ _08293_ _08294_ VGND VGND VPWR VPWR _08296_ sky130_fd_sc_hd__o211a_1
X_10278_ _00214_ _00216_ _00212_ VGND VGND VPWR VPWR _00217_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12017_ net210 _01817_ _01943_ _01942_ VGND VGND VPWR VPWR _01956_ sky130_fd_sc_hd__a31o_1
X_17874_ _08216_ _08219_ VGND VGND VPWR VPWR _08220_ sky130_fd_sc_hd__and2b_1
X_16825_ _07055_ _07064_ _07065_ VGND VGND VPWR VPWR _07066_ sky130_fd_sc_hd__a21oi_1
Xmax_cap1 net536 VGND VGND VPWR VPWR net535 sky130_fd_sc_hd__clkbuf_1
X_16756_ _06900_ _06989_ net274 VGND VGND VPWR VPWR _06990_ sky130_fd_sc_hd__or3b_1
XFILLER_0_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13968_ net440 net444 net117 VGND VGND VPWR VPWR _03940_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_45_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15707_ _05833_ _05834_ _05835_ VGND VGND VPWR VPWR _05836_ sky130_fd_sc_hd__o21ba_1
X_12919_ _02754_ _02857_ VGND VGND VPWR VPWR _02858_ sky130_fd_sc_hd__nand2_1
X_13899_ _03178_ _03863_ _03865_ VGND VGND VPWR VPWR _03866_ sky130_fd_sc_hd__a21o_1
X_16687_ _06910_ _06913_ VGND VGND VPWR VPWR _06914_ sky130_fd_sc_hd__or2b_1
XFILLER_0_119_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18426_ _06136_ _08777_ VGND VGND VPWR VPWR _08827_ sky130_fd_sc_hd__xor2_1
X_15638_ _05757_ _05759_ VGND VGND VPWR VPWR _05760_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18357_ _08737_ _08738_ _08745_ _08748_ _08750_ VGND VGND VPWR VPWR _08751_ sky130_fd_sc_hd__o32a_1
X_15569_ _05638_ _05683_ VGND VGND VPWR VPWR _05684_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17308_ _07578_ _07579_ _07596_ VGND VGND VPWR VPWR _07597_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18288_ _08624_ _08626_ _08674_ VGND VGND VPWR VPWR _08675_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17239_ net330 _06352_ _07519_ _07520_ VGND VGND VPWR VPWR _07521_ sky130_fd_sc_hd__nand4_2
XFILLER_0_31_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09992_ _05556_ _05589_ _05644_ VGND VGND VPWR VPWR _07261_ sky130_fd_sc_hd__nor3_1
XFILLER_0_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11250_ _01059_ _01172_ _01186_ VGND VGND VPWR VPWR _01189_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10201_ _09491_ _09527_ VGND VGND VPWR VPWR _09533_ sky130_fd_sc_hd__and2b_1
X_11181_ _01114_ _01118_ VGND VGND VPWR VPWR _01120_ sky130_fd_sc_hd__and2_1
X_10132_ _08768_ _08790_ VGND VGND VPWR VPWR _08801_ sky130_fd_sc_hd__or2_1
X_10063_ _07811_ _07822_ VGND VGND VPWR VPWR _08042_ sky130_fd_sc_hd__xnor2_1
X_14940_ _04883_ _04991_ VGND VGND VPWR VPWR _04992_ sky130_fd_sc_hd__or2_1
X_14871_ _04913_ _04915_ VGND VGND VPWR VPWR _04916_ sky130_fd_sc_hd__nor2_1
X_16610_ _06827_ _06826_ VGND VGND VPWR VPWR _06829_ sky130_fd_sc_hd__xor2_1
X_13822_ _03776_ _03787_ VGND VGND VPWR VPWR _03788_ sky130_fd_sc_hd__nand2_1
X_17590_ net307 _06992_ VGND VGND VPWR VPWR _07907_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16541_ _06696_ _06701_ VGND VGND VPWR VPWR _06753_ sky130_fd_sc_hd__xnor2_2
X_13753_ _03711_ _03718_ VGND VGND VPWR VPWR _03719_ sky130_fd_sc_hd__nand2_1
X_10965_ net565 _00409_ _00903_ VGND VGND VPWR VPWR _00904_ sky130_fd_sc_hd__a21bo_1
X_12704_ _02547_ _02635_ _02642_ VGND VGND VPWR VPWR _02643_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19260_ clknet_4_3_0_clock _00142_ VGND VGND VPWR VPWR prev_d_error\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13684_ _03635_ _03642_ _03648_ VGND VGND VPWR VPWR _03649_ sky130_fd_sc_hd__o21ai_1
X_16472_ net303 _06311_ _06676_ _06379_ _06366_ VGND VGND VPWR VPWR _06677_ sky130_fd_sc_hd__a32o_1
X_10896_ net401 _05138_ _05149_ VGND VGND VPWR VPWR _00835_ sky130_fd_sc_hd__and3_1
X_18211_ i_error\[10\] _08589_ VGND VGND VPWR VPWR _08590_ sky130_fd_sc_hd__xnor2_4
X_12635_ _02525_ _02526_ VGND VGND VPWR VPWR _02574_ sky130_fd_sc_hd__or2_1
X_15423_ _05503_ _05504_ _05488_ _05502_ VGND VGND VPWR VPWR _05524_ sky130_fd_sc_hd__o211ai_1
X_19191_ net1 net409 net497 _09593_ VGND VGND VPWR VPWR _00150_ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18142_ _07048_ _07152_ VGND VGND VPWR VPWR _08514_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15354_ _05333_ _05388_ _05419_ _05447_ VGND VGND VPWR VPWR _05448_ sky130_fd_sc_hd__a31oi_2
X_12566_ net221 _01854_ _02383_ VGND VGND VPWR VPWR _02505_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14305_ _04292_ _04293_ VGND VGND VPWR VPWR _04294_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11517_ _01448_ _01453_ _01455_ VGND VGND VPWR VPWR _01456_ sky130_fd_sc_hd__o21ai_1
X_15285_ _05284_ _05371_ VGND VGND VPWR VPWR _05372_ sky130_fd_sc_hd__nand2_1
X_18073_ _07798_ _07883_ VGND VGND VPWR VPWR _08439_ sky130_fd_sc_hd__xor2_4
X_12497_ _02428_ _02433_ _02435_ _01975_ VGND VGND VPWR VPWR _02436_ sky130_fd_sc_hd__o31a_1
XFILLER_0_124_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14236_ net451 net456 net120 net116 VGND VGND VPWR VPWR _04218_ sky130_fd_sc_hd__and4_1
XFILLER_0_1_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17024_ net329 _06314_ _06317_ VGND VGND VPWR VPWR _07285_ sky130_fd_sc_hd__and3_1
X_11448_ _01355_ _01386_ VGND VGND VPWR VPWR _01387_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14167_ _04081_ _04128_ _04140_ VGND VGND VPWR VPWR _04142_ sky130_fd_sc_hd__nor3_1
X_11379_ net402 _06172_ _01258_ _01259_ VGND VGND VPWR VPWR _01318_ sky130_fd_sc_hd__a22o_1
X_13118_ _03056_ _03061_ _03063_ VGND VGND VPWR VPWR _03064_ sky130_fd_sc_hd__nor3_1
X_18975_ _09429_ _09430_ VGND VGND VPWR VPWR _09431_ sky130_fd_sc_hd__xnor2_1
X_14098_ _03938_ _03942_ _04069_ VGND VGND VPWR VPWR _04070_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13049_ _02956_ _02958_ VGND VGND VPWR VPWR _02988_ sky130_fd_sc_hd__xnor2_2
X_17926_ _08274_ _08276_ VGND VGND VPWR VPWR _08277_ sky130_fd_sc_hd__and2_1
XFILLER_0_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17857_ _08187_ _08199_ _08200_ VGND VGND VPWR VPWR _08201_ sky130_fd_sc_hd__or3_1
X_16808_ _06936_ _07042_ VGND VGND VPWR VPWR _07047_ sky130_fd_sc_hd__xnor2_2
X_17788_ net298 net295 _02932_ _07570_ VGND VGND VPWR VPWR _08125_ sky130_fd_sc_hd__and4_1
XFILLER_0_49_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16739_ _06947_ _06954_ _06956_ VGND VGND VPWR VPWR _06971_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18409_ _06154_ _08807_ VGND VGND VPWR VPWR _08808_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09975_ _07052_ _07063_ VGND VGND VPWR VPWR _07074_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10750_ _00684_ _00688_ VGND VGND VPWR VPWR _00689_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10681_ _00604_ _00607_ _00610_ VGND VGND VPWR VPWR _00620_ sky130_fd_sc_hd__nor3_1
X_12420_ _02306_ _02344_ _02343_ VGND VGND VPWR VPWR _02359_ sky130_fd_sc_hd__o21a_1
XFILLER_0_152_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12351_ _02194_ _02193_ VGND VGND VPWR VPWR _02290_ sky130_fd_sc_hd__and2b_1
XFILLER_0_50_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11302_ _01236_ _01239_ _01240_ VGND VGND VPWR VPWR _01241_ sky130_fd_sc_hd__a21oi_2
X_15070_ _05123_ _05133_ _05134_ VGND VGND VPWR VPWR _05135_ sky130_fd_sc_hd__nand3_2
X_12282_ _02218_ _02220_ VGND VGND VPWR VPWR _02221_ sky130_fd_sc_hd__xor2_4
XFILLER_0_121_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14021_ net411 net151 net146 net416 VGND VGND VPWR VPWR _03993_ sky130_fd_sc_hd__a22oi_1
X_11233_ _01052_ _01058_ _01057_ VGND VGND VPWR VPWR _01172_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11164_ _00991_ _01012_ _01011_ VGND VGND VPWR VPWR _01103_ sky130_fd_sc_hd__o21a_1
X_10115_ _08559_ _08603_ VGND VGND VPWR VPWR _08614_ sky130_fd_sc_hd__xor2_1
X_18760_ _09086_ _09192_ _09193_ VGND VGND VPWR VPWR _09194_ sky130_fd_sc_hd__a21o_1
X_15972_ _06008_ _06126_ VGND VGND VPWR VPWR _06127_ sky130_fd_sc_hd__and2_2
X_11095_ _01031_ _01033_ VGND VGND VPWR VPWR _01034_ sky130_fd_sc_hd__nor2_1
X_17711_ _08038_ _08039_ VGND VGND VPWR VPWR _08040_ sky130_fd_sc_hd__and2_1
X_14923_ _04807_ _04809_ VGND VGND VPWR VPWR _04974_ sky130_fd_sc_hd__or2_1
X_10046_ net368 net520 _05149_ VGND VGND VPWR VPWR _07855_ sky130_fd_sc_hd__and3_1
X_18691_ _09108_ _09116_ _09117_ VGND VGND VPWR VPWR _09118_ sky130_fd_sc_hd__o21bai_1
X_17642_ _07872_ _07960_ _07959_ _07952_ VGND VGND VPWR VPWR _07964_ sky130_fd_sc_hd__a211oi_1
X_14854_ net465 net485 net139 net122 VGND VGND VPWR VPWR _04898_ sky130_fd_sc_hd__and4_1
X_13805_ _03733_ _03735_ VGND VGND VPWR VPWR _03771_ sky130_fd_sc_hd__xor2_1
X_17573_ net328 _06467_ _07886_ _07887_ VGND VGND VPWR VPWR _07889_ sky130_fd_sc_hd__nand4_2
X_11997_ _01933_ _01934_ _01935_ VGND VGND VPWR VPWR _01936_ sky130_fd_sc_hd__nor3_1
X_14785_ net458 net143 net139 net461 VGND VGND VPWR VPWR _04822_ sky130_fd_sc_hd__a22oi_1
X_19312_ clknet_4_1_0_clock _00013_ VGND VGND VPWR VPWR kd_1\[4\] sky130_fd_sc_hd__dfxtp_1
X_16524_ _06731_ _06734_ VGND VGND VPWR VPWR _06735_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13736_ _03689_ _03679_ _03687_ VGND VGND VPWR VPWR _03702_ sky130_fd_sc_hd__nor3_1
X_10948_ net363 _00243_ VGND VGND VPWR VPWR _00887_ sky130_fd_sc_hd__and2_1
XFILLER_0_156_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19243_ clknet_4_13_0_clock _00125_ VGND VGND VPWR VPWR i_error\[11\] sky130_fd_sc_hd__dfxtp_1
X_16455_ _06555_ _06581_ VGND VGND VPWR VPWR _06659_ sky130_fd_sc_hd__xor2_1
XFILLER_0_155_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13667_ _03449_ _03629_ _03522_ VGND VGND VPWR VPWR _03630_ sky130_fd_sc_hd__a21oi_1
X_10879_ _00815_ VGND VGND VPWR VPWR _00818_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_144_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15406_ _05488_ _05502_ _05503_ _05504_ VGND VGND VPWR VPWR _05505_ sky130_fd_sc_hd__a211o_1
X_12618_ _02556_ _02554_ VGND VGND VPWR VPWR _02557_ sky130_fd_sc_hd__xnor2_1
X_19174_ net502 _09048_ VGND VGND VPWR VPWR _09584_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13598_ net269 net252 _02409_ _01908_ VGND VGND VPWR VPWR _03557_ sky130_fd_sc_hd__and4_1
X_16386_ _06555_ _06556_ VGND VGND VPWR VPWR _06583_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_53_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18125_ _08488_ _08492_ VGND VGND VPWR VPWR _08496_ sky130_fd_sc_hd__and2_1
X_12549_ _02483_ _02487_ VGND VGND VPWR VPWR _02488_ sky130_fd_sc_hd__nand2_1
X_15337_ net427 net432 net198 net193 VGND VGND VPWR VPWR _05429_ sky130_fd_sc_hd__and4_1
XFILLER_0_53_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18056_ _08308_ _08406_ _08410_ VGND VGND VPWR VPWR _08420_ sky130_fd_sc_hd__or3_1
XANTENNA_1 _01698_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15268_ _05250_ _05251_ VGND VGND VPWR VPWR _05353_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17007_ _07263_ _07265_ VGND VGND VPWR VPWR _07266_ sky130_fd_sc_hd__or2_1
X_14219_ _04188_ _04198_ VGND VGND VPWR VPWR _04199_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15199_ _05178_ _05276_ VGND VGND VPWR VPWR _05277_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09760_ net562 _04687_ _04698_ VGND VGND VPWR VPWR _04709_ sky130_fd_sc_hd__o21ai_4
X_18958_ net418 net117 VGND VGND VPWR VPWR _09412_ sky130_fd_sc_hd__nand2_1
X_17909_ _08248_ _08250_ VGND VGND VPWR VPWR _08258_ sky130_fd_sc_hd__nand2_1
X_09691_ net53 _03881_ _03914_ net389 VGND VGND VPWR VPWR _00070_ sky130_fd_sc_hd__a22o_1
X_18889_ _02168_ _02169_ _09332_ _09333_ VGND VGND VPWR VPWR _09336_ sky130_fd_sc_hd__a2bb2o_1
Xrebuffer13 _08751_ VGND VGND VPWR VPWR net572 sky130_fd_sc_hd__clkbuf_1
Xrebuffer24 _08686_ VGND VGND VPWR VPWR net531 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09958_ net361 _05083_ VGND VGND VPWR VPWR _06887_ sky130_fd_sc_hd__and2_1
X_09889_ _05391_ _05952_ _06117_ VGND VGND VPWR VPWR _06128_ sky130_fd_sc_hd__o21ba_1
X_11920_ _01706_ _01858_ VGND VGND VPWR VPWR _01859_ sky130_fd_sc_hd__xnor2_4
X_11851_ net231 _01772_ _01779_ net227 VGND VGND VPWR VPWR _01790_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_68_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10802_ _00726_ _00727_ _00740_ VGND VGND VPWR VPWR _00741_ sky130_fd_sc_hd__o21ai_4
X_14570_ net461 net125 VGND VGND VPWR VPWR _04585_ sky130_fd_sc_hd__nand2_1
X_11782_ _01714_ _00516_ _01715_ _01719_ _01720_ VGND VGND VPWR VPWR _01721_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13521_ _03472_ _03477_ _03479_ VGND VGND VPWR VPWR _03480_ sky130_fd_sc_hd__o21ai_4
X_10733_ _00668_ _00671_ VGND VGND VPWR VPWR _00672_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13452_ _03390_ _03406_ _03388_ VGND VGND VPWR VPWR _03411_ sky130_fd_sc_hd__o21a_1
X_16240_ _06420_ _06421_ VGND VGND VPWR VPWR _06422_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10664_ _00521_ _00602_ VGND VGND VPWR VPWR _00603_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12403_ _02310_ _02340_ VGND VGND VPWR VPWR _02342_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13383_ net199 _03065_ _03335_ VGND VGND VPWR VPWR _03337_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16171_ _06345_ VGND VGND VPWR VPWR _06346_ sky130_fd_sc_hd__clkbuf_4
X_10595_ net383 _05171_ VGND VGND VPWR VPWR _00534_ sky130_fd_sc_hd__nand2_2
XFILLER_0_50_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12334_ _02271_ _02272_ VGND VGND VPWR VPWR _02273_ sky130_fd_sc_hd__and2_1
X_15122_ _05190_ _05191_ VGND VGND VPWR VPWR _05192_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15053_ _05114_ _05115_ VGND VGND VPWR VPWR _05117_ sky130_fd_sc_hd__nor2_1
X_12265_ _02185_ _02174_ VGND VGND VPWR VPWR _02204_ sky130_fd_sc_hd__or2b_1
XPHY_EDGE_ROW_128_Right_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14004_ _03974_ _03975_ VGND VGND VPWR VPWR _03976_ sky130_fd_sc_hd__nor2_1
X_11216_ _01153_ _01154_ VGND VGND VPWR VPWR _01155_ sky130_fd_sc_hd__and2b_1
X_12196_ _01992_ _01993_ _02133_ VGND VGND VPWR VPWR _02135_ sky130_fd_sc_hd__or3_1
X_18812_ net422 net117 VGND VGND VPWR VPWR _09251_ sky130_fd_sc_hd__nand2_1
Xoutput82 net82 VGND VGND VPWR VPWR out_clocked[11] sky130_fd_sc_hd__buf_2
Xoutput93 net93 VGND VGND VPWR VPWR out_clocked[4] sky130_fd_sc_hd__buf_2
X_11147_ net346 _00818_ _01027_ VGND VGND VPWR VPWR _01086_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_50_Left_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18743_ _09173_ _09174_ VGND VGND VPWR VPWR _09176_ sky130_fd_sc_hd__and2b_1
X_15955_ _06048_ _06049_ VGND VGND VPWR VPWR _06109_ sky130_fd_sc_hd__xnor2_1
X_11078_ _01016_ VGND VGND VPWR VPWR _01017_ sky130_fd_sc_hd__inv_2
X_10029_ _07624_ _07646_ VGND VGND VPWR VPWR _07668_ sky130_fd_sc_hd__nor2_1
X_14906_ _04930_ _04954_ VGND VGND VPWR VPWR _04955_ sky130_fd_sc_hd__nand2_1
X_18674_ _08935_ _09075_ _09077_ VGND VGND VPWR VPWR _09100_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_144_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15886_ _03879_ _06032_ VGND VGND VPWR VPWR _06033_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17625_ _07941_ _07916_ _07944_ VGND VGND VPWR VPWR _07946_ sky130_fd_sc_hd__and3_1
X_14837_ _04877_ _04878_ VGND VGND VPWR VPWR _04879_ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17556_ _07820_ _07836_ _07838_ VGND VGND VPWR VPWR _07870_ sky130_fd_sc_hd__and3_1
X_14768_ net481 net121 _04482_ VGND VGND VPWR VPWR _04803_ sky130_fd_sc_hd__and3_1
XFILLER_0_86_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16507_ net272 _06621_ _06624_ VGND VGND VPWR VPWR _06716_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13719_ _03678_ _03673_ _03676_ VGND VGND VPWR VPWR _03685_ sky130_fd_sc_hd__nor3_1
XFILLER_0_156_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17487_ _07782_ _07793_ VGND VGND VPWR VPWR _07794_ sky130_fd_sc_hd__xnor2_2
X_14699_ _04520_ _04726_ VGND VGND VPWR VPWR _04727_ sky130_fd_sc_hd__nor2_1
X_19226_ clknet_4_5_0_clock _00108_ VGND VGND VPWR VPWR prev_error\[13\] sky130_fd_sc_hd__dfxtp_1
X_16438_ _06639_ VGND VGND VPWR VPWR _06640_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19157_ _09559_ _09124_ _09573_ net490 VGND VGND VPWR VPWR _00133_ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16369_ net281 _06311_ VGND VGND VPWR VPWR _06564_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18108_ _08466_ _08476_ VGND VGND VPWR VPWR _08477_ sky130_fd_sc_hd__and2b_1
XFILLER_0_14_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19088_ _09523_ _00325_ _09530_ net489 VGND VGND VPWR VPWR _00100_ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18039_ _08379_ _08397_ _08398_ _08400_ _08357_ VGND VGND VPWR VPWR _08401_ sky130_fd_sc_hd__a32o_1
XFILLER_0_111_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout305 net306 VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__clkbuf_4
Xfanout316 net317 VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout327 net330 VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__buf_2
X_09812_ net6 net64 VGND VGND VPWR VPWR _05281_ sky130_fd_sc_hd__and2b_1
Xfanout338 net339 VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__clkbuf_4
Xfanout349 net350 VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__buf_1
XFILLER_0_94_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09743_ net78 net20 VGND VGND VPWR VPWR _04522_ sky130_fd_sc_hd__or2b_1
XFILLER_0_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09674_ net43 _03614_ _03647_ net290 VGND VGND VPWR VPWR _00041_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10380_ _00249_ _00250_ VGND VGND VPWR VPWR _00319_ sky130_fd_sc_hd__xor2_1
XFILLER_0_20_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_107_Left_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12050_ net223 _01931_ VGND VGND VPWR VPWR _01989_ sky130_fd_sc_hd__or2_1
X_11001_ _00850_ _00851_ VGND VGND VPWR VPWR _00940_ sky130_fd_sc_hd__xor2_2
X_15740_ net469 net473 net196 net192 VGND VGND VPWR VPWR _05872_ sky130_fd_sc_hd__and4_1
X_12952_ _02885_ _02890_ VGND VGND VPWR VPWR _02891_ sky130_fd_sc_hd__nand2_1
X_11903_ _01840_ _01841_ VGND VGND VPWR VPWR _01842_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15671_ _05790_ _05795_ VGND VGND VPWR VPWR _05796_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_116_Left_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12883_ net224 _02090_ VGND VGND VPWR VPWR _02822_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17410_ _07697_ _07698_ _07708_ VGND VGND VPWR VPWR _07709_ sky130_fd_sc_hd__nor3b_1
X_14622_ _04421_ _04641_ VGND VGND VPWR VPWR _04642_ sky130_fd_sc_hd__or2_1
X_11834_ net234 _01772_ _01770_ VGND VGND VPWR VPWR _01773_ sky130_fd_sc_hd__a21oi_1
X_18390_ _08776_ _08786_ VGND VGND VPWR VPWR _08787_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17341_ _07630_ _07631_ _07532_ _07603_ VGND VGND VPWR VPWR _07633_ sky130_fd_sc_hd__a211oi_1
X_14553_ net413 net175 _04565_ VGND VGND VPWR VPWR _04567_ sky130_fd_sc_hd__and3_1
X_11765_ prev_error\[11\] VGND VGND VPWR VPWR _01704_ sky130_fd_sc_hd__inv_4
XFILLER_0_82_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13504_ _03386_ _03408_ _03407_ VGND VGND VPWR VPWR _03463_ sky130_fd_sc_hd__a21o_1
X_10716_ _00625_ _00599_ VGND VGND VPWR VPWR _00655_ sky130_fd_sc_hd__or2b_1
X_17272_ net291 _07156_ VGND VGND VPWR VPWR _07557_ sky130_fd_sc_hd__nand2_1
X_14484_ net458 net129 _04490_ VGND VGND VPWR VPWR _04491_ sky130_fd_sc_hd__a21boi_1
X_11696_ net399 _00615_ VGND VGND VPWR VPWR _01635_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19011_ _09469_ VGND VGND VPWR VPWR _09470_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16223_ _06402_ VGND VGND VPWR VPWR _06404_ sky130_fd_sc_hd__clkbuf_4
X_13435_ _03392_ _03393_ VGND VGND VPWR VPWR _03394_ sky130_fd_sc_hd__nor2_1
X_10647_ _00584_ _00585_ VGND VGND VPWR VPWR _00586_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer4 _09099_ VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13366_ _03242_ _03243_ VGND VGND VPWR VPWR _03319_ sky130_fd_sc_hd__xnor2_2
X_16154_ _06324_ VGND VGND VPWR VPWR _06328_ sky130_fd_sc_hd__buf_2
XFILLER_0_12_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10578_ net337 _00516_ VGND VGND VPWR VPWR _00517_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_125_Left_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15105_ _05172_ _05173_ VGND VGND VPWR VPWR _05174_ sky130_fd_sc_hd__nor2_1
X_12317_ _02252_ _02255_ VGND VGND VPWR VPWR _02256_ sky130_fd_sc_hd__nor2_1
X_16085_ _06180_ _06182_ _06181_ _08570_ VGND VGND VPWR VPWR _06252_ sky130_fd_sc_hd__a2bb2o_1
X_13297_ _03156_ _03158_ _03157_ VGND VGND VPWR VPWR _03250_ sky130_fd_sc_hd__a21o_1
XFILLER_0_139_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12248_ _02178_ _02183_ _02181_ VGND VGND VPWR VPWR _02187_ sky130_fd_sc_hd__o21ai_1
X_15036_ _04955_ _04996_ VGND VGND VPWR VPWR _05098_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12179_ _02030_ _02117_ VGND VGND VPWR VPWR _02118_ sky130_fd_sc_hd__nor2_1
X_16987_ _07224_ _07231_ _07243_ VGND VGND VPWR VPWR _07244_ sky130_fd_sc_hd__or3b_2
XFILLER_0_64_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18726_ _06102_ _06070_ _06101_ VGND VGND VPWR VPWR _09157_ sky130_fd_sc_hd__nand3_1
XFILLER_0_155_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15938_ _05946_ _06081_ _06082_ _03851_ VGND VGND VPWR VPWR _06090_ sky130_fd_sc_hd__o22ai_1
XPHY_EDGE_ROW_134_Left_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18657_ _08919_ _09075_ _09077_ VGND VGND VPWR VPWR _09081_ sky130_fd_sc_hd__nand3_1
X_15869_ _02464_ _03884_ VGND VGND VPWR VPWR _06014_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17608_ _07925_ _07926_ VGND VGND VPWR VPWR _07927_ sky130_fd_sc_hd__nor2_1
X_18588_ _09004_ _09003_ VGND VGND VPWR VPWR _09005_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17539_ net311 _06721_ _07803_ _07850_ VGND VGND VPWR VPWR _07851_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_74_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19209_ clknet_4_15_0_clock _00091_ VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout124 net125 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__buf_2
Xfanout135 net136 VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__buf_2
Xfanout146 kd_2\[11\] VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__buf_2
Xfanout157 net159 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__buf_2
Xfanout168 net169 VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_2
Xfanout179 net180 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__buf_2
X_09726_ net15 net73 VGND VGND VPWR VPWR _04335_ sky130_fd_sc_hd__xnor2_2
X_09657_ _03603_ VGND VGND VPWR VPWR _03614_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11550_ net391 _00323_ _01488_ VGND VGND VPWR VPWR _01489_ sky130_fd_sc_hd__and3_1
X_10501_ net392 VGND VGND VPWR VPWR _00440_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11481_ _01416_ _01419_ VGND VGND VPWR VPWR _01420_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13220_ _03141_ _03172_ VGND VGND VPWR VPWR _03173_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10432_ net375 _05413_ _00279_ VGND VGND VPWR VPWR _00371_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13151_ net239 _02089_ _01907_ net244 VGND VGND VPWR VPWR _03100_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10363_ net384 net539 VGND VGND VPWR VPWR _00302_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12102_ _01780_ _02040_ VGND VGND VPWR VPWR _02041_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13082_ net224 _02331_ _02898_ VGND VGND VPWR VPWR _03024_ sky130_fd_sc_hd__a21oi_1
X_10294_ net356 _05996_ _06183_ net354 VGND VGND VPWR VPWR _00233_ sky130_fd_sc_hd__a22oi_1
X_16910_ net271 _07157_ VGND VGND VPWR VPWR _07159_ sky130_fd_sc_hd__nand2_1
X_12033_ _01777_ _01926_ VGND VGND VPWR VPWR _01972_ sky130_fd_sc_hd__xor2_2
X_17890_ _08235_ _08236_ VGND VGND VPWR VPWR _08237_ sky130_fd_sc_hd__nand2_1
X_16841_ _07004_ _07082_ VGND VGND VPWR VPWR _07083_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16772_ _06921_ _06919_ VGND VGND VPWR VPWR _07007_ sky130_fd_sc_hd__or2_1
X_13984_ net448 net120 VGND VGND VPWR VPWR _03956_ sky130_fd_sc_hd__nand2_1
X_18511_ _08775_ _08918_ _08919_ _08826_ VGND VGND VPWR VPWR _08920_ sky130_fd_sc_hd__a2bb2o_1
X_15723_ _05810_ _05852_ VGND VGND VPWR VPWR _05854_ sky130_fd_sc_hd__nand2_1
X_12935_ _02773_ _02871_ VGND VGND VPWR VPWR _02874_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18442_ _08833_ _08837_ _08841_ _08843_ VGND VGND VPWR VPWR _08844_ sky130_fd_sc_hd__o22a_1
X_15654_ _05771_ _05756_ _05769_ VGND VGND VPWR VPWR _05778_ sky130_fd_sc_hd__and3_1
XFILLER_0_157_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12866_ _02777_ _02792_ VGND VGND VPWR VPWR _02805_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_146_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14605_ _04614_ _04617_ _04619_ VGND VGND VPWR VPWR _04624_ sky130_fd_sc_hd__nor3_1
X_18373_ _08754_ _08755_ _08758_ _08762_ _08764_ VGND VGND VPWR VPWR _08769_ sky130_fd_sc_hd__a32o_1
X_11817_ prev_error\[18\] _05072_ VGND VGND VPWR VPWR _01756_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15585_ _05698_ _05701_ VGND VGND VPWR VPWR _05702_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12797_ _02645_ _02656_ VGND VGND VPWR VPWR _02736_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17324_ _07608_ _07609_ _07612_ VGND VGND VPWR VPWR _07615_ sky130_fd_sc_hd__a21o_1
X_14536_ _04455_ _04547_ VGND VGND VPWR VPWR _04548_ sky130_fd_sc_hd__nand2_1
X_11748_ _01682_ _01686_ _01684_ VGND VGND VPWR VPWR _01687_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17255_ net308 net305 _06467_ _06619_ VGND VGND VPWR VPWR _07539_ sky130_fd_sc_hd__and4_1
X_14467_ _04470_ _04471_ VGND VGND VPWR VPWR _04472_ sky130_fd_sc_hd__or2_1
X_11679_ net394 net390 _00809_ _00814_ VGND VGND VPWR VPWR _01618_ sky130_fd_sc_hd__and4_1
XFILLER_0_70_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16206_ _06383_ _06384_ VGND VGND VPWR VPWR _06385_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13418_ _03374_ _03280_ VGND VGND VPWR VPWR _03375_ sky130_fd_sc_hd__xnor2_1
X_17186_ net316 _06352_ _07462_ VGND VGND VPWR VPWR _07463_ sky130_fd_sc_hd__nand3_1
X_14398_ _04386_ _04388_ _04395_ VGND VGND VPWR VPWR _04396_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16137_ _06307_ _06308_ VGND VGND VPWR VPWR _06309_ sky130_fd_sc_hd__and2_2
X_13349_ _03228_ _03301_ VGND VGND VPWR VPWR _03302_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16068_ _08097_ _05193_ _04896_ net339 VGND VGND VPWR VPWR _06233_ sky130_fd_sc_hd__o211ai_1
X_15019_ _05066_ _05077_ VGND VGND VPWR VPWR _05079_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_142_Left_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18709_ _08775_ _08881_ VGND VGND VPWR VPWR _09138_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09709_ net563 net80 VGND VGND VPWR VPWR _04148_ sky130_fd_sc_hd__and2_1
X_10981_ _00917_ _00919_ VGND VGND VPWR VPWR _00920_ sky130_fd_sc_hd__or2b_1
X_12720_ _02634_ _02657_ VGND VGND VPWR VPWR _02659_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12651_ _02497_ _02498_ VGND VGND VPWR VPWR _02590_ sky130_fd_sc_hd__xor2_1
XFILLER_0_37_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11602_ _01472_ _01518_ VGND VGND VPWR VPWR _01541_ sky130_fd_sc_hd__nor2_1
X_12582_ _02518_ _02488_ _02519_ VGND VGND VPWR VPWR _02521_ sky130_fd_sc_hd__and3_1
X_15370_ _05383_ _05464_ VGND VGND VPWR VPWR _05465_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14321_ _04221_ _04310_ VGND VGND VPWR VPWR _04311_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11533_ net374 _00814_ VGND VGND VPWR VPWR _01472_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17040_ _07279_ _07281_ _07280_ VGND VGND VPWR VPWR _07302_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_135_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14252_ net434 net136 _03963_ _03964_ VGND VGND VPWR VPWR _04235_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_80_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11464_ _01391_ _01396_ VGND VGND VPWR VPWR _01403_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13203_ _03149_ _03154_ _03155_ VGND VGND VPWR VPWR _03156_ sky130_fd_sc_hd__o21ai_2
X_10415_ _00269_ _00353_ VGND VGND VPWR VPWR _00354_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14183_ _04124_ VGND VGND VPWR VPWR _04160_ sky130_fd_sc_hd__inv_2
X_11395_ _01317_ _01330_ VGND VGND VPWR VPWR _01334_ sky130_fd_sc_hd__xor2_1
X_13134_ _03072_ _03053_ VGND VGND VPWR VPWR _03082_ sky130_fd_sc_hd__or2b_1
X_10346_ _00214_ _00216_ VGND VGND VPWR VPWR _00285_ sky130_fd_sc_hd__xor2_1
X_18991_ _09447_ VGND VGND VPWR VPWR _09448_ sky130_fd_sc_hd__buf_6
X_13065_ _02989_ _02584_ VGND VGND VPWR VPWR _03006_ sky130_fd_sc_hd__nor2_1
X_17942_ _08244_ _08253_ _08252_ VGND VGND VPWR VPWR _08294_ sky130_fd_sc_hd__o21ai_1
X_10277_ _09521_ _00215_ VGND VGND VPWR VPWR _00216_ sky130_fd_sc_hd__or2_1
X_12016_ _01884_ _01954_ VGND VGND VPWR VPWR _01955_ sky130_fd_sc_hd__nand2_1
X_17873_ _08210_ _08216_ _08217_ VGND VGND VPWR VPWR _08219_ sky130_fd_sc_hd__or3_1
X_16824_ _06966_ _06968_ VGND VGND VPWR VPWR _07065_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_136_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16755_ net278 _06890_ VGND VGND VPWR VPWR _06989_ sky130_fd_sc_hd__nand2_1
X_13967_ net435 net119 VGND VGND VPWR VPWR _03939_ sky130_fd_sc_hd__nand2_1
X_15706_ net466 net483 net191 net176 VGND VGND VPWR VPWR _05835_ sky130_fd_sc_hd__and4_1
X_12918_ _02752_ _02753_ VGND VGND VPWR VPWR _02857_ sky130_fd_sc_hd__or2_1
X_16686_ _06552_ _06912_ _06542_ VGND VGND VPWR VPWR _06913_ sky130_fd_sc_hd__a21o_1
X_13898_ _03087_ _03864_ VGND VGND VPWR VPWR _03865_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18425_ _08824_ _08825_ VGND VGND VPWR VPWR _08826_ sky130_fd_sc_hd__xnor2_2
X_15637_ _05703_ _05758_ VGND VGND VPWR VPWR _05759_ sky130_fd_sc_hd__xnor2_1
X_12849_ _02686_ _02787_ VGND VGND VPWR VPWR _02788_ sky130_fd_sc_hd__and2b_1
XFILLER_0_152_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18356_ _08611_ _08749_ VGND VGND VPWR VPWR _08750_ sky130_fd_sc_hd__nand2_2
X_15568_ net479 net166 _05636_ _05637_ VGND VGND VPWR VPWR _05683_ sky130_fd_sc_hd__o2bb2a_1
X_17307_ _07588_ _07595_ VGND VGND VPWR VPWR _07596_ sky130_fd_sc_hd__xnor2_1
X_14519_ _04527_ _04528_ net421 net165 VGND VGND VPWR VPWR _04529_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_154_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18287_ _08627_ _08673_ VGND VGND VPWR VPWR _08674_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15499_ _05605_ _05606_ VGND VGND VPWR VPWR _05607_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17238_ net321 net514 _06344_ net323 VGND VGND VPWR VPWR _07520_ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17169_ _07425_ _07443_ VGND VGND VPWR VPWR _07444_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09991_ _07228_ _07239_ VGND VGND VPWR VPWR _07250_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10200_ _09499_ _09521_ VGND VGND VPWR VPWR _09527_ sky130_fd_sc_hd__or2_1
X_11180_ _01114_ _01118_ VGND VGND VPWR VPWR _01119_ sky130_fd_sc_hd__nor2_1
X_10131_ _07140_ _08779_ _07173_ VGND VGND VPWR VPWR _08790_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10062_ _08009_ _07921_ _07954_ VGND VGND VPWR VPWR _08031_ sky130_fd_sc_hd__and3_1
X_14870_ _04913_ _04914_ net436 net173 VGND VGND VPWR VPWR _04915_ sky130_fd_sc_hd__and4bb_1
X_13821_ _03772_ _03775_ _03774_ VGND VGND VPWR VPWR _03787_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16540_ _06745_ _06742_ VGND VGND VPWR VPWR _06752_ sky130_fd_sc_hd__xor2_1
X_13752_ _03705_ _03710_ _03709_ VGND VGND VPWR VPWR _03718_ sky130_fd_sc_hd__o21ai_1
X_10964_ net351 _00515_ VGND VGND VPWR VPWR _00903_ sky130_fd_sc_hd__nand2_1
X_12703_ net204 _02546_ _02410_ net207 VGND VGND VPWR VPWR _02642_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16471_ net308 _06324_ _06319_ net306 VGND VGND VPWR VPWR _06676_ sky130_fd_sc_hd__a22o_1
X_13683_ _03645_ _03646_ VGND VGND VPWR VPWR _03648_ sky130_fd_sc_hd__or2_1
X_10895_ net397 _05292_ _05303_ VGND VGND VPWR VPWR _00834_ sky130_fd_sc_hd__and3_2
X_18210_ _08510_ _08588_ VGND VGND VPWR VPWR _08589_ sky130_fd_sc_hd__xnor2_4
X_15422_ _05519_ _05520_ _05511_ _05515_ VGND VGND VPWR VPWR _05522_ sky130_fd_sc_hd__o211a_1
X_12634_ _02561_ _02572_ VGND VGND VPWR VPWR _02573_ sky130_fd_sc_hd__nand2_1
X_19190_ net498 _09345_ VGND VGND VPWR VPWR _09593_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18141_ _07460_ _08501_ _08510_ _08512_ _08509_ VGND VGND VPWR VPWR _08513_ sky130_fd_sc_hd__a32o_2
X_15353_ _05442_ _05443_ _05445_ VGND VGND VPWR VPWR _05447_ sky130_fd_sc_hd__and3_1
X_12565_ _02490_ _02503_ _02501_ VGND VGND VPWR VPWR _02504_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14304_ _04279_ _04282_ VGND VGND VPWR VPWR _04293_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11516_ _01399_ _01454_ VGND VGND VPWR VPWR _01455_ sky130_fd_sc_hd__nor2_1
X_18072_ _08049_ _08434_ _08435_ _08436_ VGND VGND VPWR VPWR _08437_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_124_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15284_ _05265_ _05283_ _05282_ VGND VGND VPWR VPWR _05371_ sky130_fd_sc_hd__a21o_1
X_12496_ _02430_ _01973_ _02434_ VGND VGND VPWR VPWR _02435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17023_ _07279_ _07282_ VGND VGND VPWR VPWR _07284_ sky130_fd_sc_hd__or2b_1
XFILLER_0_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14235_ _03955_ _03960_ VGND VGND VPWR VPWR _04217_ sky130_fd_sc_hd__xor2_1
XFILLER_0_123_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11447_ _01369_ _01384_ _01385_ VGND VGND VPWR VPWR _01386_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_151_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14166_ _04081_ _04128_ _04140_ VGND VGND VPWR VPWR _04141_ sky130_fd_sc_hd__o21a_1
X_11378_ _01254_ _01262_ VGND VGND VPWR VPWR _01317_ sky130_fd_sc_hd__xnor2_1
X_13117_ _02937_ _03062_ VGND VGND VPWR VPWR _03063_ sky130_fd_sc_hd__and2_1
X_10329_ _00265_ _00267_ VGND VGND VPWR VPWR _00268_ sky130_fd_sc_hd__xor2_4
X_18974_ _09231_ _09239_ _09237_ VGND VGND VPWR VPWR _09430_ sky130_fd_sc_hd__a21o_1
X_14097_ _03943_ _03948_ VGND VGND VPWR VPWR _04069_ sky130_fd_sc_hd__and2b_1
X_13048_ _02969_ _02970_ VGND VGND VPWR VPWR _02987_ sky130_fd_sc_hd__xnor2_2
X_17925_ _08078_ _08275_ VGND VGND VPWR VPWR _08276_ sky130_fd_sc_hd__or2_1
X_17856_ _08070_ _08186_ _08184_ VGND VGND VPWR VPWR _08200_ sky130_fd_sc_hd__a21oi_1
X_16807_ _07044_ _07045_ VGND VGND VPWR VPWR _07046_ sky130_fd_sc_hd__and2_2
X_17787_ _08122_ _08123_ VGND VGND VPWR VPWR _08124_ sky130_fd_sc_hd__xnor2_1
X_14999_ _05044_ _05049_ _05055_ _05056_ VGND VGND VPWR VPWR _05057_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_88_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16738_ _06959_ _06965_ _06969_ VGND VGND VPWR VPWR _06970_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16669_ net271 _06891_ _06893_ VGND VGND VPWR VPWR _06894_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18408_ _06153_ _06145_ VGND VGND VPWR VPWR _08807_ sky130_fd_sc_hd__and2b_1
XFILLER_0_56_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18339_ _08618_ VGND VGND VPWR VPWR _08731_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09974_ net342 _05754_ _07041_ VGND VGND VPWR VPWR _07063_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10680_ net337 _00615_ _00616_ _00618_ VGND VGND VPWR VPWR _00619_ sky130_fd_sc_hd__a31o_1
XFILLER_0_94_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_109_Right_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12350_ net221 _01836_ VGND VGND VPWR VPWR _02289_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11301_ _01232_ _01235_ _01231_ VGND VGND VPWR VPWR _01240_ sky130_fd_sc_hd__o21a_1
XFILLER_0_50_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12281_ _01729_ _02219_ VGND VGND VPWR VPWR _02220_ sky130_fd_sc_hd__nand2_4
XFILLER_0_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14020_ net411 net416 net151 net146 VGND VGND VPWR VPWR _03992_ sky130_fd_sc_hd__and4_1
X_11232_ _01062_ _01077_ VGND VGND VPWR VPWR _01171_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11163_ _01081_ _01100_ _01101_ VGND VGND VPWR VPWR _01102_ sky130_fd_sc_hd__nand3_1
X_10114_ _08581_ _08592_ VGND VGND VPWR VPWR _08603_ sky130_fd_sc_hd__nor2_1
X_15971_ _06013_ _06124_ _06125_ VGND VGND VPWR VPWR _06126_ sky130_fd_sc_hd__a21o_1
X_11094_ _00910_ _01032_ VGND VGND VPWR VPWR _01033_ sky130_fd_sc_hd__nand2_1
X_17710_ _07938_ _08028_ _08037_ VGND VGND VPWR VPWR _08039_ sky130_fd_sc_hd__or3_1
X_10045_ _07833_ _05226_ VGND VGND VPWR VPWR _07844_ sky130_fd_sc_hd__xor2_1
X_14922_ _04969_ _04971_ VGND VGND VPWR VPWR _04972_ sky130_fd_sc_hd__nand2_1
X_18690_ _09114_ _09115_ _09111_ VGND VGND VPWR VPWR _09117_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_117_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17641_ _07962_ VGND VGND VPWR VPWR _07963_ sky130_fd_sc_hd__inv_2
X_14853_ net465 net139 net121 net485 VGND VGND VPWR VPWR _04897_ sky130_fd_sc_hd__a22oi_2
X_13804_ _03768_ _03769_ VGND VGND VPWR VPWR _03770_ sky130_fd_sc_hd__nor2_1
X_17572_ net323 _06618_ _06721_ net319 VGND VGND VPWR VPWR _07887_ sky130_fd_sc_hd__a22o_1
X_14784_ net452 net148 VGND VGND VPWR VPWR _04821_ sky130_fd_sc_hd__nand2_1
X_11996_ _01789_ _01930_ _01788_ _01790_ VGND VGND VPWR VPWR _01935_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_86_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19311_ clknet_4_1_0_clock _00012_ VGND VGND VPWR VPWR kd_1\[3\] sky130_fd_sc_hd__dfxtp_1
X_16523_ _06621_ _06732_ net270 VGND VGND VPWR VPWR _06734_ sky130_fd_sc_hd__and3b_1
X_13735_ _03699_ _03700_ VGND VGND VPWR VPWR _03701_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10947_ _00779_ _00885_ VGND VGND VPWR VPWR _00886_ sky130_fd_sc_hd__xnor2_1
X_19242_ clknet_4_13_0_clock _00124_ VGND VGND VPWR VPWR i_error\[10\] sky130_fd_sc_hd__dfxtp_2
X_16454_ _06654_ _06657_ VGND VGND VPWR VPWR _06658_ sky130_fd_sc_hd__nor2_1
X_13666_ net229 _03220_ VGND VGND VPWR VPWR _03629_ sky130_fd_sc_hd__nand2_1
X_10878_ net343 _00614_ _00816_ VGND VGND VPWR VPWR _00817_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_128_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15405_ _05418_ _05417_ _05401_ VGND VGND VPWR VPWR _05504_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12617_ _02416_ _02533_ VGND VGND VPWR VPWR _02556_ sky130_fd_sc_hd__nand2_1
X_19173_ net502 net449 net490 _09582_ VGND VGND VPWR VPWR _00141_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16385_ _06555_ _06581_ VGND VGND VPWR VPWR _06582_ sky130_fd_sc_hd__or2_1
X_13597_ _03523_ _03555_ VGND VGND VPWR VPWR _03556_ sky130_fd_sc_hd__xor2_1
XFILLER_0_143_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18124_ _08491_ _08494_ VGND VGND VPWR VPWR _08495_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15336_ _05426_ _05427_ VGND VGND VPWR VPWR _05428_ sky130_fd_sc_hd__and2_1
X_12548_ net235 _01836_ _02485_ _02486_ VGND VGND VPWR VPWR _02487_ sky130_fd_sc_hd__a31o_1
XFILLER_0_124_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18055_ _08308_ _08410_ _08413_ _08418_ _08301_ VGND VGND VPWR VPWR _08419_ sky130_fd_sc_hd__a2111o_1
X_15267_ _05330_ _05326_ VGND VGND VPWR VPWR _05352_ sky130_fd_sc_hd__or2b_1
X_12479_ _02398_ _02417_ VGND VGND VPWR VPWR _02418_ sky130_fd_sc_hd__and2b_1
XANTENNA_2 _01851_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17006_ _07158_ _07262_ _07264_ VGND VGND VPWR VPWR _07265_ sky130_fd_sc_hd__o21ai_1
X_14218_ _04196_ _04197_ VGND VGND VPWR VPWR _04198_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15198_ _05175_ _05177_ VGND VGND VPWR VPWR _05276_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14149_ _04084_ _04103_ _04121_ VGND VGND VPWR VPWR _04122_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18957_ _09228_ _09245_ _09247_ VGND VGND VPWR VPWR _09411_ sky130_fd_sc_hd__a21boi_1
X_17908_ net298 _02933_ VGND VGND VPWR VPWR _08257_ sky130_fd_sc_hd__nand2_1
X_09690_ net52 _03881_ _03914_ net391 VGND VGND VPWR VPWR _00069_ sky130_fd_sc_hd__a22o_1
X_18888_ _02168_ _02169_ _09334_ VGND VGND VPWR VPWR _09335_ sky130_fd_sc_hd__or3b_1
X_17839_ _08177_ _08178_ _08180_ VGND VGND VPWR VPWR _08181_ sky130_fd_sc_hd__o21ba_1
Xrebuffer14 net535 VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__clkbuf_1
Xrebuffer25 net531 VGND VGND VPWR VPWR net532 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09957_ _06854_ _06865_ VGND VGND VPWR VPWR _06876_ sky130_fd_sc_hd__and2b_1
X_09888_ _06018_ _06106_ VGND VGND VPWR VPWR _06117_ sky130_fd_sc_hd__xor2_1
X_11850_ net231 net227 _01772_ VGND VGND VPWR VPWR _01789_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10801_ _00728_ _00738_ _00739_ VGND VGND VPWR VPWR _00740_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_138_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11781_ prev_error\[2\] _00613_ VGND VGND VPWR VPWR _01720_ sky130_fd_sc_hd__and2b_1
X_13520_ _03365_ _03478_ VGND VGND VPWR VPWR _03479_ sky130_fd_sc_hd__nor2_1
X_10732_ _00669_ _00670_ VGND VGND VPWR VPWR _00671_ sky130_fd_sc_hd__xor2_2
XFILLER_0_48_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13451_ net104 _03345_ _03386_ _03409_ VGND VGND VPWR VPWR _03410_ sky130_fd_sc_hd__o211a_1
X_10663_ _00520_ _00512_ VGND VGND VPWR VPWR _00602_ sky130_fd_sc_hd__and2b_1
XFILLER_0_153_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12402_ _02310_ _02340_ VGND VGND VPWR VPWR _02341_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16170_ _06344_ VGND VGND VPWR VPWR _06345_ sky130_fd_sc_hd__clkbuf_4
X_10594_ _00437_ _00447_ VGND VGND VPWR VPWR _00533_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_23_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13382_ _03271_ _03334_ VGND VGND VPWR VPWR _03335_ sky130_fd_sc_hd__xor2_1
X_15121_ _05090_ _05189_ _05168_ net538 VGND VGND VPWR VPWR _05191_ sky130_fd_sc_hd__a211oi_1
X_12333_ _01765_ _02258_ VGND VGND VPWR VPWR _02272_ sky130_fd_sc_hd__xor2_1
XFILLER_0_90_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15052_ net467 net484 net148 net131 VGND VGND VPWR VPWR _05115_ sky130_fd_sc_hd__and4_1
X_12264_ _02201_ _02202_ VGND VGND VPWR VPWR _02203_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14003_ net420 net141 _03972_ _03973_ VGND VGND VPWR VPWR _03975_ sky130_fd_sc_hd__o2bb2a_1
X_11215_ net367 _00408_ _00514_ net362 VGND VGND VPWR VPWR _01154_ sky130_fd_sc_hd__a22o_1
X_12195_ _01992_ _01993_ _02133_ VGND VGND VPWR VPWR _02134_ sky130_fd_sc_hd__o21ai_2
X_18811_ _04138_ _04194_ _04128_ VGND VGND VPWR VPWR _09250_ sky130_fd_sc_hd__o21bai_2
Xoutput83 net83 VGND VGND VPWR VPWR out_clocked[12] sky130_fd_sc_hd__buf_2
X_11146_ _01082_ _01084_ VGND VGND VPWR VPWR _01085_ sky130_fd_sc_hd__xor2_1
Xoutput94 net94 VGND VGND VPWR VPWR out_clocked[5] sky130_fd_sc_hd__buf_2
X_15954_ _06060_ _06105_ _06107_ VGND VGND VPWR VPWR _06108_ sky130_fd_sc_hd__a21o_1
X_18742_ _09171_ _09172_ _09168_ VGND VGND VPWR VPWR _09174_ sky130_fd_sc_hd__a21o_1
X_11077_ _01014_ _01015_ VGND VGND VPWR VPWR _01016_ sky130_fd_sc_hd__or2b_1
X_10028_ _07624_ _07646_ VGND VGND VPWR VPWR _07657_ sky130_fd_sc_hd__and2_1
X_14905_ _04947_ _04952_ _04930_ _04953_ VGND VGND VPWR VPWR _04954_ sky130_fd_sc_hd__o211ai_2
X_18673_ _08961_ _08962_ _09096_ _08881_ _09097_ VGND VGND VPWR VPWR _09099_ sky130_fd_sc_hd__a221o_1
X_15885_ _03878_ _02770_ _03876_ VGND VGND VPWR VPWR _06032_ sky130_fd_sc_hd__nand3_1
XFILLER_0_144_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14836_ _04876_ _04868_ _04873_ VGND VGND VPWR VPWR _04878_ sky130_fd_sc_hd__and3_1
X_17624_ _07941_ _07916_ _07944_ VGND VGND VPWR VPWR _07945_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17555_ _07601_ _07867_ _07865_ _07862_ VGND VGND VPWR VPWR _07869_ sky130_fd_sc_hd__o211a_1
X_14767_ net481 net121 _04482_ VGND VGND VPWR VPWR _04802_ sky130_fd_sc_hd__a21oi_1
X_11979_ _01915_ _01917_ VGND VGND VPWR VPWR _01918_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16506_ net284 _06438_ _06714_ _06712_ VGND VGND VPWR VPWR _06715_ sky130_fd_sc_hd__a31o_1
X_13718_ _03682_ _03683_ VGND VGND VPWR VPWR _03684_ sky130_fd_sc_hd__xor2_1
XFILLER_0_73_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17486_ _07784_ _07792_ VGND VGND VPWR VPWR _07793_ sky130_fd_sc_hd__xnor2_1
X_14698_ net436 net156 _04518_ _04519_ VGND VGND VPWR VPWR _04726_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_129_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16437_ _06626_ _06638_ _06636_ VGND VGND VPWR VPWR _06639_ sky130_fd_sc_hd__a21oi_2
X_19225_ clknet_4_5_0_clock _00107_ VGND VGND VPWR VPWR prev_error\[12\] sky130_fd_sc_hd__dfxtp_2
X_13649_ _03573_ _03605_ VGND VGND VPWR VPWR _03610_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19156_ net501 net486 VGND VGND VPWR VPWR _09573_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16368_ _06379_ _06561_ _06562_ VGND VGND VPWR VPWR _06563_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_5_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18107_ _08470_ _08475_ VGND VGND VPWR VPWR _08476_ sky130_fd_sc_hd__nand2_1
X_15319_ _05306_ _05408_ VGND VGND VPWR VPWR _05409_ sky130_fd_sc_hd__nor2_1
X_19087_ net499 prev_error\[5\] VGND VGND VPWR VPWR _09530_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16299_ _06397_ _06450_ _06486_ VGND VGND VPWR VPWR _06487_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_2_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18038_ _08397_ _08399_ VGND VGND VPWR VPWR _08400_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout306 net307 VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__clkbuf_4
X_09811_ _05248_ _05259_ VGND VGND VPWR VPWR _05270_ sky130_fd_sc_hd__nand2_1
Xfanout317 ki\[4\] VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__clkbuf_4
Xfanout328 net330 VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__clkbuf_4
Xfanout339 kp\[17\] VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__clkbuf_4
X_09742_ net20 net78 VGND VGND VPWR VPWR _04511_ sky130_fd_sc_hd__and2b_1
X_09673_ net42 _03614_ _03647_ net291 VGND VGND VPWR VPWR _00040_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11000_ _00924_ _00937_ _00938_ VGND VGND VPWR VPWR _00939_ sky130_fd_sc_hd__a21boi_2
X_12951_ net236 _01909_ _02889_ _02886_ VGND VGND VPWR VPWR _02890_ sky130_fd_sc_hd__a31o_1
X_11902_ net208 _01836_ _01839_ VGND VGND VPWR VPWR _01841_ sky130_fd_sc_hd__a21oi_1
X_15670_ _05557_ _05791_ _05794_ VGND VGND VPWR VPWR _05795_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_59_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12882_ _02818_ _02820_ VGND VGND VPWR VPWR _02821_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14621_ _04418_ _04420_ VGND VGND VPWR VPWR _04641_ sky130_fd_sc_hd__nor2_1
X_11833_ _01764_ VGND VGND VPWR VPWR _01772_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17340_ _07532_ _07603_ _07630_ _07631_ VGND VGND VPWR VPWR _07632_ sky130_fd_sc_hd__o211a_1
X_14552_ net417 net182 VGND VGND VPWR VPWR _04565_ sky130_fd_sc_hd__and2_1
X_11764_ prev_error\[15\] _05193_ VGND VGND VPWR VPWR _01703_ sky130_fd_sc_hd__and2b_1
XFILLER_0_95_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13503_ _03456_ _03444_ _03455_ VGND VGND VPWR VPWR _03462_ sky130_fd_sc_hd__nor3_2
X_17271_ net298 _07093_ VGND VGND VPWR VPWR _07556_ sky130_fd_sc_hd__nand2_1
X_10715_ _00565_ _00653_ VGND VGND VPWR VPWR _00654_ sky130_fd_sc_hd__xnor2_4
X_14483_ net451 net133 VGND VGND VPWR VPWR _04490_ sky130_fd_sc_hd__nand2_1
X_11695_ _01633_ _01632_ VGND VGND VPWR VPWR _01634_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19010_ _09467_ _09468_ VGND VGND VPWR VPWR _09469_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16222_ _06401_ VGND VGND VPWR VPWR _06402_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13434_ net229 _02745_ VGND VGND VPWR VPWR _03393_ sky130_fd_sc_hd__nand2_2
XFILLER_0_64_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10646_ net364 _06623_ _00488_ VGND VGND VPWR VPWR _00585_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer5 _08432_ VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__buf_6
X_16153_ _06320_ _06325_ VGND VGND VPWR VPWR _06327_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13365_ _03315_ _03317_ VGND VGND VPWR VPWR _03318_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10577_ _00515_ VGND VGND VPWR VPWR _00516_ sky130_fd_sc_hd__buf_4
XFILLER_0_24_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15104_ net427 net189 net184 net432 VGND VGND VPWR VPWR _05173_ sky130_fd_sc_hd__a22oi_1
X_12316_ _02251_ _02250_ VGND VGND VPWR VPWR _02255_ sky130_fd_sc_hd__and2b_1
X_16084_ _08845_ _06203_ _06887_ VGND VGND VPWR VPWR _06251_ sky130_fd_sc_hd__o21bai_1
X_13296_ _03246_ _03247_ _03248_ VGND VGND VPWR VPWR _03249_ sky130_fd_sc_hd__nor3_2
XFILLER_0_51_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15035_ _05093_ _05087_ _05096_ VGND VGND VPWR VPWR _05097_ sky130_fd_sc_hd__a21o_1
X_12247_ _02174_ _02185_ VGND VGND VPWR VPWR _02186_ sky130_fd_sc_hd__or2b_1
X_12178_ _02033_ _02112_ _02116_ VGND VGND VPWR VPWR _02117_ sky130_fd_sc_hd__o21a_1
X_11129_ _01067_ _00664_ VGND VGND VPWR VPWR _01068_ sky130_fd_sc_hd__and2_1
X_16986_ _07238_ _07242_ VGND VGND VPWR VPWR _07243_ sky130_fd_sc_hd__xnor2_1
X_18725_ _08925_ _09075_ _09077_ VGND VGND VPWR VPWR _09156_ sky130_fd_sc_hd__nand3b_1
X_15937_ _06086_ _06088_ VGND VGND VPWR VPWR _06089_ sky130_fd_sc_hd__and2_1
X_15868_ _06009_ _06010_ _06012_ VGND VGND VPWR VPWR _06013_ sky130_fd_sc_hd__a21o_1
X_18656_ _09075_ _09077_ _09079_ VGND VGND VPWR VPWR _09080_ sky130_fd_sc_hd__a21o_1
X_14819_ _04016_ net190 VGND VGND VPWR VPWR _04859_ sky130_fd_sc_hd__nor2_1
X_17607_ net295 _07182_ VGND VGND VPWR VPWR _07926_ sky130_fd_sc_hd__nand2_1
X_15799_ _05827_ _05935_ _05936_ _05733_ VGND VGND VPWR VPWR _05937_ sky130_fd_sc_hd__o211a_1
X_18587_ _06121_ _09000_ VGND VGND VPWR VPWR _09004_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17538_ net332 _06408_ _06619_ net315 VGND VGND VPWR VPWR _07850_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_156_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17469_ _07703_ _07706_ VGND VGND VPWR VPWR _07774_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19208_ clknet_4_15_0_clock _00090_ VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19139_ _09559_ _09039_ _09562_ net494 VGND VGND VPWR VPWR _00124_ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout125 net126 VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
Xfanout136 kd_2\[14\] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_4
Xfanout147 kd_2\[11\] VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__buf_2
Xfanout158 net159 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_2
Xfanout169 kd_2\[7\] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_2
X_09725_ net16 net74 VGND VGND VPWR VPWR _04324_ sky130_fd_sc_hd__xnor2_4
X_09656_ _03080_ _03592_ VGND VGND VPWR VPWR _03603_ sky130_fd_sc_hd__and2b_2
XFILLER_0_77_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10500_ net396 VGND VGND VPWR VPWR _00439_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11480_ _01417_ _01418_ VGND VGND VPWR VPWR _01419_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10431_ net375 _05413_ _00279_ VGND VGND VPWR VPWR _00370_ sky130_fd_sc_hd__a21o_1
XFILLER_0_122_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13150_ _03097_ _03098_ VGND VGND VPWR VPWR _03099_ sky130_fd_sc_hd__nand2_1
X_10362_ _07338_ _07371_ VGND VGND VPWR VPWR _00301_ sky130_fd_sc_hd__and2b_1
X_12101_ net234 _01779_ _01770_ VGND VGND VPWR VPWR _02040_ sky130_fd_sc_hd__a21o_1
X_13081_ _03005_ _03021_ _02965_ _03022_ VGND VGND VPWR VPWR _03023_ sky130_fd_sc_hd__o211ai_4
X_10293_ net354 _05996_ _00231_ VGND VGND VPWR VPWR _00232_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12032_ _01969_ _01970_ VGND VGND VPWR VPWR _01971_ sky130_fd_sc_hd__and2_1
XFILLER_0_109_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16840_ _06398_ _06891_ _07003_ VGND VGND VPWR VPWR _07082_ sky130_fd_sc_hd__o21ba_1
X_16771_ _06978_ _07005_ VGND VGND VPWR VPWR _07006_ sky130_fd_sc_hd__xnor2_1
X_13983_ _03915_ _03919_ VGND VGND VPWR VPWR _03955_ sky130_fd_sc_hd__nor2_4
X_15722_ _05806_ _05808_ VGND VGND VPWR VPWR _05852_ sky130_fd_sc_hd__or2_1
X_18510_ _06266_ _08827_ VGND VGND VPWR VPWR _08919_ sky130_fd_sc_hd__or2_1
X_12934_ _02772_ _02872_ VGND VGND VPWR VPWR _02873_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15653_ _05774_ _05775_ VGND VGND VPWR VPWR _05777_ sky130_fd_sc_hd__nand2_1
X_18441_ _08585_ _08842_ VGND VGND VPWR VPWR _08843_ sky130_fd_sc_hd__nand2_2
X_12865_ _02798_ _02803_ VGND VGND VPWR VPWR _02804_ sky130_fd_sc_hd__xor2_2
X_14604_ _04485_ _04622_ VGND VGND VPWR VPWR _04623_ sky130_fd_sc_hd__xnor2_1
X_18372_ _08739_ _08744_ _08751_ _08766_ VGND VGND VPWR VPWR _08767_ sky130_fd_sc_hd__a2bb2o_1
X_11816_ prev_error\[18\] _05061_ VGND VGND VPWR VPWR _01755_ sky130_fd_sc_hd__or2_4
X_15584_ _05624_ _05700_ VGND VGND VPWR VPWR _05701_ sky130_fd_sc_hd__xnor2_1
X_12796_ _02732_ _02734_ VGND VGND VPWR VPWR _02735_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17323_ _07608_ _07609_ _07612_ VGND VGND VPWR VPWR _07614_ sky130_fd_sc_hd__nand3_2
X_14535_ _04450_ _04452_ _04454_ VGND VGND VPWR VPWR _04547_ sky130_fd_sc_hd__or3_1
X_11747_ _01130_ _01133_ VGND VGND VPWR VPWR _01686_ sky130_fd_sc_hd__or2b_1
XFILLER_0_154_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17254_ net302 _06721_ VGND VGND VPWR VPWR _07538_ sky130_fd_sc_hd__nand2_1
X_14466_ _04469_ _04437_ _04466_ VGND VGND VPWR VPWR _04471_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11678_ _01615_ _01616_ VGND VGND VPWR VPWR _01617_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_126_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16205_ _06382_ _06327_ _06331_ VGND VGND VPWR VPWR _06384_ sky130_fd_sc_hd__nand3_1
X_13417_ net237 _02409_ VGND VGND VPWR VPWR _03374_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17185_ net566 _06431_ _06434_ VGND VGND VPWR VPWR _07462_ sky130_fd_sc_hd__and3_2
X_10629_ net387 _00567_ _05512_ _05523_ VGND VGND VPWR VPWR _00568_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14397_ _04393_ _04394_ VGND VGND VPWR VPWR _04395_ sky130_fd_sc_hd__and2_1
X_16136_ _01784_ _06269_ _06306_ VGND VGND VPWR VPWR _06308_ sky130_fd_sc_hd__or3_4
X_13348_ _03225_ _03227_ VGND VGND VPWR VPWR _03301_ sky130_fd_sc_hd__or2_1
X_16067_ net339 _04896_ _05193_ _08097_ VGND VGND VPWR VPWR _06232_ sky130_fd_sc_hd__a211o_1
X_13279_ _03151_ _03153_ VGND VGND VPWR VPWR _03232_ sky130_fd_sc_hd__nor2_1
X_15018_ _05066_ _05077_ VGND VGND VPWR VPWR _05078_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16969_ _07218_ _07223_ VGND VGND VPWR VPWR _07224_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18708_ _09082_ _09083_ _06136_ VGND VGND VPWR VPWR _09137_ sky130_fd_sc_hd__a21o_1
X_18639_ _06109_ _06056_ _06108_ VGND VGND VPWR VPWR _09061_ sky130_fd_sc_hd__nand3_1
XFILLER_0_91_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09708_ _04126_ VGND VGND VPWR VPWR _04137_ sky130_fd_sc_hd__buf_1
XFILLER_0_69_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10980_ _00897_ _00918_ VGND VGND VPWR VPWR _00919_ sky130_fd_sc_hd__xnor2_1
X_09639_ net52 _03358_ _03391_ net258 VGND VGND VPWR VPWR _00012_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12650_ _02587_ _02588_ VGND VGND VPWR VPWR _02589_ sky130_fd_sc_hd__or2b_1
XFILLER_0_78_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11601_ _01526_ _01527_ _01539_ VGND VGND VPWR VPWR _01540_ sky130_fd_sc_hd__nand3_2
XFILLER_0_154_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12581_ _02518_ _02488_ _02519_ VGND VGND VPWR VPWR _02520_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14320_ net448 net123 _04220_ VGND VGND VPWR VPWR _04310_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11532_ net370 _00810_ VGND VGND VPWR VPWR _01471_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14251_ _04231_ _04233_ VGND VGND VPWR VPWR _04234_ sky130_fd_sc_hd__nor2_1
X_11463_ _01393_ _01395_ VGND VGND VPWR VPWR _01402_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13202_ _02994_ _03001_ VGND VGND VPWR VPWR _03155_ sky130_fd_sc_hd__xor2_1
X_10414_ _00271_ _00349_ _00352_ VGND VGND VPWR VPWR _00353_ sky130_fd_sc_hd__o21a_2
X_14182_ _04097_ _04101_ _04156_ _04157_ VGND VGND VPWR VPWR _04158_ sky130_fd_sc_hd__o211ai_4
X_11394_ _01295_ _01332_ VGND VGND VPWR VPWR _01333_ sky130_fd_sc_hd__or2_1
X_13133_ _03076_ _03079_ VGND VGND VPWR VPWR _03081_ sky130_fd_sc_hd__and2b_1
X_10345_ _00282_ _00283_ VGND VGND VPWR VPWR _00284_ sky130_fd_sc_hd__and2b_1
X_18990_ _09446_ _09356_ VGND VGND VPWR VPWR _09447_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_104_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13064_ _02988_ _03004_ VGND VGND VPWR VPWR _03005_ sky130_fd_sc_hd__and2b_1
X_17941_ _08244_ _08252_ _08253_ VGND VGND VPWR VPWR _08293_ sky130_fd_sc_hd__or3_1
X_10276_ net350 _06194_ _09514_ VGND VGND VPWR VPWR _00215_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12015_ _01882_ _01886_ VGND VGND VPWR VPWR _01954_ sky130_fd_sc_hd__or2b_1
X_17872_ _08133_ _08215_ _08214_ _08204_ VGND VGND VPWR VPWR _08217_ sky130_fd_sc_hd__o211a_1
X_16823_ _07061_ _07062_ VGND VGND VPWR VPWR _07064_ sky130_fd_sc_hd__nand2_1
X_16754_ _06984_ _06987_ VGND VGND VPWR VPWR _06988_ sky130_fd_sc_hd__xnor2_1
X_13966_ net435 net123 _03924_ _03923_ net119 VGND VGND VPWR VPWR _03938_ sky130_fd_sc_hd__a32o_1
Xmax_cap3 _07692_ VGND VGND VPWR VPWR net537 sky130_fd_sc_hd__buf_1
X_15705_ net462 net195 VGND VGND VPWR VPWR _05834_ sky130_fd_sc_hd__nand2_1
X_12917_ _02853_ _02855_ VGND VGND VPWR VPWR _02856_ sky130_fd_sc_hd__nand2_1
X_16685_ _06545_ _06911_ VGND VGND VPWR VPWR _06912_ sky130_fd_sc_hd__xnor2_1
X_13897_ _02985_ _03086_ VGND VGND VPWR VPWR _03864_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18424_ _08542_ _08578_ VGND VGND VPWR VPWR _08825_ sky130_fd_sc_hd__and2b_1
XFILLER_0_152_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15636_ _05705_ _05704_ VGND VGND VPWR VPWR _05758_ sky130_fd_sc_hd__nor2_1
X_12848_ net259 _01798_ _02684_ _02685_ VGND VGND VPWR VPWR _02787_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15567_ _05680_ _05681_ net478 net171 VGND VGND VPWR VPWR _05682_ sky130_fd_sc_hd__and4bb_1
X_18355_ _08610_ _08536_ _08608_ _08609_ VGND VGND VPWR VPWR _08749_ sky130_fd_sc_hd__or4_1
X_12779_ _02716_ _02717_ VGND VGND VPWR VPWR _02718_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14518_ net429 net161 net155 net567 VGND VGND VPWR VPWR _04528_ sky130_fd_sc_hd__a22oi_1
X_17306_ _07593_ _07594_ VGND VGND VPWR VPWR _07595_ sky130_fd_sc_hd__nor2_1
X_15498_ _05526_ _05549_ _05604_ VGND VGND VPWR VPWR _05606_ sky130_fd_sc_hd__a21oi_1
X_18286_ _08671_ _08672_ VGND VGND VPWR VPWR _08673_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14449_ _04450_ _04451_ net409 net175 VGND VGND VPWR VPWR _04452_ sky130_fd_sc_hd__and4bb_1
X_17237_ net323 net319 _06408_ _06344_ VGND VGND VPWR VPWR _07519_ sky130_fd_sc_hd__nand4_2
XFILLER_0_25_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17168_ _07428_ _07442_ VGND VGND VPWR VPWR _07443_ sky130_fd_sc_hd__xor2_2
XFILLER_0_4_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16119_ _06273_ _02087_ _06287_ _06288_ VGND VGND VPWR VPWR _06289_ sky130_fd_sc_hd__and4_1
X_09990_ _07206_ _07217_ VGND VGND VPWR VPWR _07239_ sky130_fd_sc_hd__nand2_1
X_17099_ _07335_ _07341_ VGND VGND VPWR VPWR _07367_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10130_ _07151_ VGND VGND VPWR VPWR _08779_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10061_ _07921_ _07954_ _08009_ VGND VGND VPWR VPWR _08020_ sky130_fd_sc_hd__a21oi_2
X_13820_ _03752_ _03784_ VGND VGND VPWR VPWR _03786_ sky130_fd_sc_hd__xnor2_1
X_13751_ _03714_ _03716_ VGND VGND VPWR VPWR _03717_ sky130_fd_sc_hd__nor2_1
X_10963_ net357 net351 _00798_ _00515_ VGND VGND VPWR VPWR _00902_ sky130_fd_sc_hd__and4_1
XFILLER_0_98_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12702_ _02640_ VGND VGND VPWR VPWR _02641_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16470_ _06365_ _06674_ VGND VGND VPWR VPWR _06675_ sky130_fd_sc_hd__and2_1
X_13682_ _03635_ _03642_ VGND VGND VPWR VPWR _03646_ sky130_fd_sc_hd__xnor2_1
X_10894_ _00734_ _00735_ VGND VGND VPWR VPWR _00833_ sky130_fd_sc_hd__xnor2_1
X_15421_ _05511_ _05515_ _05519_ _05520_ VGND VGND VPWR VPWR _05521_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_128_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12633_ _02559_ _02560_ VGND VGND VPWR VPWR _02572_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15352_ _05444_ _05419_ VGND VGND VPWR VPWR _05445_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18140_ _08502_ _08511_ VGND VGND VPWR VPWR _08512_ sky130_fd_sc_hd__nand2_1
X_12564_ _02501_ _02502_ VGND VGND VPWR VPWR _02503_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14303_ _04289_ _04290_ VGND VGND VPWR VPWR _04292_ sky130_fd_sc_hd__or2_1
X_11515_ _01397_ _01398_ VGND VGND VPWR VPWR _01454_ sky130_fd_sc_hd__and2_1
X_18071_ _07969_ _07977_ VGND VGND VPWR VPWR _08436_ sky130_fd_sc_hd__nand2_1
X_15283_ _05365_ _05366_ _05368_ VGND VGND VPWR VPWR _05370_ sky130_fd_sc_hd__or3_1
X_12495_ net259 net254 _01764_ _01974_ VGND VGND VPWR VPWR _02434_ sky130_fd_sc_hd__o211a_1
X_17022_ _07280_ _07279_ _07281_ VGND VGND VPWR VPWR _07282_ sky130_fd_sc_hd__or3_1
X_14234_ _04213_ _04215_ VGND VGND VPWR VPWR _04216_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11446_ _01371_ _01383_ VGND VGND VPWR VPWR _01385_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14165_ _04129_ _04139_ VGND VGND VPWR VPWR _04140_ sky130_fd_sc_hd__xor2_1
X_11377_ _01270_ _01269_ _01248_ VGND VGND VPWR VPWR _01316_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_22_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13116_ net202 _02935_ _02927_ _02936_ VGND VGND VPWR VPWR _03062_ sky130_fd_sc_hd__a22o_1
X_10328_ _00182_ _00266_ VGND VGND VPWR VPWR _00267_ sky130_fd_sc_hd__nor2_2
X_18973_ net407 net127 VGND VGND VPWR VPWR _09429_ sky130_fd_sc_hd__nand2_1
X_14096_ _04065_ _04066_ _04035_ _04046_ VGND VGND VPWR VPWR _04068_ sky130_fd_sc_hd__a211oi_1
X_13047_ _02977_ _02979_ VGND VGND VPWR VPWR _02986_ sky130_fd_sc_hd__xnor2_1
X_17924_ net331 _07181_ VGND VGND VPWR VPWR _08275_ sky130_fd_sc_hd__nand2_1
X_10259_ _07778_ _00197_ _07349_ VGND VGND VPWR VPWR _00198_ sky130_fd_sc_hd__o21ai_1
X_17855_ _08193_ _08198_ VGND VGND VPWR VPWR _08199_ sky130_fd_sc_hd__xnor2_1
X_16806_ _06935_ _07043_ VGND VGND VPWR VPWR _07045_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17786_ _07926_ _08018_ _08017_ VGND VGND VPWR VPWR _08123_ sky130_fd_sc_hd__o21a_1
X_14998_ _05051_ _05052_ _05054_ VGND VGND VPWR VPWR _05056_ sky130_fd_sc_hd__nand3_1
XFILLER_0_72_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16737_ _06966_ _06968_ VGND VGND VPWR VPWR _06969_ sky130_fd_sc_hd__and2_1
X_13949_ _03916_ _03920_ VGND VGND VPWR VPWR _03921_ sky130_fd_sc_hd__nor2_2
XFILLER_0_72_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16668_ _06888_ _06892_ VGND VGND VPWR VPWR _06893_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18407_ _08803_ net571 _08800_ VGND VGND VPWR VPWR _08806_ sky130_fd_sc_hd__o21a_1
XFILLER_0_119_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15619_ net469 net183 net179 net473 VGND VGND VPWR VPWR _05739_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_9_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16599_ _06815_ _06812_ VGND VGND VPWR VPWR _06817_ sky130_fd_sc_hd__and2b_1
XFILLER_0_57_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18338_ _08728_ _08729_ VGND VGND VPWR VPWR _08730_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18269_ _06554_ _06572_ _06549_ VGND VGND VPWR VPWR _08654_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_72_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout5 _04995_ VGND VGND VPWR VPWR net539 sky130_fd_sc_hd__clkbuf_4
X_09973_ net342 _05754_ _07041_ VGND VGND VPWR VPWR _07052_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11300_ _01237_ _01106_ _01238_ VGND VGND VPWR VPWR _01239_ sky130_fd_sc_hd__o21a_1
X_12280_ prev_error\[7\] _00226_ VGND VGND VPWR VPWR _02219_ sky130_fd_sc_hd__or2_1
X_11231_ _01104_ _01105_ _01121_ VGND VGND VPWR VPWR _01170_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_121_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11162_ _01079_ _01080_ _01061_ _01078_ VGND VGND VPWR VPWR _01101_ sky130_fd_sc_hd__o211ai_4
X_10113_ net342 _05182_ _08570_ VGND VGND VPWR VPWR _08592_ sky130_fd_sc_hd__and3_1
X_15970_ _06009_ _06010_ _06012_ VGND VGND VPWR VPWR _06125_ sky130_fd_sc_hd__and3_1
X_11093_ _00913_ VGND VGND VPWR VPWR _01032_ sky130_fd_sc_hd__inv_2
X_10044_ net360 _05182_ VGND VGND VPWR VPWR _07833_ sky130_fd_sc_hd__nand2_1
X_14921_ _04967_ _04970_ VGND VGND VPWR VPWR _04971_ sky130_fd_sc_hd__and2_1
Xhold50 i_error\[9\] VGND VGND VPWR VPWR net557 sky130_fd_sc_hd__dlygate4sd3_1
X_17640_ _07955_ _07956_ VGND VGND VPWR VPWR _07962_ sky130_fd_sc_hd__nor2_1
X_14852_ _04890_ _04889_ VGND VGND VPWR VPWR _04895_ sky130_fd_sc_hd__xor2_1
XFILLER_0_89_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13803_ _03760_ _03765_ VGND VGND VPWR VPWR _03769_ sky130_fd_sc_hd__xnor2_1
X_14783_ net461 net143 VGND VGND VPWR VPWR _04820_ sky130_fd_sc_hd__nand2_1
X_17571_ net319 _06618_ _07885_ VGND VGND VPWR VPWR _07886_ sky130_fd_sc_hd__nand3_2
X_11995_ net223 _01932_ _01930_ VGND VGND VPWR VPWR _01934_ sky130_fd_sc_hd__and3_1
X_19310_ clknet_4_1_0_clock _00011_ VGND VGND VPWR VPWR kd_1\[2\] sky130_fd_sc_hd__dfxtp_1
X_16522_ _06710_ _06730_ VGND VGND VPWR VPWR _06732_ sky130_fd_sc_hd__xnor2_1
X_13734_ _03697_ _03698_ VGND VGND VPWR VPWR _03700_ sky130_fd_sc_hd__or2_1
X_10946_ _00782_ _00780_ VGND VGND VPWR VPWR _00885_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19241_ clknet_4_13_0_clock _00123_ VGND VGND VPWR VPWR i_error\[9\] sky130_fd_sc_hd__dfxtp_1
X_13665_ _03622_ _03627_ _03620_ VGND VGND VPWR VPWR _03628_ sky130_fd_sc_hd__o21ai_1
X_16453_ _06653_ _06655_ VGND VGND VPWR VPWR _06657_ sky130_fd_sc_hd__or2_1
X_10877_ net340 _00815_ VGND VGND VPWR VPWR _00816_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12616_ _01847_ _02410_ VGND VGND VPWR VPWR _02555_ sky130_fd_sc_hd__nor2_1
X_15404_ _05418_ _05401_ _05417_ VGND VGND VPWR VPWR _05503_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19172_ net502 _09062_ VGND VGND VPWR VPWR _09582_ sky130_fd_sc_hd__nand2_1
X_16384_ _06361_ _06395_ VGND VGND VPWR VPWR _06581_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13596_ _03547_ _03546_ VGND VGND VPWR VPWR _03555_ sky130_fd_sc_hd__and2_1
XFILLER_0_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15335_ _05425_ _05420_ _05422_ VGND VGND VPWR VPWR _05427_ sky130_fd_sc_hd__or3_1
X_18123_ _08488_ _08492_ VGND VGND VPWR VPWR _08494_ sky130_fd_sc_hd__xnor2_2
X_12547_ _02372_ _02484_ VGND VGND VPWR VPWR _02486_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15266_ _05230_ _05322_ _05323_ VGND VGND VPWR VPWR _05351_ sky130_fd_sc_hd__or3_1
X_18054_ _08265_ _08300_ VGND VGND VPWR VPWR _08418_ sky130_fd_sc_hd__and2_1
X_12478_ _02401_ _02403_ _02416_ VGND VGND VPWR VPWR _02417_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_151_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_3 _02638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14217_ _04195_ _04129_ VGND VGND VPWR VPWR _04197_ sky130_fd_sc_hd__and2b_1
X_17005_ net284 _07095_ _07157_ net278 VGND VGND VPWR VPWR _07264_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11429_ net370 _00615_ _01366_ _01367_ VGND VGND VPWR VPWR _01368_ sky130_fd_sc_hd__a31o_1
X_15197_ net419 net198 _05274_ VGND VGND VPWR VPWR _05275_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14148_ _04104_ _04120_ VGND VGND VPWR VPWR _04121_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14079_ _04049_ _04050_ net408 net144 VGND VGND VPWR VPWR _04051_ sky130_fd_sc_hd__and4b_1
X_18956_ _09247_ _09248_ _09261_ _09260_ VGND VGND VPWR VPWR _09410_ sky130_fd_sc_hd__a31oi_1
X_17907_ _08244_ _08254_ _08201_ _08255_ VGND VGND VPWR VPWR _08256_ sky130_fd_sc_hd__o211a_1
X_18887_ _09332_ _09333_ VGND VGND VPWR VPWR _09334_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17838_ net326 _06889_ _08179_ VGND VGND VPWR VPWR _08180_ sky130_fd_sc_hd__and3_1
Xrebuffer26 _01690_ VGND VGND VPWR VPWR net533 sky130_fd_sc_hd__dlygate4sd1_1
X_17769_ _07991_ _08102_ _08103_ VGND VGND VPWR VPWR _08104_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09956_ net348 _05193_ _06821_ _06843_ VGND VGND VPWR VPWR _06865_ sky130_fd_sc_hd__a22o_1
X_09887_ _06084_ _06095_ VGND VGND VPWR VPWR _06106_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_142_Right_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10800_ _00731_ _00737_ VGND VGND VPWR VPWR _00739_ sky130_fd_sc_hd__nor2_1
X_11780_ _01716_ _01717_ _01718_ VGND VGND VPWR VPWR _01719_ sky130_fd_sc_hd__a21o_2
XFILLER_0_68_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10731_ _00573_ _00572_ VGND VGND VPWR VPWR _00670_ sky130_fd_sc_hd__and2b_1
XFILLER_0_138_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13450_ _03407_ _03386_ _03408_ VGND VGND VPWR VPWR _03409_ sky130_fd_sc_hd__nand3_2
XFILLER_0_94_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10662_ net568 _00600_ VGND VGND VPWR VPWR _00601_ sky130_fd_sc_hd__nand2_2
XFILLER_0_35_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12401_ net199 _02311_ _02338_ _02339_ VGND VGND VPWR VPWR _02340_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_63_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13381_ _03272_ _03331_ _03333_ VGND VGND VPWR VPWR _03334_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_106_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10593_ _00474_ _00479_ VGND VGND VPWR VPWR _00532_ sky130_fd_sc_hd__xor2_4
X_15120_ _05168_ net538 _05090_ _05189_ VGND VGND VPWR VPWR _05190_ sky130_fd_sc_hd__o211a_1
X_12332_ _01975_ _01980_ VGND VGND VPWR VPWR _02271_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15051_ net467 net148 net130 net484 VGND VGND VPWR VPWR _05114_ sky130_fd_sc_hd__a22oi_2
X_12263_ _02191_ _02200_ VGND VGND VPWR VPWR _02202_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14002_ _03972_ _03973_ net420 net141 VGND VGND VPWR VPWR _03974_ sky130_fd_sc_hd__and4bb_1
X_11214_ net366 net362 _00408_ _00514_ VGND VGND VPWR VPWR _01153_ sky130_fd_sc_hd__and4_1
X_12194_ _02131_ _02132_ VGND VGND VPWR VPWR _02133_ sky130_fd_sc_hd__and2_1
X_18810_ _09247_ _09248_ VGND VGND VPWR VPWR _09249_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11145_ _01009_ _01083_ VGND VGND VPWR VPWR _01084_ sky130_fd_sc_hd__nand2_1
Xoutput84 net84 VGND VGND VPWR VPWR out_clocked[13] sky130_fd_sc_hd__buf_2
Xoutput95 net95 VGND VGND VPWR VPWR out_clocked[6] sky130_fd_sc_hd__buf_2
X_18741_ _09168_ _09171_ _09172_ VGND VGND VPWR VPWR _09173_ sky130_fd_sc_hd__and3_1
X_15953_ _06053_ _06055_ VGND VGND VPWR VPWR _06107_ sky130_fd_sc_hd__xnor2_1
X_11076_ _00943_ _00944_ VGND VGND VPWR VPWR _01015_ sky130_fd_sc_hd__xor2_2
X_10027_ _07393_ _07635_ _07360_ VGND VGND VPWR VPWR _07646_ sky130_fd_sc_hd__o21ai_1
X_14904_ _04912_ _04927_ _04928_ VGND VGND VPWR VPWR _04953_ sky130_fd_sc_hd__nand3_1
X_18672_ _08799_ _08881_ VGND VGND VPWR VPWR _09097_ sky130_fd_sc_hd__nor2_1
X_15884_ _05993_ _06030_ VGND VGND VPWR VPWR _06031_ sky130_fd_sc_hd__nor2_1
X_17623_ _07831_ _07942_ VGND VGND VPWR VPWR _07944_ sky130_fd_sc_hd__or2_1
X_14835_ _04868_ _04873_ _04876_ VGND VGND VPWR VPWR _04877_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17554_ _07862_ _07865_ _07867_ _07601_ VGND VGND VPWR VPWR _07868_ sky130_fd_sc_hd__a211oi_2
X_11978_ _01903_ _01916_ VGND VGND VPWR VPWR _01917_ sky130_fd_sc_hd__and2_1
X_14766_ net467 net135 VGND VGND VPWR VPWR _04801_ sky130_fd_sc_hd__nand2_1
X_16505_ _06712_ _06713_ VGND VGND VPWR VPWR _06714_ sky130_fd_sc_hd__nor2_1
X_13717_ net247 _02746_ VGND VGND VPWR VPWR _03683_ sky130_fd_sc_hd__nand2_1
X_10929_ _00861_ _00859_ VGND VGND VPWR VPWR _00868_ sky130_fd_sc_hd__xor2_1
X_14697_ _04722_ _04724_ VGND VGND VPWR VPWR _04725_ sky130_fd_sc_hd__nor2_1
X_17485_ _07790_ _07791_ VGND VGND VPWR VPWR _07792_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19224_ clknet_4_5_0_clock _00106_ VGND VGND VPWR VPWR prev_error\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16436_ _06636_ _06637_ VGND VGND VPWR VPWR _06638_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13648_ _03554_ _03608_ _03550_ VGND VGND VPWR VPWR _03609_ sky130_fd_sc_hd__or3_1
XFILLER_0_144_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19155_ net505 net547 net495 _09572_ VGND VGND VPWR VPWR _00132_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13579_ _03526_ _03535_ VGND VGND VPWR VPWR _03538_ sky130_fd_sc_hd__nor2_1
X_16367_ net290 _06328_ _06379_ net287 VGND VGND VPWR VPWR _06562_ sky130_fd_sc_hd__a22o_1
X_18106_ _08470_ _08473_ _08474_ VGND VGND VPWR VPWR _08475_ sky130_fd_sc_hd__nand3_1
X_15318_ net482 net149 _05304_ _05305_ VGND VGND VPWR VPWR _05408_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_41_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19086_ _09523_ _00410_ _09529_ net489 VGND VGND VPWR VPWR _00099_ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16298_ _06451_ _06485_ VGND VGND VPWR VPWR _06486_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18037_ net322 _08275_ _08395_ _03065_ _07291_ VGND VGND VPWR VPWR _08399_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15249_ _05320_ _05309_ _05318_ VGND VGND VPWR VPWR _05332_ sky130_fd_sc_hd__nand3_1
XFILLER_0_78_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09810_ _05237_ _05116_ VGND VGND VPWR VPWR _05259_ sky130_fd_sc_hd__or2b_1
Xfanout307 ki\[7\] VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__clkbuf_4
Xfanout318 net321 VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__buf_2
Xfanout329 net330 VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__buf_2
X_09741_ _04390_ _04357_ _04478_ _04489_ VGND VGND VPWR VPWR _04500_ sky130_fd_sc_hd__a31o_2
XFILLER_0_94_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18939_ net206 _01930_ VGND VGND VPWR VPWR _09391_ sky130_fd_sc_hd__nand2_1
X_09672_ net41 _03614_ _03647_ net295 VGND VGND VPWR VPWR _00039_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09939_ _06568_ _06667_ VGND VGND VPWR VPWR _06678_ sky130_fd_sc_hd__or2_1
X_12950_ _02886_ _02888_ VGND VGND VPWR VPWR _02889_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11901_ net208 _01836_ _01839_ VGND VGND VPWR VPWR _01840_ sky130_fd_sc_hd__and3_1
X_12881_ _02817_ _02819_ VGND VGND VPWR VPWR _02820_ sky130_fd_sc_hd__or2b_1
X_14620_ _04593_ _04592_ VGND VGND VPWR VPWR _04640_ sky130_fd_sc_hd__or2b_1
X_11832_ net234 _01770_ VGND VGND VPWR VPWR _01771_ sky130_fd_sc_hd__and2_1
X_14551_ _04559_ _04561_ _04563_ VGND VGND VPWR VPWR _04564_ sky130_fd_sc_hd__o21ai_1
X_11763_ _01701_ _04874_ VGND VGND VPWR VPWR _01702_ sky130_fd_sc_hd__nand2_2
XFILLER_0_56_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13502_ _03459_ _03460_ VGND VGND VPWR VPWR _03461_ sky130_fd_sc_hd__nand2_1
X_10714_ _00626_ _00652_ _00650_ VGND VGND VPWR VPWR _00653_ sky130_fd_sc_hd__a21oi_4
X_14482_ net452 net456 net133 net129 VGND VGND VPWR VPWR _04488_ sky130_fd_sc_hd__and4_1
X_17270_ _07553_ _07554_ VGND VGND VPWR VPWR _07555_ sky130_fd_sc_hd__or2_1
X_11694_ _01606_ _01613_ VGND VGND VPWR VPWR _01633_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13433_ net232 _02639_ VGND VGND VPWR VPWR _03392_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16221_ _06400_ VGND VGND VPWR VPWR _06401_ sky130_fd_sc_hd__buf_4
X_10645_ net364 _06623_ _00488_ VGND VGND VPWR VPWR _00584_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16152_ net299 net296 _06324_ VGND VGND VPWR VPWR _06325_ sky130_fd_sc_hd__and3_1
X_13364_ _03313_ _03316_ VGND VGND VPWR VPWR _03317_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10576_ _00514_ VGND VGND VPWR VPWR _00515_ sky130_fd_sc_hd__buf_4
Xrebuffer6 net512 VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__clkbuf_1
X_12315_ _02118_ _02253_ VGND VGND VPWR VPWR _02254_ sky130_fd_sc_hd__nor2_1
X_15103_ net427 net432 net189 net184 VGND VGND VPWR VPWR _05172_ sky130_fd_sc_hd__and4_1
X_16083_ _06245_ _06248_ VGND VGND VPWR VPWR _06250_ sky130_fd_sc_hd__xnor2_1
X_13295_ _03186_ _03197_ VGND VGND VPWR VPWR _03248_ sky130_fd_sc_hd__xnor2_1
X_15034_ _05092_ _05095_ VGND VGND VPWR VPWR _05096_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_2_Left_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12246_ _02011_ _02184_ _01978_ VGND VGND VPWR VPWR _02185_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_39_Left_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12177_ _02113_ _02115_ VGND VGND VPWR VPWR _02116_ sky130_fd_sc_hd__or2b_1
X_11128_ net405 _05897_ _06150_ VGND VGND VPWR VPWR _01067_ sky130_fd_sc_hd__and3_1
X_16985_ _07240_ _07241_ VGND VGND VPWR VPWR _07242_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18724_ _08961_ _08962_ _08788_ _08881_ _09154_ VGND VGND VPWR VPWR _09155_ sky130_fd_sc_hd__a221o_1
X_15936_ _05943_ _06087_ VGND VGND VPWR VPWR _06088_ sky130_fd_sc_hd__nor2_2
X_11059_ _00996_ _00997_ VGND VGND VPWR VPWR _00998_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18655_ _08826_ _09078_ _08880_ VGND VGND VPWR VPWR _09079_ sky130_fd_sc_hd__mux2_1
X_15867_ _03889_ _06011_ VGND VGND VPWR VPWR _06012_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17606_ net298 _07156_ VGND VGND VPWR VPWR _07925_ sky130_fd_sc_hd__nand2_1
X_14818_ _04856_ _04857_ VGND VGND VPWR VPWR _04858_ sky130_fd_sc_hd__nand2_1
X_18586_ _08898_ _09002_ _08964_ VGND VGND VPWR VPWR _09003_ sky130_fd_sc_hd__mux2_2
XFILLER_0_148_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15798_ _05676_ _05731_ _05825_ _05826_ VGND VGND VPWR VPWR _05936_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_59_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17537_ _07803_ _07802_ net311 _06721_ VGND VGND VPWR VPWR _07849_ sky130_fd_sc_hd__and4b_1
XFILLER_0_157_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14749_ _04780_ _04781_ VGND VGND VPWR VPWR _04782_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17468_ _07257_ _07724_ _07725_ _07721_ VGND VGND VPWR VPWR _07773_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_6_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19207_ clknet_4_15_0_clock _00089_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dfxtp_1
X_16419_ _06618_ VGND VGND VPWR VPWR _06619_ sky130_fd_sc_hd__buf_2
XFILLER_0_42_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17399_ _07308_ _07695_ _07696_ VGND VGND VPWR VPWR _07697_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19138_ net504 i_error\[10\] VGND VGND VPWR VPWR _09562_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19069_ _09515_ _09518_ VGND VGND VPWR VPWR _00091_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout126 net127 VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_2
Xfanout137 kd_2\[13\] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_4
Xfanout148 net150 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_4
Xfanout159 kd_2\[9\] VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_2
X_09724_ _04225_ _04269_ _04291_ _04302_ net13 VGND VGND VPWR VPWR _04313_ sky130_fd_sc_hd__o32a_4
X_09655_ net31 _03047_ VGND VGND VPWR VPWR _03592_ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10430_ _00361_ _00368_ VGND VGND VPWR VPWR _00369_ sky130_fd_sc_hd__or2b_1
XFILLER_0_150_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10361_ _07778_ _00197_ VGND VGND VPWR VPWR _00300_ sky130_fd_sc_hd__xor2_1
XFILLER_0_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12100_ _02036_ _02037_ _02038_ VGND VGND VPWR VPWR _02039_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_103_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13080_ _02961_ _02964_ _02963_ VGND VGND VPWR VPWR _03022_ sky130_fd_sc_hd__a21o_1
X_10292_ net357 _05897_ _06150_ VGND VGND VPWR VPWR _00231_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12031_ _01967_ _01968_ VGND VGND VPWR VPWR _01970_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16770_ _06896_ _06979_ _07001_ _07004_ VGND VGND VPWR VPWR _07005_ sky130_fd_sc_hd__a31oi_4
X_13982_ _03921_ _03953_ VGND VGND VPWR VPWR _03954_ sky130_fd_sc_hd__xor2_1
X_15721_ _05848_ _05850_ VGND VGND VPWR VPWR _05851_ sky130_fd_sc_hd__or2b_1
X_12933_ _02773_ _02871_ VGND VGND VPWR VPWR _02872_ sky130_fd_sc_hd__nor2_1
X_18440_ _08542_ _08579_ _08583_ _08584_ VGND VGND VPWR VPWR _08842_ sky130_fd_sc_hd__o22ai_1
X_15652_ net447 net195 _05760_ _05764_ VGND VGND VPWR VPWR _05775_ sky130_fd_sc_hd__a211o_1
X_12864_ _02598_ _02799_ _02802_ VGND VGND VPWR VPWR _02803_ sky130_fd_sc_hd__o21ba_1
X_14603_ net461 net129 VGND VGND VPWR VPWR _04622_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18371_ _08750_ _08748_ _08759_ _08765_ VGND VGND VPWR VPWR _08766_ sky130_fd_sc_hd__a211o_1
X_11815_ _01700_ _01752_ _01753_ VGND VGND VPWR VPWR _01754_ sky130_fd_sc_hd__o21a_1
XFILLER_0_157_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12795_ _02660_ _02733_ VGND VGND VPWR VPWR _02734_ sky130_fd_sc_hd__nor2_1
X_15583_ _05626_ _05625_ VGND VGND VPWR VPWR _05700_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17322_ _07226_ _07611_ VGND VGND VPWR VPWR _07612_ sky130_fd_sc_hd__xor2_2
XFILLER_0_141_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14534_ _04540_ _04542_ _04545_ VGND VGND VPWR VPWR _04546_ sky130_fd_sc_hd__o21ai_1
X_11746_ _01682_ _01684_ VGND VGND VPWR VPWR _01685_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17253_ net311 _06468_ _07461_ _07535_ VGND VGND VPWR VPWR _07537_ sky130_fd_sc_hd__a31o_1
X_14465_ _04437_ _04466_ _04469_ VGND VGND VPWR VPWR _04470_ sky130_fd_sc_hd__a21oi_1
X_11677_ _01598_ _01597_ VGND VGND VPWR VPWR _01616_ sky130_fd_sc_hd__and2b_1
XFILLER_0_36_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16204_ _06327_ _06331_ _06382_ VGND VGND VPWR VPWR _06383_ sky130_fd_sc_hd__a21o_1
XFILLER_0_141_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13416_ net237 _02546_ _03370_ _03372_ VGND VGND VPWR VPWR _03373_ sky130_fd_sc_hd__a31oi_1
X_10628_ net405 _05138_ _05149_ VGND VGND VPWR VPWR _00567_ sky130_fd_sc_hd__and3_2
X_14396_ _03895_ _04389_ _04392_ VGND VGND VPWR VPWR _04394_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17184_ net332 _06351_ _06437_ net316 VGND VGND VPWR VPWR _07461_ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13347_ _03297_ _03299_ VGND VGND VPWR VPWR _03300_ sky130_fd_sc_hd__nand2_1
X_16135_ _06269_ _06306_ _01784_ VGND VGND VPWR VPWR _06307_ sky130_fd_sc_hd__o21ai_4
X_10559_ _08086_ _00325_ VGND VGND VPWR VPWR _00498_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_47_Left_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16066_ _08834_ _06207_ _07382_ VGND VGND VPWR VPWR _06231_ sky130_fd_sc_hd__o21a_1
X_13278_ _03163_ _03164_ VGND VGND VPWR VPWR _03231_ sky130_fd_sc_hd__xnor2_1
X_12229_ _02119_ _02167_ VGND VGND VPWR VPWR _02168_ sky130_fd_sc_hd__xnor2_2
X_15017_ _05074_ _05075_ _05076_ VGND VGND VPWR VPWR _05077_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_75_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16968_ _07219_ _07220_ _07222_ VGND VGND VPWR VPWR _07223_ sky130_fd_sc_hd__a21bo_1
X_18707_ _09106_ _09134_ _09135_ VGND VGND VPWR VPWR _09136_ sky130_fd_sc_hd__a21boi_4
X_15919_ _03857_ _06068_ VGND VGND VPWR VPWR _06069_ sky130_fd_sc_hd__nor2_1
X_16899_ _07115_ _07145_ _07146_ VGND VGND VPWR VPWR _07147_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_56_Left_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18638_ _09053_ _09059_ VGND VGND VPWR VPWR _09060_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18569_ _06131_ _08978_ VGND VGND VPWR VPWR _08984_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_65_Left_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_74_Left_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09707_ _04115_ VGND VGND VPWR VPWR _04126_ sky130_fd_sc_hd__buf_4
X_09638_ net51 _03358_ _03391_ net262 VGND VGND VPWR VPWR _00011_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11600_ _01535_ _01538_ VGND VGND VPWR VPWR _01539_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12580_ _02386_ _02388_ VGND VGND VPWR VPWR _02519_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11531_ net377 _00815_ VGND VGND VPWR VPWR _01470_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_83_Left_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14250_ _04231_ _04232_ net434 net137 VGND VGND VPWR VPWR _04233_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11462_ _01387_ _01399_ _01341_ _01400_ VGND VGND VPWR VPWR _01401_ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13201_ _03151_ _03153_ VGND VGND VPWR VPWR _03154_ sky130_fd_sc_hd__and2_1
X_10413_ _00350_ _00351_ VGND VGND VPWR VPWR _00352_ sky130_fd_sc_hd__or2b_1
X_14181_ _04155_ _04067_ _04153_ _04154_ VGND VGND VPWR VPWR _04157_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_150_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11393_ _01290_ _01294_ VGND VGND VPWR VPWR _01332_ sky130_fd_sc_hd__and2_1
X_13132_ _03077_ _03078_ VGND VGND VPWR VPWR _03079_ sky130_fd_sc_hd__nor2_1
X_10344_ _00277_ _00276_ VGND VGND VPWR VPWR _00283_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13063_ _02994_ _03001_ _03002_ VGND VGND VPWR VPWR _03004_ sky130_fd_sc_hd__o21ai_2
X_17940_ _08283_ _08290_ _08291_ VGND VGND VPWR VPWR _08292_ sky130_fd_sc_hd__nor3_2
X_10275_ _00212_ _00213_ VGND VGND VPWR VPWR _00214_ sky130_fd_sc_hd__nand2_1
X_12014_ _01848_ _01861_ VGND VGND VPWR VPWR _01953_ sky130_fd_sc_hd__nor2_1
X_17871_ _08204_ _08214_ _08215_ _08133_ VGND VGND VPWR VPWR _08216_ sky130_fd_sc_hd__a211oi_1
XPHY_EDGE_ROW_92_Left_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16822_ _07051_ _07054_ VGND VGND VPWR VPWR _07062_ sky130_fd_sc_hd__xor2_1
Xfanout490 net491 VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__buf_2
X_16753_ _06894_ _06985_ VGND VGND VPWR VPWR _06987_ sky130_fd_sc_hd__nor2_1
X_13965_ _03926_ _03929_ _03936_ VGND VGND VPWR VPWR _03937_ sky130_fd_sc_hd__a21oi_1
Xmax_cap4 _05188_ VGND VGND VPWR VPWR net538 sky130_fd_sc_hd__buf_1
X_15704_ net466 net191 net176 net483 VGND VGND VPWR VPWR _05833_ sky130_fd_sc_hd__a22oi_1
X_12916_ _02849_ _02854_ VGND VGND VPWR VPWR _02855_ sky130_fd_sc_hd__and2_1
X_16684_ net312 _06319_ VGND VGND VPWR VPWR _06911_ sky130_fd_sc_hd__nand2_1
X_13896_ _03268_ _03860_ _03862_ VGND VGND VPWR VPWR _03863_ sky130_fd_sc_hd__a21o_1
X_18423_ _08772_ _08774_ _08577_ VGND VGND VPWR VPWR _08824_ sky130_fd_sc_hd__o21a_1
X_15635_ net462 net187 _05746_ _05745_ VGND VGND VPWR VPWR _05757_ sky130_fd_sc_hd__a31o_1
X_12847_ net264 _01798_ _02785_ VGND VGND VPWR VPWR _02786_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18354_ _08740_ _08747_ _08620_ VGND VGND VPWR VPWR _08748_ sky130_fd_sc_hd__o21a_1
X_15566_ net469 net179 net176 net474 VGND VGND VPWR VPWR _05681_ sky130_fd_sc_hd__a22oi_1
X_12778_ _02712_ _02713_ _02715_ VGND VGND VPWR VPWR _02717_ sky130_fd_sc_hd__nand3_1
X_17305_ net281 _07183_ _07592_ VGND VGND VPWR VPWR _07594_ sky130_fd_sc_hd__a21oi_1
X_14517_ net429 net567 net161 net155 VGND VGND VPWR VPWR _04527_ sky130_fd_sc_hd__and4_1
XFILLER_0_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11729_ _01456_ _01459_ _01405_ _01667_ VGND VGND VPWR VPWR _01668_ sky130_fd_sc_hd__a211o_1
X_18285_ _08668_ _08670_ VGND VGND VPWR VPWR _08672_ sky130_fd_sc_hd__and2_1
X_15497_ _05526_ _05549_ _05604_ VGND VGND VPWR VPWR _05605_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17236_ _07467_ _07468_ _07466_ VGND VGND VPWR VPWR _07518_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_154_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14448_ net413 net170 net165 net417 VGND VGND VPWR VPWR _04451_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_3_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17167_ _07430_ _07441_ VGND VGND VPWR VPWR _07442_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_142_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14379_ _04343_ _04373_ _04286_ _04374_ VGND VGND VPWR VPWR _04375_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_12_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16118_ _01705_ _01736_ _01871_ VGND VGND VPWR VPWR _06288_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_110_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17098_ _07238_ _07242_ _07236_ VGND VGND VPWR VPWR _07366_ sky130_fd_sc_hd__a21bo_1
X_16049_ _06210_ _06211_ VGND VGND VPWR VPWR _06212_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10060_ _07976_ _07998_ VGND VGND VPWR VPWR _08009_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13750_ _03707_ _03713_ VGND VGND VPWR VPWR _03716_ sky130_fd_sc_hd__and2_1
X_10962_ _00822_ _00900_ VGND VGND VPWR VPWR _00901_ sky130_fd_sc_hd__nand2_1
X_12701_ _02639_ VGND VGND VPWR VPWR _02640_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13681_ _03643_ _03644_ VGND VGND VPWR VPWR _03645_ sky130_fd_sc_hd__xor2_1
X_10893_ _00742_ _00741_ _00725_ VGND VGND VPWR VPWR _00832_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_156_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15420_ _05492_ _05516_ _05518_ VGND VGND VPWR VPWR _05520_ sky130_fd_sc_hd__and3_1
X_12632_ _02565_ _02563_ VGND VGND VPWR VPWR _02571_ sky130_fd_sc_hd__xor2_1
XFILLER_0_109_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12563_ _02500_ _02495_ _02499_ VGND VGND VPWR VPWR _02502_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15351_ _05333_ _05388_ VGND VGND VPWR VPWR _05444_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14302_ _04288_ _04256_ _04286_ VGND VGND VPWR VPWR _04290_ sky130_fd_sc_hd__nor3_1
XFILLER_0_81_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11514_ _01450_ _01452_ VGND VGND VPWR VPWR _01453_ sky130_fd_sc_hd__and2_1
XFILLER_0_136_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18070_ _08048_ _08432_ VGND VGND VPWR VPWR _08435_ sky130_fd_sc_hd__and2b_1
XFILLER_0_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12494_ _02430_ _02432_ VGND VGND VPWR VPWR _02433_ sky130_fd_sc_hd__and2_1
X_15282_ _05362_ _05367_ VGND VGND VPWR VPWR _05368_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17021_ net320 _06352_ net270 VGND VGND VPWR VPWR _07281_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14233_ _04212_ _04153_ _04157_ VGND VGND VPWR VPWR _04215_ sky130_fd_sc_hd__and3_1
X_11445_ _01371_ _01383_ VGND VGND VPWR VPWR _01384_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14164_ _04136_ _04138_ VGND VGND VPWR VPWR _04139_ sky130_fd_sc_hd__xnor2_1
X_11376_ _01248_ _01270_ _01269_ VGND VGND VPWR VPWR _01315_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_156_Right_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10327_ _00181_ _00177_ _00180_ VGND VGND VPWR VPWR _00266_ sky130_fd_sc_hd__nor3_1
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13115_ net211 _02746_ _03060_ VGND VGND VPWR VPWR _03061_ sky130_fd_sc_hd__and3_1
X_18972_ _04213_ _09270_ _09271_ _09275_ _09277_ VGND VGND VPWR VPWR _09427_ sky130_fd_sc_hd__a32o_1
X_14095_ _04035_ _04046_ _04065_ _04066_ VGND VGND VPWR VPWR _04067_ sky130_fd_sc_hd__o211a_1
X_13046_ _02982_ _02984_ VGND VGND VPWR VPWR _02985_ sky130_fd_sc_hd__nor2_1
X_17923_ net331 _06890_ _07182_ net314 VGND VGND VPWR VPWR _08274_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10258_ _00193_ _00196_ VGND VGND VPWR VPWR _00197_ sky130_fd_sc_hd__xnor2_1
X_17854_ _08087_ _08194_ _08197_ VGND VGND VPWR VPWR _08198_ sky130_fd_sc_hd__o21ba_1
X_10189_ _08097_ _06645_ _08372_ VGND VGND VPWR VPWR _09428_ sky130_fd_sc_hd__o21ai_1
X_16805_ _06935_ _07043_ VGND VGND VPWR VPWR _07044_ sky130_fd_sc_hd__nand2_1
X_17785_ net291 _02932_ VGND VGND VPWR VPWR _08122_ sky130_fd_sc_hd__nand2_1
X_14997_ _05051_ _05052_ _05054_ VGND VGND VPWR VPWR _05055_ sky130_fd_sc_hd__a21o_1
X_16736_ _06882_ _06967_ VGND VGND VPWR VPWR _06968_ sky130_fd_sc_hd__nor2_1
X_13948_ _03909_ _03919_ VGND VGND VPWR VPWR _03920_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16667_ net278 _06723_ _06803_ net274 VGND VGND VPWR VPWR _06892_ sky130_fd_sc_hd__a22oi_1
X_13879_ _03670_ _03715_ _03717_ _03844_ VGND VGND VPWR VPWR _03845_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_9_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18406_ _08792_ _08794_ _08620_ VGND VGND VPWR VPWR _08805_ sky130_fd_sc_hd__nand3_1
X_15618_ net469 net473 net183 net179 VGND VGND VPWR VPWR _05738_ sky130_fd_sc_hd__and4_1
X_16598_ _06812_ _06815_ VGND VGND VPWR VPWR _06816_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18337_ _08682_ _08686_ _08727_ VGND VGND VPWR VPWR _08729_ sky130_fd_sc_hd__and3_1
X_15549_ _05634_ _05661_ VGND VGND VPWR VPWR _05662_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18268_ _08650_ _08652_ VGND VGND VPWR VPWR _08653_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17219_ _07478_ _07479_ _07498_ VGND VGND VPWR VPWR _07499_ sky130_fd_sc_hd__and3_2
XFILLER_0_31_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18199_ i_error\[6\] _08574_ _08575_ VGND VGND VPWR VPWR _08577_ sky130_fd_sc_hd__nand3_1
Xfanout6 _07571_ VGND VGND VPWR VPWR net540 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_123_Right_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09972_ net344 net520 _05149_ VGND VGND VPWR VPWR _07041_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11230_ _01152_ _01166_ _01168_ VGND VGND VPWR VPWR _01169_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_132_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11161_ _01098_ _01099_ VGND VGND VPWR VPWR _01100_ sky130_fd_sc_hd__nor2_1
X_10112_ net342 _05193_ _08570_ VGND VGND VPWR VPWR _08581_ sky130_fd_sc_hd__a21oi_1
X_11092_ _01025_ _01028_ _01030_ VGND VGND VPWR VPWR _01031_ sky130_fd_sc_hd__a21o_1
X_10043_ _07272_ _07778_ VGND VGND VPWR VPWR _07822_ sky130_fd_sc_hd__xor2_1
X_14920_ _04798_ _04959_ _04966_ VGND VGND VPWR VPWR _04970_ sky130_fd_sc_hd__o21ai_1
Xhold40 i_error\[18\] VGND VGND VPWR VPWR net547 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 kp\[7\] VGND VGND VPWR VPWR net558 sky130_fd_sc_hd__dlygate4sd3_1
X_14851_ _04789_ _04893_ VGND VGND VPWR VPWR _04894_ sky130_fd_sc_hd__nand2_1
X_13802_ _03756_ _03767_ VGND VGND VPWR VPWR _03768_ sky130_fd_sc_hd__nand2_1
X_17570_ net323 _06718_ _06719_ VGND VGND VPWR VPWR _07885_ sky130_fd_sc_hd__and3_2
X_14782_ _04816_ _04817_ VGND VGND VPWR VPWR _04818_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11994_ net223 _01930_ _01932_ VGND VGND VPWR VPWR _01933_ sky130_fd_sc_hd__a21oi_1
X_16521_ _06710_ _06730_ VGND VGND VPWR VPWR _06731_ sky130_fd_sc_hd__and2b_1
X_13733_ _03697_ _03698_ VGND VGND VPWR VPWR _03699_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_11_Left_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10945_ _00877_ _00882_ _00883_ VGND VGND VPWR VPWR _00884_ sky130_fd_sc_hd__o21a_1
XFILLER_0_86_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19240_ clknet_4_13_0_clock _00122_ VGND VGND VPWR VPWR i_error\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16452_ _06651_ _06652_ VGND VGND VPWR VPWR _06655_ sky130_fd_sc_hd__nor2_1
X_13664_ net237 _02935_ _03623_ _03626_ VGND VGND VPWR VPWR _03627_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_38_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10876_ _00814_ VGND VGND VPWR VPWR _00815_ sky130_fd_sc_hd__clkbuf_4
X_15403_ _05488_ _05499_ _05500_ VGND VGND VPWR VPWR _05502_ sky130_fd_sc_hd__nand3_1
XFILLER_0_144_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12615_ _02540_ _02553_ VGND VGND VPWR VPWR _02554_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19171_ _09550_ _09074_ _09581_ net491 VGND VGND VPWR VPWR _00140_ sky130_fd_sc_hd__o211a_1
X_16383_ _06486_ _06578_ VGND VGND VPWR VPWR _06580_ sky130_fd_sc_hd__and2_1
X_13595_ _03501_ _03548_ VGND VGND VPWR VPWR _03554_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18122_ _08476_ _08466_ VGND VGND VPWR VPWR _08492_ sky130_fd_sc_hd__xnor2_2
X_15334_ _05420_ _05422_ _05425_ VGND VGND VPWR VPWR _05426_ sky130_fd_sc_hd__o21ai_1
X_12546_ _02372_ _02484_ VGND VGND VPWR VPWR _02485_ sky130_fd_sc_hd__xor2_1
XFILLER_0_124_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18053_ _08403_ _08404_ _08414_ _08415_ VGND VGND VPWR VPWR _08417_ sky130_fd_sc_hd__a211o_1
XFILLER_0_123_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15265_ _05345_ _05349_ VGND VGND VPWR VPWR _05350_ sky130_fd_sc_hd__and2_1
X_12477_ _02405_ _02414_ _02415_ VGND VGND VPWR VPWR _02416_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_124_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_4 net563 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17004_ net274 _07183_ VGND VGND VPWR VPWR _07263_ sky130_fd_sc_hd__nand2_1
X_14216_ _03902_ _03907_ _04195_ VGND VGND VPWR VPWR _04196_ sky130_fd_sc_hd__o21a_1
XFILLER_0_151_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11428_ net377 net374 _00408_ _00514_ VGND VGND VPWR VPWR _01367_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_20_Left_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15196_ net423 net198 _05272_ _05273_ VGND VGND VPWR VPWR _05274_ sky130_fd_sc_hd__a31o_1
XFILLER_0_111_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14147_ _04118_ _04119_ VGND VGND VPWR VPWR _04120_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11359_ _01297_ _01239_ VGND VGND VPWR VPWR _01298_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14078_ net415 net140 net134 net418 VGND VGND VPWR VPWR _04050_ sky130_fd_sc_hd__a22o_1
X_18955_ _09257_ _09408_ VGND VGND VPWR VPWR _09409_ sky130_fd_sc_hd__xnor2_1
X_13029_ _02907_ _02905_ VGND VGND VPWR VPWR _02968_ sky130_fd_sc_hd__and2b_1
X_17906_ _08187_ _08200_ _08199_ VGND VGND VPWR VPWR _08255_ sky130_fd_sc_hd__o21ai_1
X_18886_ _09330_ _09331_ VGND VGND VPWR VPWR _09333_ sky130_fd_sc_hd__nand2_1
X_17837_ _08177_ _08178_ VGND VGND VPWR VPWR _08179_ sky130_fd_sc_hd__xor2_1
Xrebuffer16 _07966_ VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__clkbuf_1
Xrebuffer27 _08738_ VGND VGND VPWR VPWR net534 sky130_fd_sc_hd__clkbuf_1
X_17768_ _07984_ _07985_ _07990_ VGND VGND VPWR VPWR _08103_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16719_ _06847_ _06948_ VGND VGND VPWR VPWR _06949_ sky130_fd_sc_hd__xnor2_1
X_17699_ _07936_ _07939_ VGND VGND VPWR VPWR _08027_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_147_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09955_ net348 _05193_ _06821_ _06843_ VGND VGND VPWR VPWR _06854_ sky130_fd_sc_hd__and4_1
X_09886_ net342 _06073_ _05336_ net344 VGND VGND VPWR VPWR _06095_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_79_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10730_ net371 _05996_ VGND VGND VPWR VPWR _00669_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10661_ _00513_ _04291_ VGND VGND VPWR VPWR _00600_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_126_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12400_ _02321_ _02336_ _02313_ VGND VGND VPWR VPWR _02339_ sky130_fd_sc_hd__o21a_1
X_13380_ _03303_ _03332_ VGND VGND VPWR VPWR _03333_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10592_ _00434_ _00530_ VGND VGND VPWR VPWR _00531_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12331_ _01973_ _01974_ VGND VGND VPWR VPWR _02270_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15050_ _05111_ _05112_ VGND VGND VPWR VPWR _05113_ sky130_fd_sc_hd__and2_1
X_12262_ _02191_ _02200_ VGND VGND VPWR VPWR _02201_ sky130_fd_sc_hd__or2_1
X_14001_ net425 net137 net136 net430 VGND VGND VPWR VPWR _03973_ sky130_fd_sc_hd__a22oi_1
X_11213_ _01144_ _01150_ _01151_ VGND VGND VPWR VPWR _01152_ sky130_fd_sc_hd__o21ai_1
X_12193_ _02127_ _02130_ VGND VGND VPWR VPWR _02132_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11144_ _01006_ _01008_ VGND VGND VPWR VPWR _01083_ sky130_fd_sc_hd__or2_1
Xoutput85 net85 VGND VGND VPWR VPWR out_clocked[14] sky130_fd_sc_hd__clkbuf_4
Xoutput96 net96 VGND VGND VPWR VPWR out_clocked[7] sky130_fd_sc_hd__buf_2
XFILLER_0_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18740_ _08924_ _09075_ _09077_ VGND VGND VPWR VPWR _09172_ sky130_fd_sc_hd__nand3_1
X_15952_ _06065_ _06103_ _06104_ VGND VGND VPWR VPWR _06105_ sky130_fd_sc_hd__a21o_1
X_11075_ _00991_ _01013_ VGND VGND VPWR VPWR _01014_ sky130_fd_sc_hd__nor2_1
X_10026_ _05479_ _05853_ VGND VGND VPWR VPWR _07635_ sky130_fd_sc_hd__xnor2_2
X_14903_ _04948_ _04950_ VGND VGND VPWR VPWR _04952_ sky130_fd_sc_hd__and2_1
X_18671_ _08803_ _08743_ VGND VGND VPWR VPWR _09096_ sky130_fd_sc_hd__nor2_1
X_15883_ _05992_ _05981_ _05982_ VGND VGND VPWR VPWR _06030_ sky130_fd_sc_hd__nor3_1
X_17622_ _07828_ _07830_ VGND VGND VPWR VPWR _07942_ sky130_fd_sc_hd__nor2_1
X_14834_ _04766_ _04875_ VGND VGND VPWR VPWR _04876_ sky130_fd_sc_hd__nand2_1
X_17553_ _07548_ _07549_ _07600_ VGND VGND VPWR VPWR _07867_ sky130_fd_sc_hd__o21a_1
X_14765_ _04794_ _04799_ VGND VGND VPWR VPWR _04800_ sky130_fd_sc_hd__nand2_1
X_11977_ _01897_ _01900_ _01902_ VGND VGND VPWR VPWR _01916_ sky130_fd_sc_hd__or3_1
XFILLER_0_58_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16504_ net289 _06410_ _06402_ net286 VGND VGND VPWR VPWR _06713_ sky130_fd_sc_hd__a22oi_1
X_13716_ _03431_ _03680_ _03681_ VGND VGND VPWR VPWR _03682_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10928_ _00760_ _00863_ VGND VGND VPWR VPWR _00867_ sky130_fd_sc_hd__xor2_1
X_17484_ _06398_ _07571_ _07788_ VGND VGND VPWR VPWR _07791_ sky130_fd_sc_hd__o21ba_1
X_14696_ _04722_ _04723_ net436 net161 VGND VGND VPWR VPWR _04724_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_156_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19223_ clknet_4_5_0_clock _00105_ VGND VGND VPWR VPWR prev_error\[10\] sky130_fd_sc_hd__dfxtp_2
X_16435_ _06628_ _06632_ _06635_ VGND VGND VPWR VPWR _06637_ sky130_fd_sc_hd__and3_1
X_13647_ _03556_ _03607_ VGND VGND VPWR VPWR _03608_ sky130_fd_sc_hd__nand2_2
X_10859_ _00408_ VGND VGND VPWR VPWR _00798_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19154_ net506 _09442_ VGND VGND VPWR VPWR _09572_ sky130_fd_sc_hd__nand2_1
X_16366_ net290 net287 _06328_ VGND VGND VPWR VPWR _06561_ sky130_fd_sc_hd__and3_1
X_13578_ _03511_ _03514_ VGND VGND VPWR VPWR _03537_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18105_ _08457_ _08469_ _08467_ _08468_ VGND VGND VPWR VPWR _08474_ sky130_fd_sc_hd__a211o_1
XFILLER_0_26_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15317_ _05405_ _05406_ net482 net153 VGND VGND VPWR VPWR _05407_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_81_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12529_ _02463_ _02467_ VGND VGND VPWR VPWR _02468_ sky130_fd_sc_hd__nor2_1
X_19085_ net498 prev_error\[4\] VGND VGND VPWR VPWR _09529_ sky130_fd_sc_hd__or2_1
XFILLER_0_140_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16297_ net270 _06452_ _06484_ _06482_ VGND VGND VPWR VPWR _06485_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_2_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18036_ _08234_ _08378_ VGND VGND VPWR VPWR _08398_ sky130_fd_sc_hd__nand2_1
X_15248_ _05326_ _05330_ VGND VGND VPWR VPWR _05331_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15179_ _05153_ _05254_ VGND VGND VPWR VPWR _05255_ sky130_fd_sc_hd__or2_1
Xfanout308 ki\[6\] VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__clkbuf_4
Xfanout319 net321 VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__clkbuf_4
X_09740_ net76 net18 VGND VGND VPWR VPWR _04489_ sky130_fd_sc_hd__and2b_1
X_18938_ _09389_ _09313_ _02146_ VGND VGND VPWR VPWR _09390_ sky130_fd_sc_hd__o21a_1
.ends

